`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 5248 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/9huKRhRMtvnNqb3Z+UU7TahEoHV+T8U3P3ufru7l1O
3DlgtZzb9QxCbOjthp9+wDkjygH0eUfDrEl1ovhZG631fscPLVJ+KF4bO5YocKzY
CriN4E1RhE4IKyONpxBwkCdqBPfFHBU5X/qMZVrgQ3ehvLcmGascO46ga6yQMRBj
Jlom/YkL90duOnNtfZ1Oqj28VEO6uR54BHfkD5L4TetdJrw03Nkf26ntO9bz65NW
PDh1inhOhZ2rP056KKWXxTutKNhNj8coGkvgvBaxmcfURKWUjL35ocLOfBPWVp5Q
a2EmY63V7yp0YRmazuXyEOBT4CaLvAP+ZmoUjaIwjKbYXhx6K2wkcXEhWxTskqvV
Qkq+/yaDoRDrgaWczVlcgnSlllnrLcdIhW9kgLhJkRL/3XF2DUPiIYRQdcIhd3nl
WEbN1epJdDu7/c/CgN81UYzA+yXWHHYTx55X9stoBk5WCSbSjwaDLpYhz36Rsyut
9ihgZ8o91xkRX599rnr8vZ/6sb9Zl4uBcLwDa/gPqP3OPUFHIzd//pz+Fvq9gEGI
v2hpBK7VBHyL6kzTHqmt7XId49lNmYzanZW1XdgvQBzDJBmVyMlxa4Z3SbM+j00K
lIy8tzEAeiRnWMU90GgUTVnlO4przoKU2FDAxD2unJIrnbLXudCC5vnkeT83YHWg
KUR9vQEI/rhS/fbGUp5PDwQOQTeZzGjIn6rlu/n9nHv2jgAzEmbGDr6M8kLQzF5U
7pK3SI5gXLvftM241Hf1J+GZ/Zmi1tCvfqjdXinfgD8btnJvVERq2FoLUJqjhbEj
yE1da5CJHA1hYploW2fG3tVDoOYCFbFPprtk7NihJzU2ie/wrdaGkb3Ekl9bcf73
GnNoomsCTD39tU9ZMOjYIa4zysLwanGHE2vmMGHf+Fny8haK6pgrA+CCtcm5KITS
uNPqIj3xPkq8F9LThdKrGNqB/yysyqMSSX40Ea/OiyCag6PGatAd9Zk10iXmF8Ky
xPo7tSXE3O1avW2e2PkKjMrNnM4+qZkLSeVx4WhMpMlN6uoXZxIq9LuRABNxdFI1
xSPzEGn7cTMTCuKdZ+J4PtD043Ykf7ExNAFRpLfcKN1ZCIvtYvUltb+yyQPme3Nr
robMwFjDhgl6SC4WBP92m81dRR8v4JmAt72Cvj/J9QcUxGxtmpSKGVAy4Q+3uz1t
wuPWt5IC0PUHyFs6I3xH+zGcqeQ8Q0lE0frRsQRcVuiZTw1pUry2mv3Fg+4ewNZ5
tdyS1vWjG12McCtYcixdl2g24ASjpRQ0IssAFUR8Rx6Vm+bmFQQvAtcpLKkG4RmN
sE3wtP/dpS/Tp2/0E5aKfH23cFWXuK06gyiOewjb+1jWAclZG6KT0tEgWoHC31ed
KUN1aWU2YOoEnOmBMwLK/Y/2ni5pPGqWnEK5Zoqa4s8usTbBDCTuDATW3xSe/x1s
fIE8JBWquU/pbGc8HN9gcU8/sy09fiXvdOzspYMPl6Lvs7SOxZjLGyu3gbFqNOzj
QNLWvM159xpcg/MY9kKZt/bGPHnNzeY6mi+2A6xXYZL8UD8sHuXs9MEhs7TrA2yp
Sx+JqW59/c6CH0ojw0NQhvLXpfXin9ZrzZqhI955B3G4saVC+vOKYL1dCLzubdtt
The+q95qtj5+7zSNFm35lXa6YP8cVCT+erIeAgIjY16Am6vUai9bZfkiSC+7XWk9
mAFE3afYxaXhIHJGBB61bidylEwdANp8/0OkG1lQ95+s7y2vHUKaKRYkk376fMR+
qIRSli9ZHzVOS2GNvOzpiQ3tbUBDhSgY7c9+CjKosj+yxw14xz1CBzn2tTTHv9eW
seDhBh7yfRt4JdiUPUQgM/s6W3SSfaWqdWywT/hnE8RskfEXALuoQ4FS8aeh1ceI
uboC8sEZRlCyBkn5SJ7iZ5s8yJDPZE+ou7OvM749FURidNInT/eX8KsOiEkSlGfR
YOV4T1MTBo3RnMIF/BgTzd39UvqJuMCxhaTmfaPrdfRgr/In32Wv4/rQ2zj3xGy4
sS/U7KYPxTLlbkQDdCV4tMzXY77pSyjXDQaxMk28qq1rHnnQ94GO2z2s/3vEZDKL
Itvpdceb5vzPuGpzBdyBlE5xrue6Q+ciP+FP4oDmw/bIC3t8fIvTP9IrTeFmqSHW
+z3Jn+opc1sNufEg9qzA0mB6X3pnuwWFcHrfZYyOcG5zcXq8K86QOPqEEOBbjnQZ
KToWrGDXK973sjMj0cS55tsc0kyzTyRudTi+R694AV/EnW5EgNMxWrTzGIkHzIDk
8tJAuYviboeSPmU+f3Hdt4U1eucP2RPvTkJdKWZhrjGWdtZv7Qill60zRD5AlFMu
0g+kjb94aKZ+Iy2yQmeWYs7OPHr+eAn7svOSHnU2Nv9dJOEIFLwf3e6Hpr9Bqjc+
bLbXW/F0lvXUw8f0kZvmm27z2q6/+Trz/w9JTXQl1EClz24k99ZLd7Ehpei0Sp7o
2vQd3AnKF4P0BTH9J9KCr1Cq7DqeONBSywyhMs6owwU/nq5hQ2wE2D9S1z9Iks95
9WjYZEbSdtJ+pzTNvEEsGZKYoGo2sstRUHZ9a4Kqjjs2WD3TUOhn28RlZnsWPAGE
49nl8hwXU/kMm1fHyyOkBx+iXC6LDuw7FwJQ1797lDcTG8trXAmpmeyCslxITOh/
kF+0fjb0GTMRtHaUvfaEFUNkUwg7LyOySl0o9ZsRp61uAh5LHi+elJiZQCyc8izO
9U1X4eY7T8Zh0G1/XzbgZwxOX1laHEnl57ZAc81yw6RTMguVStVhWCOeatg0eTbI
wkEHrfoCpN97++LPg8Y9otUCDIIbrU8+0PKsCZYib/9qOr9jyn1JE8POCnt/3ZIm
MG0fKNUJY0rkcGvJppIJGhK5amG0IgJaq/prZQRyWLgiPoSXCBk6LpmElb0yIExa
EnjH+SCB6c1YmjG/6YG/6EBvXXZDLhaEbax6EQ0SrtQi8wt0eQoDY08xMbke9bZX
pcBrl/4lF70+B8fUI8Sv9Fi9hwGYqUxSjUs1022Qzw2751IG1+83dexP6FTeI9ud
3FK18KXMh6179QzuY1uY5CISheIFpXiYj4flkvA1YufW7q4n4/8SQn1bW1SRs9pp
dwrUcyYiH6NWuCMxZcFwihNH+iMfV+fD2ihkZ8n5xyWRA3fU7KIeH5D24R73uMmE
2s1ifWQn/zN4tE7qowYQvS00lR+Q04VNZupqUzesBAvDO38fDIoV9z+MBTf8b2/t
MFnebL9Yn9hH+BYztVGzNSU+wayqhcYtts+VWyJUYvKgKha+IhbdDfDjI1ed8HTa
asoz8RSDX+AtexykeXwy4Fkw9EJhMyMAG+0ZKRQz/tmVXsqbPMJUIx1Fr++3X++v
l7e4K/uZWMUr+sTS+QV1S9z/UhPExot1L2uLRwP9Zw3r5AO28O1c2/xsoaVfd9CE
pDxjFLOEmwiYVJKCe5Y1CDlDh2Id36w/Q9s1z+2wfqqL+klldokUc6nwww2GFbic
0O8pF8X2R8BVraJ1DLkJqBkA0dU4U4ZyFIiGj+DTFQiD/lpRmCeNgUSN/xWPWI51
wQjkEir9HT93xRpwIY4KYglQGLHXJWJdekVhmEFkohJZi9dPDIS7+xZgdCAsf8Xl
nxtoDUwBBoKyajIb3MdXZq/3OcfZcWFxVzPDsXpeqMgQu1rzgkirx9DjrVweQm/1
XVyY08Z2letJ8/MpWw6+jT83FciEhOEtma4M+4y3lT3NR1PFs1rFNt8eD5hQ2+mt
6ZBdRLxQ58O3YgBuvmUk0r0CSEmWEpP7n+jG8eypeUMrtYV3hUvr3mTWlyThFHTE
3L/1oK2ItxwMbrf1HW8kK0QLAcl3/XyfQN6Kb8HSe5s2HB3W9DrdLXfMfNrCF3FD
5LCaM4XhZwC3+BcKuvytdBTlEZSGbDE5CGgTHdI7m9MdtqPQW2Yq2E2ADutq4QLc
4IP3cUd1MWdzimS9NX4Unm4FtzwiXgcoiuZHhegfCiYGka/NEn4HBWxQswapZHRH
fW5oaob3HovVJ0z08p0xjvmEINBG2MOHlfKtoqnvvzMWHHxmJ3WxCZLivMagHijY
1rFc8cby5IaJ4slkrWN+eOaL4J1TDJGAupGCTNnGFChXOMKzBuaQINJZ/V/9l5no
JoRfXFySaU4I8Yotv5jIZpRHFfmFZSUzMmWVOawfZ8/yJ2LdXt4U9cjyBPamVaHs
QPBETi7X0LBkyPf8wSqyV10usmHsLaTsVjBK1y+JZt2jJ4aP02cbQOZS5jeLm9H7
hsl6D+uk2Tw1rccNJKUlUl+/IkDeB4SZPgEUJWtCPLh0WlX/a3Yy+iSmOb9YHFNV
LsnnRb/XYkIKFYxyHUGgCtNJlJELYEPQnQuSBAgLdcdAeqE+P5pYflCFLHNkpKnf
NPydT2Hcr8xpFxbhXJ51Bp0q098hm1MtO2gC+8AwML9IBJqppvP1y+oPlD0yZwQY
Ujpy0/5gdUqNCHKB/+hbE7UdZ9nzHgcorYbi2eDKNJ96WHgaDJSG33EvFIyzDhcs
Ca3Mtng8wZp6myggBUTEmV3NXnt006nZxHueDLVpSAnAR2Am0Vbzvo1toylABYPU
4XEx+utzUe3YIkZS6Ym8JXliGAjYUhwynz7syJswmeb6RvrDxeNhGM7zplKQaaEK
cg4E2OtWKHiXRCLeuNyWcVyA6yx55PdU1WRng29cIx/y8vHk3KAR/H59SfRpkuIJ
T1qSVaOo0FIsze98vrPn/CDYshVg6F8LLALZl27LZHS6lvZF4tyWioWWyKMFxGRx
5UoPL1HjD6VezECd7CMWF8nd2EBbimT4VRjUgwRzi8ESYL5emrTVdcxSQB1DKltW
R3HJDNPBDHHi3xmsvD9kVm2ITPu3x08EH97+H01zglqT1IcdYGfOSJw85kn7WhQj
Bp3llJIJOwi/MJGcHY6ZxioR8I/ymnezv55SiLef55woiYhz/230HsuPSrYJI4BY
u9y+/QDRdy9epBlOk/EYoJ+Y9f6tMy/AHs7dO2TdCvuVT6wXQ3O98vM/kkuBsEuy
y6NdiKS5zlLadjOZvNZdt95j8aAb8Wuk1iIJHoycH214kidBZMHy9V4TplG0c3i7
QoSPXD5w7ggcb4B75fNq9kogdAoqxEj3kkLYrhymi6uXV6Pkq+f7jwmFQyBhwhQj
e1IPZQidVpGdUggCOuMCYpVqSQeFyjlplcwYSCHxyvtwZPNYo4s5OWH3mHLvOR5C
l8GCLLGTi3nce5pkaPfb5dT2bjN3oYDmt14phwhc6K66roTV4MKvrwHPoMJrr/ao
huXMdq3N8aJUMfK0YSSvy5MubNpI3konBuKh7UCA3B/f17SAvlnPCAUED18jQh9l
ikMzzXAXLXoym0drs6+67cllgWDNeK9Mkuft6drQkJ/Li9ysMyxJeGr60YfLTI5w
eTlww/iV9f5QVkdfEcRO8oczjQG4h80VHFNFuCTrx5Hy6l0t5H/9mFdE7m9ETzud
w6LcUwnNKufvZwizUh9rThZXB5IkrdG1tkcyvggNt+vRWsRsj/q72TnZRNq1sUW2
69cT2A8NcuEWSoWT0nHewbuRlFuBOlvAEjfAxwLEOgSChU/CZ2Sytfiqv0IOOPf4
vYTanC1npvdzLTm1EtxTuvDJ5B8J6Wkm8STD7SDIXN4w60k6bkM0zJJYh8T1fG0n
7uY6514bJhRZSGxDtKkgfMwQYXKKxoJJ/sirJhvo4n11N9G1yQfg8I8hDI27AgAy
o+LyzOLeSi0vCXIJ2MHBw+TPKwrr6Sm7rpF8f2fdklqpWYISuKFsTczclaXIgCzf
1vx3ieSsjQb7SMeLwQZ+T3Dv92ivRimD+JiiZNFQ8rjGpqxfS+ER5XN2xw0MFUGP
hA/BhBCRLqb9TJd/nQCyoVm/fPPcCIHsp197JysAl7cyuS11ur4toeuzVJjPIJik
8LN41xC812MYppwvD237l+Gz1HzzUxrVUIUpB1s0QNZrRpaIwI/ej5EgBKqlfOIi
GaR1xpqWQNI9qcGk2KzQhyYQoQiYlgielb5fS90plJhmz1s+/v80Aitm8thMf3qB
jqZ8qFiUg11NJw+0c4Txy5hl+lq4FEranqx8kDNyfDHT/2074gP+G2kyqMv7SCpI
2spKWWHhhBPIyz8b6oGeBVRSz/7s0sQAxECidWxA/DAxNtHBS0/ppmqMbRxwctTF
AUN7wtCinRgUqeLraOpiiUbPI5Z2QUWQwKGs9pjDWCuc6ae1sgLdPqxxV0X47AI0
iXH9t+NltTxECpLtRKWByqo+Luv6TSC0pVZUBsZeH283b8RhTSxnqhYFOY+Mef2e
DcnVWi0F6qd4C0Hl1mGQCUYeRmN837k28ffybd7qrD1Ad1eRjv2nBPNdspx76e4k
yqJhZwlapYNX6mOzpL0px6oHGk3NAJZcXoCT28zr9tXgVfTyd0N5bQIpZelgqrqV
8bKRfn2j5uEsqdEQzxfAxMMRqbWTkZca8uM955Y9kv0IdqgUBOtzpTmG/Eat6sXp
zuaq/Ik3eZq0WA9iIjfYqWhWlPz5yV+Q8k0CI0EXxeNwIXnppboyhn5QONFv/PfE
1pE+vSgf8oddvhRUAkAdmfvt/ke5dtaRSQWm21aOmVLWNI9Lv2DPtoNYLo2qpqjG
vZ29jeIELkZ2B3mJWpr1vtErx6zyjvp6J0Ff8Izs++qPhV0HfZNaWq7CB7a9VkM5
SqamedMzbrc+s0psTCVZ1x9/5Y08x5Pmd8i4e4N/tDY0GIK+pfcCpj+LdXO8gq1C
OJov8NJcUOnpzcHppugTOlJ7sWKftsEM7RpKs5+op3zPJbwE5Vw9lddWYCkBjvQh
k1OGIABjt5GpEkOFlMlIGSgwqZARftQvo22GMMTh4GYwDiG2mxQA58mYpkAP9WAr
WIMGufEUg3giCUAzauGq0UyRXeSV/6g+ftDNoDtpH7WSUlM+T1spgi4DagOXcMM5
pmo8BqrHD1m4/v8lta69zQ==
`protect end_protected