`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 2992 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/9huKRhRMtvnNqb3Z+UU7TahEoHV+T8U3P3ufru7l1O
3DlgtZzb9QxCbOjthp9+wDkjygH0eUfDrEl1ovhZG61ReK1tTLd+kH/e61F8qT9U
S20w+cDXONds/HAmuNx5SpGnGfBlc0gYgxLGziboppk7uR+DStqRVbDClWQvNL+b
q2dqg8Fdxu1HyZ5PsZbIQkGeDMcEdbmhDOT7FtGJLlspwmmqwpuR0iP6i8IqUQIh
jI9vI5q5lArAzCfpVTfs4ftPxAAqYcggxmUqDijQ9/86tEsFf66NMeG6+7TNZM5i
BuQZ5PJLuL9cKUtbyccq8779/ROv+W6VPTTaZEErnNHcQkUXMpvk3NhZ5siuflVo
GAtqWjzXP0mRT/51A2M5SeqOdDme74D+wBawy7ZOYiboVRTQAGLfGik6lw28ywwV
gEmdxRbqsLbiVg6o4OcICXOKDdryNjBseRN9Wu8q6nWEb2kKyRur1Aeh1pphwXuC
Kwvtm8iWIu8ssTzpVdJ5yfdTSEO5vWpNZjhv4mnTwoZ+H+l6y+43UE7/GHakrHa/
Q0Ld8n3/kIUlLQH+O/a9uqhBMpjMxGpm7WaJ2on7mnixQ/BIDbMr1TeOwPvkJqs2
Xwo6L2knacB+gNqYah18p2enB2NMreBmUyaWibu4PESUytq5/C7ncl3GSLbEHOgq
Sxpj/Iqlq5VHlVlx50727903KqJW0B1l+tOzqM99qLWgV25+9tZ2Gry9V7eM/ifT
+kFLfdAJHkJhyFLo3BKfgpCblDem5b9LBEO+87sg8xIOiKR8Yvn60TJeSLrNaKCz
vRwtEGbe7VSTLSrUqAyAZYB1/4zDvDS2TB2Ym6/6kBUVGb0GlBF+wqXfCBa6QUTP
yNfiTve5ljfyYbOlMrjBCW+CIkFLkTygDeygk+/fqE8SHscHVh76Pihwt6lwb03g
X7vCNMrVXsb4513V9bO2BdMFcv2DV2KXlmdeBIk8WZDdL9p6aWq7VYFp1G2asygI
ABnsIi/iHKtaNMOMP4jkNGrSyuzJSMEUYvSR4KBB1zx2+4DhZCU5eJs5rIUC8inR
diepjn4rA6NyAK2/JbqhgGmW9vlDdc8IGocSIWztwP8lKb54HsiouosFLSenFOLE
QUnj89r3sHMDGZ+BbxDcaBfhjuMcNpii9Ieu3ibqrQNqRZo8snYNsPC9PuUeDDXr
GrbrUuF1OLwCNK9+RpKyu/SGsEoiwFyyvs8d1fzCct6Odp4ureXEowr6vy4W6/uf
sAPAt/KtqaMptOxCZg9Ghxy5k5S2xtiPpEd6iO+suNPfVOgLPQO2FRrquED6nI3h
djXwa/Aklnq1E6q8lNdrlxSD5Ed3+E5rs6Ou+P4/+urrm2YrTr+Qo631IgEKRhh3
uoYuNISe6mjLQW8pKTjXA673tBmghovZpU+eNladVL8Edsy5diTYZAARjEFcZ3Yg
y4AeahkoGNUZX/rsCv3uJdrIugYu5StGnpuKho0VrhCMLOnO3JdDPgrbWusJiK1S
d584wCChNRO3gHp3xFXqUBQfarOQ5ibY3Zcjz0T6+P1PKrf1inhn7FBAlzQ94GXI
8XjMnY9IAfSqjCo5RXxCQ4oAouXVYLU3zLNw6GMsv6JBsv8d7OcfmiVKA2X1PmZy
6/N6HJXPlBlpt0lzxSl2S3JcA4VHmo1VMfTz5bnMPB+OWiQlLOMnSDnfFG19Om5Q
keDGgCZosiBK5kSAij88L8fJxfl/ERaLoVxcJV49ZncGTj5kqXSIT2NyqOhP3AeA
hTz+wti9beJSIo0l+NTWZUj9hdi2ynSBp43CHGkxuMpLeLlukbpAjTByapNw5LoM
EJZoKPW955Z7J9xh8kXQ4U896+0cTfHJ2ej1ZeVHV6CAb4/PKp2Q7W2zU1gwDKE0
xhqi2yNXyQVlt5blPUtiC/84ImQWzxDT8EpxAuq29C/tA+kv6XWKLmJNTOTLkRZ1
DiVbpRGxDf+PfYeCB50/Wo/jJ979WilVVsx+jGWhc43mCZ6YKPAMPwYA/suYhmDU
RC9Br9RuUQqFPZVw3Vhf3PK81+lVLADfBFB1SyP+ESmwulBQYcPcYXQDwNWo2hRA
k3jC1Sj37NrxgFtd0TVa/gE2Z5yLez9VtZmwwrW45aMTjaNbmHVbUfjLHjRkZuvs
ZTTP7R9E975Z2YMwqL9wOczoPTyyNA78Cho0ATSHTTsIj0dwsB4hVRNStk+2RF+P
agtEZPzwcuJj9BM7Jm+hSmzbN5vgoi9CRuzuDiv1/Pn+B2KsLsB7APtiNhEKvlzd
mJh8EuLSqvk63a4UfcEOQSH8u5fHEtljcjgQU8mQhFxbMG934o3Dhg5kKHLsMr+m
bpSHU5INLHUN+MXewD2l8M6o9Za03/o+l3gbyyXtIj/Paz/Qs26O7OWy7nzGwPTz
T8OX00bbb8/llZrJRsJCDhuqSi48oIH4l6tWi6W9hsCc0JJrj15o2FxWl3bU0GTi
bxp503VomNeUBnGWy6MYQ6dUQvjjcxK2dMAv6KTkzGiWHLfJ4eR6ZyGQvT5i+lbI
3zsMggHDteiVmTS0AXPsXSqNPbocmOMlQ1s6ZBUmg7zp4KJ97Xm3nD+I3+KweAPx
uXDY1xK9jP3h4gXJzW1whqOuF58IMoUKgbtHzR46tr6JGo7lGPzwz1wUzNWeq9CZ
SCMV/uq4+YamvlSRYxwL3ULJjx3I3Hpy0o+2L0BJGS8h82NqyFqn3ojulg3lmhyq
gFmbxHMcPlK+X1OO9SPgHRWFVrwyIgXukGz3xbibzxMYFBRQA+PUS0w6OJZcIiEJ
HMO51enNr+kzrAbYi/KtZil6qZ5s6gZR/NIMkxW/VF27afZNZ8VQ0di5bkw1U+gh
O3HJBhrhzJ3TDMwKkO8bbkrsZQ2qe+UTF6JkUgt+x6wtMxkYGYF2zXlO7gk+oe71
rmPrW9G0MemVf5kmVwbgHA3u/qDMHxG23CZPHzi7nIjIGTqZK/ciB949n98Jypgv
Mh9Gan+PJXIGMD0UV+2JUWusZRlbe7p7iM78C+nCyso+mQ20APDaE8HUdKw+uU7V
exT21GPjSaRDTswe533FTjykOLt6pEGEeWAety6X18nZ2qqUDOtBFK05ggf1HBNH
3Yxs30bWfz9Fb4WEH9EabXd/k+ZpAdK/xQjfWLd1GxnPcN+S4DXVUSJi0ExlEW4I
mOke8y3dcbiLNsPhlAfYYs8cryFMxB0DZHYE3uSqYhCjTpgMANJoyjiKBVCOJrZ6
Xfj5JSqPm9/FXMk0e8RmYSrNEhJObV3tF7q7KIYqnO5YL/vGMZhui7jYqtdoXGx7
URj5DfXpgPrVSWu93NF1ERW8NxQmwU3qqC4OnReyLCaZHQBEe7m0/smcjeOMfUO9
SM+jclsvfgd6hkop/oAoNnjGE5UmfXHa0qkjFZGSEnRsyyTtaBBj/YwPKWA7wW2j
PW+ksCkhdVUJhJTVThEOVu3RGBOhVN4SlcWkcvEnjvxwnYJnBN7k2uXe+PKweE+J
yDiRoPDQkDhmSqfPAciLtLRtmW/1QUAjWJBQpV57JSn/SopFO/avDbNjHSMRWBb5
5Kt1StcxTEEOmROphIv6fgUactNrYWPDaztrrkDTjISTqYAINQaI5+Pbhns2mfh4
xP5XO26MeZVvXw89XFxavhnOQyP87Ujl3c0lBbkI9339507B+s406mLbw43Zy5U7
gDHbP/slCsaF5T3TwImaiieBs0bLCUMhAHVZK1InOX4b7aUjHL3vacWKljjeUnKH
6rutxxHdmcVbzPuLAbDfcQEp7iD2MS7o3okROTc2iSWRre934xwsI3JSelU0K6vL
vkEyYc4ERw5ddxIXchi1fPdrDoHs2bj124LPLNPxXL6j2nZTvyvu/p3Tmcm/e/rg
kmE+uXmRuFtcXUL3C5qBVbUURjRUFq99lx4IEV4a9FhLJnbCFZNll+TK7VWkPQwO
osx5hXijGx3TwKhEusRT3w==
`protect end_protected