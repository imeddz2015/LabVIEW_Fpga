`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 16304 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/9huKRhRMtvnNqb3Z+UU7TahEoHV+T8U3P3ufru7l1O
3DlgtZzb9QxCbOjthp9+wDkjygH0eUfDrEl1ovhZG631Oq2L3PXfuycKED6mt0PQ
ewh5AQgcR+Pel9EawLeVhs+7TN4E2NdLSs5nyOonF7p0zBQCnKbTvgEdcvYBOWpz
+gVdm+nlA73iahqWro3L4rVSGSCHEGYAApuysJaIpFS/ryhCzu5kVKn/s6d8YUIn
4VMfM+yHY38cZYoD0qt+WT10WrnZRVhEUWLI2VRKdrvC4s2NH3giIoZigIuInC36
qMT/GVnzrBV0fgBzzMOGFiIDsDtzrNpPPUuwpPkHYwwRe1QHiJjYs12Hbm3WA5vz
qD5mto6YJe1vEWq7+Z3KtV4Il4+dlaQl74jZ1NtV7ks8KCHk/3YYJtAwHmeHMj7R
SuVPP/zVS1qoSSDdTcE/CLX1w7nmq4ueGDYEdeYsIx5Pl29NHFOYpglA4pOpGJz1
WDtya0ptMyJ7Lo9Skrm9yZOgdWVp2wkhl42aJ1VtKMArjs1nDDe7OzY2v00acYXx
ktDZIdHXqOLWNHJe+0gukXUg6UXIm0WyegPjIIgNNIFspmXW6BUmb26YmwbDZvVU
dgq9oNmCqfXmwQfGpOAHH7Sri540MZKgqxOch95nNNDWEbypF4COXmDQRL2VUuFt
8W6ZL02gCPlWBLEyFsLc8VLWi8f0vllJg5oHGafuKV0aRJYCHnw1Gx4ZdPWaOb4u
BruniSqehrWWSAwqTxthj/ssAa7+/W+DZd+4m0MtogbjC6e6mzhUCVWD24OzuCT9
FN/TLaSa+CDAP4Gw92Lr0pkE6YxWcnTm1XqTK8y6LcQAeOOEBPha7gZAyv0qsMCm
CEHbzts/+Pj57BvScdT7dWF89FdJ8+dAZm+2JV4eR+JNCumI8Aa2uW2oxQX3QaCE
BX7aNUY5Tx/7XNKp5yMAhgVBYrotfOZYk+Rb3eCvxWhdJmsAMY+7QK9d9a+COkpd
AGr3YogSc4geFwJ7Xo5nECBc9EetSDtQZzx4ZuXktWw8X3B6/bI/UpAD1gfIiDfu
ifIXIdtGSG7EbJJsSimq/sG5UiW/6N8+MM0SzTs8u7wl+RRlOEpiZayz9ZpsbNxh
Y1YLq2PGzQkm2LU27eXag88MV6DLzjXwJMXbbQCMqMHMGyDiQMgWH3Nudo+t1+wn
ZyFrHGRVV8A8NPyWuscybqgDOONOc47TGgBq4qv/CrdtqcA4CA/wBREBU7WB9QMY
hoZy5oXrDGeLnejJqlHfZ/owHWoyP4/VD/Pwn/HcwprcR88hDVYxdvu49qsTGxx/
MaUyWBY6FYAH9drVlZzH5PmibkmD+3/Gdt62Ru5gsFKONanjNHF5eSqZsV1T/4s+
soxbfsBFbgwfUL5B/x0wKFT4CbxfyxS5YgEkVapEolF0MKccSXH8qH3cquOfNqxC
XzpFoViA+3IZiyo7vxvCSnpJYan0t/Y2JDPrSJ1gE9FqrbeXfWLnyRGzWFHXz1Hj
Xyha4r4pyLOVy6DW/O82imkLgjniXXEHgRsGzdJ9+b7Wag/YGND04vEyappUWHTj
jz9NZTSF2fhStUbnmuR8bfH6/G202jNQIZ031u+rkke/iMI/KPRu12HxDw7OcwRq
AtOhSCtXjiEGt+b7b6lFdw9KcnONx6D4fQNPGEDM4mypJ9mrD4coR803Zi4mgKPQ
2jdGtFSOaFkR7/F4X1jruVgycq4FNsewsHyMS9Umu1gTfRZO7oP4NVcZvbyL0sGp
nvvk5WndHMJebEguq5J+TKfp3POTIbLUxsTmVsawgJ1lXpYDhnoA5PNKlLtJWc/C
b9s9Yl7iL2LTK5hSCGlxt2P7MFSP9h453HDQg1vsLxz5P4/DTmovNC0VBX5OX6hI
ks9vbE8CC4F6pmPIIbT+FMCYpDrPX1vqTnh/8+gpz44rF804x8CCy3FeW+TJRxsH
QauQyE/pF1RnqEXGUpcscB9Lh+xzafwFkorBdgGyryOjEJJh4hZq4fY8xXVcGrbq
lQUleK7u29WY63ITUcoOLC4kgSB6ZyRQ5aIfZnGU56HQtOBOMo2QudYOzM56MVvR
Wrw7i6GofQ/gYgOPfFzH2fovvSnnOTbu+ig1bYEAtmYM0uUp87ZnESIFhVv0OnSI
ie9ee8gZbmTMgJeOfoBz5prQwFQI3EzGR/U11rxV6o1HNHu3Y8YzWb3vFfdFuGuf
ezEHb37JecYti7Nb+7uoEsGwnN3yGVrEL+u5rcCrRi2oiYHJxequcMBDsTAdn+iQ
XxeSPOe1+lYtJ5XyY0RLCXITU1CEYIJEvbryhuApKVBaq9XzhJVgknwFU2CbV+jE
WAhgwz2oJ3AjgZQj+s+Kvgf9vctZIkb4n+dr3kRiMaffTXT8S4ZtNai6WDuMJ/iK
EWMaKv+DqlTEQF/VPh40kqn5kONZnmqvmmxyHBajjnQrVuCbljrVdc1P6WD2zy4X
Pw9mkiz9AbOpOQonens0Sy0L978sP8em3JvVM1Gbn/PsD2ABN0PhtZ5LFvMYx8V2
m95MPtxS7JbkxvFbWWMttwEs8qMeTw1rEqYrOE2XUON4J83z2ajHttGKHNyafSv2
9F7wNYjHDOUba9yVRpke1ODblq38vRrIRzZxSnOJYkXYEqYBKsV55kZheI3TnCoa
2TGX885rUnSHKTli3gn4xdnfIW6v8u28NxX/Ka7xB1ZthyAFQDQDnw/Hv72P4WJg
ALeIr43DM/ifZOR3lRbn5Y0pwukfcKSoxeBWEHuqiMAqXXrfKW50NgdiN+FsH/te
H5btbXsqQx2tvdvWCfN14JfatgEMm0KUDdXwGlFVVV+nO3Oo/J0Hus4Y2Qxem8Hs
F6+I0345kqnEJateTsrUSfV21ePR0ywYQ+ZzINGtfWfhhsdJk+am1o+gyiMdH4CS
czozyTP6SFg6EYYAzOK1oKMPj9LWYnPb+J81IXTeXUTK9xz/LxQqlqfyuPGjzvAb
QgT3LCLF+TzWfyzwy1SIos+w+pQk/bsdXe8MBvHo8XLin4nAYRtrvpO/a9X/y1f9
0IbcWe3Lmw5ID+cM3cSuzFJgPo+zh8zsqxa4gDmJ2E+96/5Qka/HhISFDtMWLb9u
j0DBYgDxEWge+b6/lA+ycpPY6/E9AfIPKcviujJjyVV8WxXrdhpe45CpYu+QWoXW
wE0TUbuJsh9Kn41vxKVxyA+hii4ECbycsGN5USO30z9QvACPxFMyB0IFQANgNZH1
9bPV8cpHqN4MNx6Ygso/FoHLScOFoQHQ+PHIPRfal8BTpsqnRVrOe8z1Az6p0J8Z
sdRzCkFI7d9bsry8cnvhhoBhZL/1HBEEmpSdDrCycxrPbrTqJ7Gr64sDwpVgd7Jf
2ahiVo6sHQK2XKC+PhO8dVbK5ez5CQTtTORED0r6D+sty7rZJ+HrWaY+VfHmGw4r
GTS6kK2ezLopajLDgvYa91BWNe09ib1RVSUHCq4Y/KsWBxlTK3qgADAYTzDuq7KP
ft5YuoB5R7MH55f9iLmiVysztSd2GMjxZgpQKnI4fvuhJLNQ/p0w5c1s9fM/hUHx
QO2Yr8l5Rvm4AVqxSr4I14iOPW7O2TXBcWKthNF1DLzb4SwDskvaCSc+l9dzPD+v
LSWzAYU76D9pqd6tswv5+kNlV8ScLrLECh4rwES17kNQwDn9rJrerJPxAImVMXPi
g/AUyL2AYw3NNzN9NrbRlEiYZMjg8zcgPLjFVW2+x3Vv/Q9l8tqvol7h5t010H5x
e0ZfVJ/u/C/PvlwEDa7t4KpjttczoelrsY7VIKAcAZFu+z+XYVrinRB8871zx3sV
yPjsdR1DKJf49FQGz9PG28dn96LT3g45nVMDzY/FVpeO0b6oUPeOB526D45uCcBV
J5EDySyc/sEJCtja1Yil8OO6vKlB4zZ3GNtIXCq03iAjc6kR1lPON6S7bk8hO+V3
ONQz4vvwiYbE2RCvMCgpSi9ybEk0L1KOfxO7brRnnS+4XMI3wg0jf+JmuSWi8kDx
gefvzysWIn0dA7eCRsc4K5boyQrZz8dq0qnzL/7x5T+5ATd9LHeooeHBhRJ8tuu4
odYTT2D1ncF7kIX+HcB9Wf7feiaMg5WbFm/kdponGLIkS1SOQF0SLkRLyxRqpfTB
rL45wgkGW7bozgtJbUpeuJfPvU+aPZcSq+xiiAOQs6pn2kAtZsA6SMq8bLiDrz1t
uPnOeUQUiD0DXnB1dm/PJ0e+lk92KjP3DOFzkpVWhaDVdYkGepVCGwenUPo71FbD
F4mFrkuwfF101S6B63ACfKzT3+tAUx4bGrWAiTa7+buKDLUmcM3j2BqU9rQjLDvB
osPlVYtJco6fVzQCwSj9aBj/V+ux++tfhLqQN/Rpay+dDk+casAgL1KjbVUuIUCk
1a1Bb6JqO3I1R87ONS2eiaBbhhyqEGsk+2Tmd1B1pR9NRy/7kViXJk0vMAU8DiZk
QCYQ9mdqu1F5yYty1fpBt+3BI6tM27AniXLPc5Hz/wfedwjaSqbQgCdOsXcMBSTv
GrAsff9H5dra/ASbL2k/uI6UIf8RL9T+EwkBUvkMjOXRwH0mrecOObJLQ9xyGrA9
sPuueoX0ueYxegRRuqQh0HchgyrmgisHJ6Q9Xqxjpz3PlSf36BgR2JK+N1ojIk3v
Q0YhIguCS/Bi7rSfiHWAI3H//Y6JT+y1LUhRpaXcVQsXNFIS39jwJgEYxmP4OXEH
U8SL4Fb16zAq0oZvPvHeYGdr5E+8I7svr+ImU/FbfMMuKxugC79EG6ssxnZ6LNPL
OERlihZfLeTpkjnPnqpf1GO/NN8XFovpTWvG0FZK6vsYGbbWpiPuHrLCrZ/7SCYz
3kun90ZduId7/aU/XDO0U2VnLHrchaWeDR6BDQr35ciBy2Fz4MLubYHrID2bAWEX
+hx9EwPC8l/Qk9JBigVR76ObpkHwK+T/8xc0vxMwmDBwzkzcPHMKUbfy0KqWIeaI
6Ppl1PVXa/HPZLNAlQFp9FY+KdeRAZjsEH4wU0ReJPONVzZy7TlLGHnfUXoAknFR
IHO4kJ7HYcaYNdcFhRTDO4naKqdq31DVgPWSBqrgZVKOPAgsbz0ddE3lq6scUOty
CRiIyyA8mYnfTiNKfkEgF1eoe/soDFbKA0kxQWB+8kh16kRui1EfcAL8XYaps53v
bP/pZEGhqkKnWU9/4n0It/frOyMVI0e1d/6lXGbIwnEXvibHXafbnSILjc2+z6Ji
KpCCu+QVbTzwUN/SQM90e/MUlUR4eAraY+yjQYCzc8Si5lFjOmrledwPFXcgvQEG
ehxTqxI7ptWTvVjBjUfhmoWlJ6qSVkag80ts30wAap94RtJe94LipNWqtUHP1PoO
YDehBHb2pMJ3RxtTphBTgVPq3t1Gdr6TF4bFnLUPnetX5uxrn49+b7YtXz+dLDMJ
JqKDMDNU+bZeZ87nZRGiB0G8Mnx9KpiXRX621A6h/QlMaGVv9eQiMsAog7Iqc1i1
2j5bZ1XgGMJYs6r5G9QHD/jryKBIU0GlsjN5CWsNUTZA3eTwj1wOMtHljZBknf+P
H6TkbSsTAqcSRfVFNO7qTdA0JnSlbOtvargiVN/0k90pFY83VS9vH1uqQWDNmwnb
pFAYmoLlufPOhQCOtDgnAezP3unfY6O0ctYOyg4Oo4frOxMuuUrrbcW3k3c6vGd2
yNia5O54zkh533wQJ6vD9o26CWJWH2HFmijQy3m3AZklFxY+BcMdmygLHJuoNy6P
AK7HQY/6xcoNoC3pxn0abte+4o4IhzJorDAvbtO5K3yj/9/m//ARQPU634oA2pdV
H1/zBbL6DMOWcjOGoQEmDUjNQRcQRdppYrSHQettGlqBsu9INopxdt66vhtNT1if
tpn+dJBbdbQLcOrIHmLT7NCF962p4/Qb0OpgFWoEEi4IPVzHv96sJHJ9/tOQ4hI8
NLqeQoEayVcuVomXepBXRPapi7b764dlyX63MHcKIhu9NzYj6HgccI63Dbt3ChC0
gSTKgNhgBdXkQgqVJmSTDJ4ODNuqf1RMZpa+VrpXYAw00LE8jk8+ZHakdor6SRWe
2sSjuD+Ahsrkp44KIULIPZgZ+JloRhvtNhJg2mk1jIJSy37M8LToUk3flQGF4TUh
CBVlJGo5Vx/V58krLUyNUuX+MvCYPU/Ek4N0c2N2R39crN8rQxglzKg6gGqSBg/f
Y7H9nIJOPcUZM5sOezb/Rd+Mr4EetwRwtkM3fscTIMzMCkl/mf3sK3cJJOSaZlTc
Mti7FYCy1ssne3j5Bh4Etdl26Zh1MY+IrXyDYMG9s0/uFNcR5ne34Kvd+42j4Pk6
Vnj1RkdfoB75EBk3TWuhoiCwT5NeHLO6txy+UoPMZZryJrg2AtVxFm7JONEsVOyG
sZqr7JNO6Ra/UZef6Ye3h6/gP95BzCRW98jsw7Nup+39pqOGkwlBx4F3jrGN3tZd
aB8LPjzBMC+tx3/jH93mDGCBy3TsycAh+1Z6TKHkg7KTg+bFS0jbhKTz6yQBmMmO
u6EWhFDSAdcydxY4bYiXXtxDPRfYvmbA/S2+/tZYUXxvu9WeXQOI0voUHaV10F2j
7pU9Z74OoedqzIGw9TKFXg6UTkLgPRYSSLj6bbCRV9frwbmVwriwOypPgAX0z4Vn
e6vIBqIyaSaJRZcFaNY5wABLYfKK8jm4oxnQAsCFZty1NXMseeaunxjboQVQXwCA
4IJWmi0VxFCUWjFhWAqSbV72aTehffrIlyUHXw3GjwwEIFuNDSLHiR7UAEsLQIc2
1GdlbxhiHWSqk37j9ksiZe4tz+y+/eT11OEC5V14HsoqL4z9kjoCcphbEQQ7Q/H2
nvwXA7Zmo+eHRiTDv5wnhdIzGotQV6uw2VF1rViUcNobYvuVYwk+8/BmzBaHt1Mx
V5glOxlli0khJj7+ZrxVYMT4yJmcPIRlGxcpSDI/vKaaU9Qulq+6iuHYcCf9f5p1
ZdrqFZ1KeVrcCLsOZt4QRBY1kTowJjy2R3bbLqzvMvPnguzKLNgzuXplGoegT2wE
qO0f/2/5dVBjHDIdlHH85ZjgE1oGHYgBUP9ms6z2rg63coiRS2CB3DEzf50l8UTn
yYM15RXQLv+3kZJXXwiYlRANyQuZDufZmQBxsh/JFFJjq6U01L2dPClgx492WxX4
I5Kd5MLcl4J15yfAzorF9QmsL3TxLvtEyTVN+ZKr9H3UhYVOWgpNT0FjOZCgVcqI
Shf+hfuZzwQVy7h+7OzlavhsSNthn9zzUen31nDBsyIZPRXhiZ1s4G+EJr1fpQgt
PngaTlIxTmulhz9WgmdBh4RILw2LHYVpM3jrRGeONt0qe3X6Zqku15A6PE8WA1GR
xzYFSzvdnJUMf7Ekbo3Dklqrgj64ndlqNPI89fM3MovUiotAe12GNYPy5clsXr/n
dqo7wMsdb2hhjUhFGiluiCvIq3qvsHjY+vmpmX7Pwnn9AXaKLVM1l0aEt6/2yOwS
QumO5yKl9Zs5TQsUjqP7gi6GZXAet1PXTDDvLNLz4oNsf6XrcuGcFlAzqmteNQK5
N0dJrqOO8VeWzUQYfP22/Wj8ZshhY2Ci04+XEn3/tmbenRSVzpzqVPjfS+sdf3e2
4kjknKNnYzFvkhwkors9WwvGLvF8WDFQmKaxcC8KVNi1Tmlw+7fJG3fKmcGmGCiP
zglD8GJPZexaijGg92/jRlj1Qu2AsyPO3hv26kCNaLY0AMCAQAvYOGim9QRa9ind
tQmYFxRlpvLFSGlKlyaPS0K5cR6ojMIRJYKyTp63EQpGPy/s5D+JSzPK/GhGm71O
WdLjyT5JdLkzM22eRdeBl/AmhQYuU0Ot4KI1J7pKULv2TG5VG7fR6NKVp/CMh7V3
wRVOPY7Q+0+RfUxNMfZqDRzyfLFVWtSty7L8ZsmWLHJIdTJap111msQsrEbOvv5g
inw5vHyLvy2CJJ/8RFMLw2sTZJ+jpQX0GfkGcTiMv3fwti+8ofdaoPuH2O2lpk0e
x+EBLX/J8Icr1AeE2DeWSK5Pe5O8xTLAmXJOeaD+jZ11cP2t52g3ehVLU0Q1ibxW
44oS6lwMoZ7z4U7klQY16p843gPzBw1f7QV03zfePkiAqC4lvB4iDs/l7wYk4bfS
SSw89v7UqYF8gbKyTC2hTYyt6DVFcILlrpdcTuKZIIZx26+H+vmH3aCi8yXnsbsS
gdCZABWM5bzeTOW2K5CRaQ1+pmJ7rQKL8hCGeAQaiaRBws8LignQJ/Oy1us3iG9c
0WVFFE3xKQ2U8ctdgLxa4kjcz6ywmV4FgUDUeiCDjEdk1ebZTGBP9xAfYi6/k/ot
Fri+IWinoaMSsG7vbZ/K8qYc0fXshv6RN+YSlFO4knnD/eemhTzCL+EXgEsiTMoV
/avU4vjZBeIJGfuAPu1jGrUipA9Ffqol0fQiD/SwdWHrJX7sOQZ1+4LDajNW83CW
djlkBOGR2d1K2iV9BhNcU3oIlf7YcGPZWd3kJA+nvv5+0MetVjoOJ0dDla54tQ6f
e7CjqjGW+wzHPohBT0EtW9TxqhPf0GhfGe8nXSGwP9Qwl2lW2dKptf/434VOM4Wn
gMd9ygJK0onvP6nIWSLXAWvIMxB7kst708FU45YG7Tto1+/WHKRSlMCKXEp/taRI
QPIMDfs8nA6dKCtaHQ6D1/VrpuQU4bz0/jEV9xh/oXpGBgKCLPE7O8XlfRXxaAD3
q9EkqENSoQRiLDZRgZEI89hVNlgTVVKUtlZr5OIBLzaVutBL4Fk34vYMWJX0atoE
EQOXIkOeN9LGwoO77JDzR6pFztYha1YkkTZTRp6rqDMXeBsmKg7J9iCPGVE95XlQ
1me1o2UwyB5GK3j81gnWqJSV2xmK6ptBuqHkqWjrM9LHtpAR+s2eLtzm02AKYpi0
x+EKTGDCxu7wn3bqp81QdGnEFd/o3BjUoHDNFM8e2WWIEf7azxCI1j9J+nEXzv7C
CIM9TWfoWGhHe+zWVJDJuMYuXBjIk6Ot57pSDQIpXNriT/bl7FHZhgXCnO99lrpF
CsmRyRM45GSRiLHzRNDwDnFb332SmIfesrW6AWxlKSKOr89qDr+pYwyRX2aO4145
So82rwzoV+s4J4NEJLbZG0z7Y7R3N2+WwZHjRg0sv9uDGEfyjbVzUmsYxkEOH5tY
6Xb1Qpf/C+XrtKTQLTx9eSM9g1NxrPDsH8SzpCcjOSCobAYAXEIYbwdfds5gJiZO
mUerT+rh+MC6F1g8j9t8HWyruSG138a+GdiT+yq8PR5G2N/jUpWisHBCODw2BjG3
DOqbiCKYq7NSEowFJh5u4M/Aj91E94AjyxbUYNjRr/bgBtOVIQYgCcURfrhZy6mZ
/xRXTCZsJbp3Cf7YOqfaQcOVsVsVCtcXWIbpXkv0Wp8GJYoahbEjuNho1GBm26cl
Vs3r66+8QFsefSx/N+K9i52++QT/RqyIejtZEhb5XxnsfGbg0AY8lZiqtaQszKHW
rRdt84gfoh/YkkOJgLDcbel6XlTffHOXJpdM3rkftGHVOcpxP/8MwKNtocAKHBR7
JsSW2fjpe5xuzF6TFbJWXnFzlR63NniZxwZgXnGamvPfVYO0XRjBcZ0mauEX6dmQ
qf3LHENnaq9iKHItZM9FsT4IRthg7mIpLLBnv2dvoqXUPsawAQI7POnu8vEoDHgD
gpRn7buobLA/e7t+mZXwoS4A5Eb+WHpnN8F+qizbj5E+Rkv3uGJKJT6ZeIqhm4q6
sNUdeIo3s0bvgWBIoxDtfMYju2EbplxEwVO6bztzYps2k6MbsOEuhD8/Xx/F4l4g
ZAdQpYwwvw8NcEnhfnU4nb/I1IsEvcgFB4gxcSMIU67fUQgUwaj1CUkoesv60Ggb
sWhZ1cP/iAIsGYthZTq6OifvUM9jDJH7JQSKUoiKMfZ3u92RTESBUrjwPsFoRI01
wK8bgJbn0A3PVZmPT6isFcDoSoDHvHmqra7Wb2rCG4NkDfAqa6GGO5CVfWubrUyb
8gxpP2cxYJnimJGLRkCzlU85foSoGAf9e1ly+iGi43fMrXnfjONAa9ZDP2Dg1Mrk
P377xcvtYm4OkvtpAOlKU4RvIZpOgCYIuyHjE+hiCqanHNpT8WgK4Y7N/7I+mI95
Ab00ahCFYkwXLWNPx4UR0/tt33QXptv79sFVq3OlhuK8vMTH+4zd0lMq7Vgais8E
AnROYJ3dRs2SyfnlFya/CR3KiMSbTuBtXBfgybbwstnLLuhNlxXQgyKwcFFx3BN2
IobQqzuGHKzA7wVfpE6m80PG2zvckWYMF7swMdFUlr1aDRXNweUICGK8DwAwC2pa
5LIUkABCPAo3vOR6OB5u0d/p1kVXuyuTQSVw3Ed72VgckoFJmggiAHj5uAL6xsdL
lpnm9gkipnQw6oaNz9CHB1buu6X3JjgpQ0+7UzZbOIGb1FOMmM28ndZ2b7TxhJ40
6me2GH/AnHa7cbd/0aEKkEIzev7P303U4M3MM2NLDN8jZw33Nu9VdZbh2IpqwdIV
xP3OFRWDvkhdcKGjIrgs9e/3PLQGv1Ri7WjPzzycKDTS1aZ0UR7vAIuXE5gIH5IQ
yt3njKt4nyk3fWaVS4CIcfODjzJ4gDH6a4sHI1irW8ddJhFzdqfjLKLiHGb2Z3vy
25GmdHyxiijN0I5CMFAal3i2DMk1WLU+j2JPfexyEBf96zLriYIJJkI+3bxpVMMw
2YX+OlysgZiPN2jYPTZx492WS5dFmSB6cyxs4R/mUp2bO+Z85lxvBBsvqwgjsxA0
XIazCq/gHlWCuCOamtjTxSGO3cjdoiXuBn99Eo/r66cgtDBBY/GiPl1DBkPalpxt
EHvYsAGVsUWoshQezGjF/5ovLl9YzrR3fjENNsCzTyarl3R1I7C62nJWDfdQIfAW
rp4ae++4k+87QYzmF2ZkjdDaiNSN6sNVx3MG0XqwC6lPAptwVZN8raYGRqs+5RyK
CpQmF+hihX/fVz8+gAKrYVVdo7ABvQPsFvXaKiBfasu5FayTpFm0WMnEvv1sJlan
XWfWbJtzG8KlaHXZ6BJei5abyQV/MLkBHbuepC/Zl8KCgJM8IE5BJRdxNheasoN+
a6Lr1tdFq2HUWBTeYsTRlaG+OBCdetk0w8mvK/4Y9IwB1wA5M+MtXgSyquDbB7gd
2J9P4Y2kuwbwzpA1rIOTht/ZANLueAktov+xliOd7pXJcnxlDOQ3oEY8S8k0zKCF
TO4UYJd78NOw2+95kfzcpkkdIFqgNvv9z2rNDBYR6BY+4+Yhvl0ZMIrUfOeEOxX4
1CfJjL/7MC0lPHMIFxnLmcjW1rEpkHY3LNbHTGcE0J3Kcv4bhJVWabzM6zppRrNt
ie5xSf+Kb4N6h3gU2nMFkDGqSZCiva6sTal4Ae0HGbgWKLJs05NY5onyr5wBbqWk
BCsqDuysDX6iE2tt1sTAuuQI40f94Bb3w4Bk8aqg6iFY2f1yV5a3P64yglpbrLLL
QYmlWfZ2kpleQ027nvb4foxQ7m1eNyEfZHOUXBh1m2ZMb1L4e84NgNhecgtHkyIf
eMhmJlIlY/KbrcJdYdLue2h0E1H5AAQk48C7KcvaRtNp6KS++aPIteILnznHCA8n
JEwMUZ29BIYFpoUljwqJs67LXZ8EaJloirJB58KZkjkNjrVGtWLA2UACqWaR/FDW
a5UU3UwgSWb2G32Uqohm2RdTAM2TZW1nxEXsuJeKgyiUPnZbrngfDjtroDKF8ToR
2qcHveXPWrMAzQ+fYqR8pwI7+Nk34QRwO3QziP9i69kEU3ggf5e6npCfDtIbI9Z9
c7YuL3ZvM4NOt5rmvvpDa/cBGqq6XjnI5mtlvwbanOVb0KlAMl0SQwcDA48tmvYF
ecdwzRbwV0IY2Ph0/0uZ3NU26lcOnjA7PKKUQtuM1ld0rwvQG3b5RIwU+eSMWMMS
xPmbcOEJ2Deg2AYOiE+1B5OGEHZ5pmixVyiCg38wFLzs8/JwAFL/As1vSLZjPvvk
w7vA8+rRkJHdcsY3T51+wDxfIxKKsiAMdaCzUPFoM2PaYQ10EmKDHFOxW5w97zMx
T3+1cadGhexyZ7s9I+6GYJdmYNh6kir5ub/uwOonBQPx7BHmf136yh8iTxveCAaE
pJ9gKLJR5kFSpF7zPykWJrTKJero4xyApFBngci71UoXA2ct/cdi+Rkz28oUL7Sa
p53XcUl0kbh/7FdsDE+6yBa6dFvb9lXPdNK9k4cMXiv3ORvf3LF8tdvb1HgUnJ9H
eRvgs6KbSPhoFCnQcRkrMTIPxKWmNBBNDCqT6jvwlpAh0lEuxU0ectYp6tqSqa7E
h4jcwUBkYAq+Xf6zN7Sgjj/h0lBY58CJEHVnwPG7AWQ3eNf4VrFQkZtS2E1lnp7D
n46hB2nPlvEUGw9Sd9rnS2zEBgpn/oNW1GvNDqnN08snhsjyDAAXa7yOD0Glu7PG
i2cBBNbnKw7DYsx9f6gHpYXg+vjy7U/dSDAvWO3ifvIUL002JPLdANJZjIHDtOT8
RWThQHSxZE8YO6LgPj5jZ7UFAc1EPqGQ2KQExOD3H/QRK3QLzdfZ0mnuHKKVy0tp
ktddMziZLGaYT5nwIyOOZ2QohVTCDmmAfSdPSdTCXgkEbBihBAiE6moDVo09Elr+
XkYA93WDKt30JqpW+6Z/gf9Gbv6Walx/rsOVW/umq28SfeehW7ylve9phhDqtm9Z
ZbmqfTIHYd/mExcW07bpqCmLu4dM/Y4hcpD7OROLepk7qsSIPCOuAXk0pPqa0gkv
/SR2knE/KvEG2Npvg+symmN/UpFCQiL/h32E5kPkV2TWQrCjYBBmbUNCVrObISOe
Qz4x4HGHAfa4w6ey2WSBhlecw0bO7CpPmugttGj7AjmmblINasS9ZJVm9rUKb8w1
XmjQrzx3Dc7FatJgg2yG1J1A1zNhafjt4S0P0FNmabMjZ4J5dBQiB7+BJmk8KjzN
ofSwwTdsJA1nZz7chfHlMmrKh4vPw8HhTZb5zvzGOGdqEvzdJZmdWUw+l3JhZZUk
bv046onHMGhDf49M6F0mS3B06yZVvoONA2MhLdW1s3J7KigaWtIuLsxxDKzIgCHT
o6lMqdN998h/kAHn1+d2PVKxkRdgCxjZKNf00QlM2Wusni9hZ5I8eyhYUdxYlrM6
c/M3gJp/WMp83V2VJ5/Dnobtph/vLftIWNG1RglihkgpTyM6mUWXhcq+6nXULj9m
G7yy1KtsmLMq6DrW7YjkVvyPHxl1cBDaDlOwroaRCIcJLu0GeMyNyGIhF+QZ97Sz
Ktk6fxvUlAqEZyNCNtCdcLMOKj3t7kJ1g/6Zly0X+K7o21MoI2Vqs9mvsElcs2Xv
4RslQuRZerU0grU219G5mxhzLy62wZE4okSDYO+C+3g+BPkDrSu+R+a6k0BQEejm
W5eDV9tjAU0DwKJw15f/bpuKG8+5fjNkzTYTNV/anOg81fX2fvlnIVkxNX55yIYh
+kwegjo2nhSIgZE8HzfGLGeh13bIH50Vjnn5DxQGcZOWKejhguod/IYR11w/ROiw
mW89CuZrzgYWFiXrT+n5fmK7VO0F3JaEy9DJu8glp1cXuj3tPZ0Gj6GfSAyXPc9j
67fVKyk2uHvxISa9NS0eH4KqdkyxPHM/KNcvO7IFjcNqZZ7HT6Mv6SMlkXrutHBG
ho2nlhcLlxOcvCQgUraZFXOwA2gMUZFPeMM/H/e85lciMLmxirx+xr2X0kU9c192
8N62KaP87fmpsGxX3M2mc73mqgYHAMQtmxjGu/UqWHSdd8TTkbzq9tkXTQv9eI2e
ord0uBo9KfSwcP5Av4+2txywaLnB2L0nZC8O03cYz/Mv7zs81pJUZvU/PoomqCWe
/MnDB5lgyrG/2Nx4r9WoJS143rCu+/EoixNYL5oDUUbmUODt0PhfzL6lngtufLoK
5eBteh0xlxinwnVccTUiJHcGyZHNAcC/JpK2XLIfRuTxF7dfiB5k4nrjen7+/dW5
ydhplicTrjNS3rXQZiSaTPUy1h3y4AZCx5gMHV2y5xsX54VZBfgbBca6bo0ErAC6
Ltd9KPaOc6hrUKugmK18mQwLXrh/Dzp5kSFk0KrrwXJ3lTILn3jLrmmK35lO+9Rk
JV1qPOGFAOVUkm6af2TSRdIbaG5n/gZAWmFNAaobtAR+77fboyzTSOTFTygLVFFh
t9Q5B/1kuDATgTN7MEmXLAX1zBj2/l1hsIfGB+p8tauUWGvJxkWMzNAQVOc0ITDX
reoC5RTgZR7gaMWuRETVVvjn2VIwM+f0Vcll4jX+EeCjl9nM20HdSesLtv7XaAMa
0zAr+e56J4fi17PXlWlsIyCW21wVnA8agIWQeukDApDXBjaPvFSstmz9EQUIzZYo
DUXzRSETzc8sQTxlm3lFK7WKy5IpZxZepfUcGiHL3ozB8CKbiYN+pZDEPUeQwNwX
s+YQCSangA6XtRwoTa+KIIFuSKBOjVbPsrbVmA9ltIW0KHSYym3tHq/JXY2MF8ys
GaphfrD3USL8tqdVb3n8ozyRfQIoXMnzcNmuRsRnelDusjiBMKiLnz/U6KZqtEPu
l0066KnEWTj4UNffoxaEOWol284IAElgqIgbw01vK4WnFVrov/Y25vXL+FY5kvzh
Iuteu1T1lAdlUJR5cuU2Bzk7n8yDQRRuS56YCJ9i5kgn06ZBmnIxAREa+zK7z9+e
6M9Ko4a/hKTrYRMs4wqTISMaFjBzG263D72Nn/0rkqKS3s+82jz0fNAAZKOQ+/D9
sGLMADj08sIxMtcZ7jmuQoUeCBsu0YtPOSHj86cM1RuLNAgPVJtaEjisZI4ugFdb
PUEVBicrKZqiJRE/Gi+gicB5xH9uryKV9odRlGcUhCw3SbA4xKdRNiBD6cBiBPFH
iAP3aglBZqVbYYqAKw+bdr/0DfXw5us68opotyUGb0NWJEtkDqL4hMensHWmss91
XPi3yb0sm0OKG53xPPsphIImJSQx1p4R3SPjeBI9aI5K9VgAi72YVE59bBBO8o1q
XpX5RVyY+O0nRy/FA1+AyEGBDCLhxE/taffVbiyZm8L6WuEyDihLJKG31wLo3cBe
/ezPka0vAxr/C8QFcUTFY6bB1LpN0NzJtVc5ByGJMvFW1s18h8CV6gY9W7kjfegK
6j3lQWbi6L+/l8TBGnU5WSGT3bLV4MoUX6NbG1yDYHdkXFBTGVfdi98hNoldIwkM
B2+XgfoKCRPbwBrG6CgB6Kt56JzHeZTzzuaVU0fulx3qNIkJkYIAde1Y9uXza9RT
Z2w1TwdjSxTQyytVned2KAOwAeiW704HM8qC7Qdu39kHfBOPR2iq9VOnjb36hbFM
9YBvtbRqk7ZeeagKqap4kQ3y0aElNfXW4LnECDFsGr5p7fP1iyu+VH9ngcPSL0YR
CBjU7QOI0ENrP/o8PVnl71MOQ1ylWrIJuEoUGKH9d/oZb/nEYGNhZKbUfCb9Bft1
An6W5gQRHHu2usQyymAkHJMtzc97ze8NB8h93h/0NehuZEgEVlktPslIHnssfHdg
oTgK98P1veLEc+rtY+xK7SA+gE9wbrRlKrKY/vr7wK2T1G6jko/XoGHzdYTSCVXW
oea6IS3teHWEQiRNeQVx3eFOUSYgVYRPpPYdsEhWEtpSXCV4mw80f3jYN0NLMcgV
cczCWIR2klGQfeigyXMcQXV0S8wa2REV4HyCxf7XQMBpGvebb3p2EebM0oLkrGRL
ttBxxQbpHwOLoNMr5/VCcCGWnGxqiGjSVgSIvjbaPm3QGV2PlHPYY2eDTGSYshJ5
7ozlUBrL8WjGI4e06dX5zT2RYGrnAzacP/m47GZF6bjOQTtgqzTISfaWpXH/nEaN
3726yLnN2XDQ+MpuERV0ZlYl60LmV7Bzo24HDz3Ib3HOZJgOoY/Cwe17JqulhiRP
LyXh9ywT/4wVn8i2O4nQV7E7e8wByhKVfM3NZ/dveGJcL2bYjx1NFJE0pBuuTv2Z
R92eKJxcF44lXbHg3WcrLRPrb7WUeeLCuNK/WNjzjcTYMMfmbu+UYGB/rtjof0ow
4o87C1EcowORFQVodoxRyJW54nNkuQDeWwnELYfnhnDbkkCZ0QFwowMfiwXeCxp8
HBFonzba9x3Vv+HG2795JLTYnJqAa0zZimoSnw1TnpgzCtg+KZO2yygCNkzr1WQT
ImMy51PbH6TNypGUohfglZevKEOJrFxVlq2Ft2PRVZ+SaHH5p/wOgvHfdlEyFDih
eYhRFzhrqCUGvSCsJiq8yHgTNGd2aT2lFURH5UcLLh2HAHp8+MIKGOWnFaOkD66b
jOgHo+u3gt8pvtluM+5KVpnkZLUupJaJ3EY2Beni9cmWI3KgZ4dCOWrBRb5WHhMA
TfZ1dckYSy6qxoWiMw90Bw2IuC+CU0C751T08tKEg/xWvuDvCoqYkCAG6Ke3TiUV
0CMc9nag649U0e+AtH8EuDDotGyEAffTGlsRsNN2XON1VEQh/XGDnvOGYbFtppTY
vuLmaPAgYtxtDotW/NfncPxpRJPEebJ6ThcConOXw9i5gFZLTUvCzclJ2qV3zP81
gUjCZoyZHRsxNl1xU9YhqdUOEJR/W34rIb+26OQD/StsPQqJnUEgKNApd3kEc4OP
x/ew92dmYie1TtVvAVp3gYGEjb8LlCGXlqkzHaqnpaUQZZaY16XzAdhgS8heG7Hq
sVjCavybibTKR7Z3g8gZjOI4pHuvGwy8Ev34STiVKJG5QBK12Ic1W7JB4xvHvI7E
YjwmcZB7M7VNW5lUncCV/7lyewwaTXAWgFWsKoi1Rwq9En81+Z9Wl+fSP6G+7vdo
JOV63a1RWC5zfoitoF6x+XG9XBtqHsFxLsw6q8i9QGl/Il4zH19yMVqK60viMzFR
bWPlU/M5AyHCGZ8vjEEnUaeYiDQ9SuwdEoQhPIR34WfSX9mf94F8EwKZWF3ICAVl
sStF77Rer3ayarMZzi171DY8Qkj5JbLEywH2rnyRJJczPrACFsKYpubVLHgERONA
AZkf2910F3lPxm6szvS5yzdHdp+yGYb9ikROqRY2RKDJoFu6zTmmyaqzR3qMypP6
QbwGTG450FK/+S3QCBpVeh+cLl9ALmAn+Oyn3mjb4mqePk+YmOI760HC+W9Sl9Df
JSh6OiuxBSZK3J4PQGOqRxf6gwnvMXftsEgsboZ9xswMjk+qsEh1qi30qiRSYkJ7
d2tJ/OJEdo/LTMCS2WSMweAi031rkuOjiLyUAqr6YodN5eW9KFndgB7EojBQv8w8
9A/G2mQJeihiiIGhyQGOCMcD9zOihCLDr6xPcltc4c3qMdBcHh/pYu/QEX5SsmXT
hNJ1zdxxiuJuVXNelO1+fm45iwkQZWJqFdE7NMf1SlZreRD+p59fSAvb+OfVyldF
OEMslLqjaGLN5oOsHFNGY+NTXSnGMzymkhURfME4oO4SX69+STH/GM0/eFRuSEw8
xZBsNDgrw9QAIafhfqZ1UkFt64WTfGyOQe3bdzO//AVfm7FUaizQ6kmJUz+GATz0
heYHiigGArIXo6NERW3DDZ00wnMM4BKd5a7KbE2VPt86QaYL7+OG2bJQy7p9hC1A
GwCliJZtpeYOm/EVrBoVyi83rTUpkvzHPOAi3OabZeTRky63fjrWmcPcqHsTu8du
FkW/4f/a8vG83TIazHAcSxhqwdcxqk10NECD4e1xuNXvdNWKqFtSm3cvZhLPltRS
sepaOlBkn+xAW5NoaEAPsO1UDMkfD8rBeeNIhiUSh43dLcIcv31jZHIU4Fm/d1He
aY85C9TebyEYOYU4bvGxTFf5ieytqlYmRwtgmoHnJsLUSzu4/q9tIouh8lmb0VTz
f1ea+T6d8NPtdRskhdEuwE+4l5rPVHkGVFcK3t0TZPY7OvzKigoFMs95fsAcRIhn
TRHw9ZqBaBiN1cYVKlNE7n268dFligI8UcXJgCXHsAoq7aq6E4Qa8W8h6a/l+k2+
by/vk9mR8NH/8JnJBoZgH1SXid8sRnNs+BkjnR1wUduiWkFOn5ggUhCnDBCNR+xj
a02HMsXaPLvOt3G8qiavFrV7Oy8SOBnX4RDrxOWa7s2RqifAB9o3TBouQPDllU9A
Icob++hySW1qA/TBRfVTU9TGcZoOS7ZDuT2lIa6gmAIWnPlcdoAi3QuERB9e94IT
lDg19BUbdTzzeYN8waml8VfFDsBbAB0epxof0m97BbhG6TbiJ5yTSmo89Xj87qXI
6Q4N5qNRiDCp/uPI8lJHNPTj/jmyIgnvY63gsbqLcEFTzHVeRgLbaP6xSMQir3kj
oOiBUOG0Cy7NWu56YD0Ckz42dqya4DBBGRH0isczenPC9OHZeNWrgh5ah/SdOKnO
VoxP5XWHOlbVTy1fWar9VLQ8RWppsiYLIYvShsUZJwNuEaP8ayG1c9iZb1UhWZIB
N07rKCsa7woxEbr+ojs2P8oHm4ROCZhlxdeBExt5hf3nzhTENGpmVAwgas4DbJsP
uGntxmWegrNL4tGoxIrbnbF0xlyWvM4Umk2Ura7a7fTlowwZytbWRNjXOZxI3klp
KcfICU6nrlnx5KvCkQ24Bhvhzv+7uTbmLvFeNhClL++K8S5oNa3mIHKAtYTADjU9
8fR0BsXL6aW+3XVkSerZ985Q4JLoprhVR0o9dsD5GbXPqlAp1dldzOjjwSqfNKPt
Ht8JQlcvfoRsPMqK/73Fjtf80Uml4yhexGqiLflKS9xOxPjGtYGMdsULx00ato43
Z7NETaH/UMhgTmJAeed6iRrZMG/rFFTaqWwmX+S55O90XUl9UUJZi+SuNSEOawtn
TLNTWRHlxvjt1jnxS/cyxWRX1QsUZb+R7aYrix2hi2sVmQnmye7EOWiTys3Ax0cA
nKLTa5FnTV2W0XxdkFUFMAtPk09plgZvQjympnl4EznXcdBu5C9biNVu1RDWMEcV
DeiDPCxGtRBcKU0hODAaL5xiv1lZAnx22qYbu6ssfbf9g+v8i1ZN0RZBUg6tnoXi
hh0Ghggrh79IywUJ09/RW/B9mvgLsm59S2liA/6DXbzAxMF8+FCWRYh/8Sfmereq
85OyNVhHPBbnH838wGCZKH99H92qVZskoZ0nWGcZcYdW7K9bMavvYCHVhaJTpSEQ
VZv4FCe7ACnNiamYbA9j6Nq0AefdlWNnV/q6so9uVAgMN+O8LnOT7qUGhqIulLs4
96GCEokekvgA25rFn4m/deuVbWRZRh7F6MrT0JybXC7ZBtbfIX7IKZn+sSOsDf5h
hilnMVEuPdY8+6mpApi3aPcIFX21ybNtb1d/fXRKCl3ZFhk/LC44DPu8SFHX56qC
cSr97pSByqDttE3kB2DSczZG1k8j6dQCrbKShPf6T12MN2eci7s5dHKAIvRfVDbP
iQcKA2hRiAYwBXA3dvthHezOVsPF131agKdmSX4jP10quUMgw6271Bha7Okn9F9f
bS7YuoakkcbYFxLsdnkeFfyc5rxTSdhdb9Ohg0Lw3swSd9raK4C1pQZgU9F/2dLk
tFyO5P6PkvvrkzDQXQ09yMDDQkfgQttae0f1h9OzNwyoY9TU4cTckoAl440xln0J
ha+QcSdmgm8My3jBGyfoaLC6KlMgoqDEfTpFr7j9r21z+olDHU7cwM+JuMxXPw7B
ngUb89FGeldO95qTg/HGDEz1Ld6dDM2CrNPZCVyTdNQh1b1eSWAtqdkxJbAHWhGe
AFHCfAtkjsCDAbkftvbKBhe7ae+xvQQFWVzNiRGJlEZO3oiPESj0rWaa0Mx3kBzu
1LFJxf0WRIAfNto88Ab3g9KRBY3/WCnpV297hNvHRbYF6vFNFIvJg3VkSn1x7vZg
QI8lUqbDXYAhVQIPu3Z5KpmkWVgAITaZvbT4Vww5HGj0amnB4h4K0Z+KYFMJWjVK
f0yqBQKNvIpldl1FXN3ibxQ3ukapGrSjCJ38FNlowrY3UeMam81PIn/URjOPS33f
JIOU/lJOzz8/zB+QssBzOksgcNKxOtSGXurAB/0vGn3jRbDvP2SeTA7UOXcmLhnE
IbyAzV+1EI4kbcZwZs1/BG/FIxZXWsC3nfxIo/7R2bXBSsAS+KI7cexoM6MsnqQM
q/P8ZlGjOK1BXHhr+V4fq1uWIkDILHadE6sA3nIvwjZag0tQXrpkVCvvybdfvOWg
sL0BF4LTxEDEo+xhBcuVDCir2aZPAjiDLgFutHAJZdIu5vA4Odpc12mBf7Sdhjv9
Awh/cCekDpsIS04Bf043panCrmPWcheJUpImpvX62YvOZriJvGfiS/WRxIphYEpF
TFUKOr6Yd480rnXeESkW8oU4odMEFs0Gjx8RFXLX+3BICgOHYqHgPvfzi2hRzE+y
YvafUwW189KXDCYQT5NDj9lpQkGEATeKHyxMv2Ec4JHcDuNOx9JEKcNuSBAbtAy+
d2bvmmke9Svq8+ZPWS/sdW3oI2YAhKLLYqxPBR9zW6nWmeRyPY2YJKfCysRY4+/H
JvqGCQ1TodtzjB1rwPLgq3RzeVJ8Gx08rpoY/fbEhXBy5W4vav0v2zmfylYWl/YJ
FZ/PLRRZmG659K4en5ZNeUy0pvytOV8sB05L3rmi1mTcZ9TnwWOwOixrTTleAoZ0
QfwICY6sLHGCAbcwQdBSFF6wAyW+Tv3hweWccjNuXZQKxCNcxziWRF0tLe9pbL44
KSoN2/8RnO3AIbwLOGG3oK77R647XLN5Gf1Re+SYiY655V7SqydCnM00j7hvFqiR
eeJlOLvSZX099bPOsWnyuYgdPnwNRoZgYAYrR2Sg2Myh28b4cwhcSyv3cYvAZkyZ
sVQ7IwRq4VoCZuWqEgBmEYuXU+COAJDIWK8zzmPVvGZkXa1goaJFeN0hvGxdxWqg
ghSBH5nu/206JQPyRgqC026tvlcsex8rec8j0tYkAkABs6EobzxhgSRsHoYHqXdA
tsARtGNI5vSBeqwX2JvN3elWq5kR/N+/hmA/DZHQ4fCWHDJNvNyHiaV3gaAEoT0b
wD4GmxqXoD8/I9y/2qfTeyeFB9xygwl18Yyo0hCD2aXCiWjc12Sofn+9hO3HQQ97
XclRtTmKd5qhqVaCdZWyvTCcVWgLYNGKusrfuTWiIZH6I97ce3pra9dFNQA2eeJa
fkvNQF2ERQhU0aUtJNRTPZHXyRFGkVCkLHlCNIafV7FlAmrGiSfu8V6PT701lGVO
tkxIyVGxYKYSVZ+JIflqfwoi781TWBYHEK6T1csx0MzjbBqSYdYqgO/3IZ0KGZI3
C0AdqMZhV4EAyI3zcXi9faBp1tUJ5wvhKNe9+aIWDeDvPBPj7aSFCzsA2ZA/x8Qm
/sx/CPlC+JeLtn135LPkaEMl1htMS3r1asBR9GwWRYPslmkG6bfpATDZbWIsKf9m
o/8lLOuNAC7QMfhbhECCLyuUqnhz3aBuOsEmcdG8FBNkNer7JqGNRW4nWrwrRcQQ
4uBa5or9dHcnYiXMDtXYJ0Jo0GqWjsvqB4TLsXIrepPCRh+wqccKBQzl79L8VNZ+
6kVwvAm9l6lv8n46uYyUYFhmuNHYyW86ZrU7qpPdjLlNOjEUmRrWZh7a3A21LHim
BNtLBfEx7Fh59kADqDPMaNz/ozty/zZxLYVP/8PwAPBclJMrQLhW+ysD50txyyKx
FGQY5bs0S3t8rOkbLXw4JwzAvnETCoxrY7RDDz03X9qB8h+CRJCBfS8DM5H9V7kd
zY70VTao5vJop9T0ksVy7jDkWy0mM0ZsMh3HadmXxnTgQDXiNKH5Xj8xPR3HC9LZ
QjHYjj4YQB9f6LYZ/3liMK36JxYsXQBYx2QC/WeVZSo=
`protect end_protected