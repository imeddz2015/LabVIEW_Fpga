`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 3136 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/9huKRhRMtvnNqb3Z+UU7TahEoHV+T8U3P3ufru7l1O
3DlgtZzb9QxCbOjthp9+wDkjygH0eUfDrEl1ovhZG63YIKCqIgpPlZ81NJ8e/Evl
9EK74ixXzOeBzzSO9nYk/p6+pM+TPM/j/HTnDtjY2pPJjyktWhWxw0q21fTq/obN
WRSb6pVZ4nOT1uwFLhz7c2y5emMxpg0yelwJhfH7LNfdMS9vqCgAPktTPl/Vc2se
gvIlfoV1eE+06zPP4G2pVpjXcwHaHArPdTJFVjU/ToaP+NtXcri6ZwvaEXA+W4a5
4eZymt2jXr6FMF5irzUpZL8GgsB47WrXVwx451r36UPYNb1U3oV9yxrz7cIUsHOo
jBQvbWSEe1GBmiRFzCY7FBDOqMyhadbLOWAQwvzbme4FQeZvGLqIm1ZQOgFefKym
B4p5dyBB+4/4YqpyRfF8h19YUXn1fYJy1gDhh43L+cIFGvTy6ggMDxACOsZ1b+mF
nm/w08q/0n72pJTxW5hAPh2qoJ+HoiYRTVZdjj1rH3Ww+L8ZOuDIgoYTZC5hRbMB
kM5TD4F70b5w9cFmdd014EpntRsVXB1PIAPIysRp6oK42tW/Dg0F+4byi8/XMzqZ
Sb5v5faB5d1lJJ0uKvNRqygtTNwgPlDV7HnFL9/OWVSW1EkL97MC0lVjtLw5sTDO
boVXMZQ3m/E9imaCkPsGPOoCAqOL+QtdDpJrGwWORVssAkT6yOF6eEpVkK1X/ogk
FhrZ/GCRU18OZsT/qApeMv9mnJ7MoZnfSK2wwHnxIPpSST9CseSIdQ93AKLu2VLF
8o9/7n67e0AkoIjVhzzExh1OXrtvATfbOLtHnDWAU0H9MA22cBUQ8u0mM8ZQXAtf
mUT18w7Ui93BCkCupe4DS1O/4e+5tEtLgsSkFDzsS0x0HpWQEHCI1FQGYqG2uNX/
XuB1ovBc0ACFbL+ZWCKp5AOFJBuMhacl4l4SKjMYZLYzv4E72y6ehYGrc7f4OP/b
SogiFLJEoTKO6IxIrO3P9878oKm49lFDYW1n7VWjkgebpnKGXmWm+1B1EXWCyybu
FtRmxCUMKQ7tBiq1Zgtdem+d93s0AkdBmD9W2fSeIO0FmFrxuCjekkWxdEtkrBZ/
M3/9RrgTz9AATRsgGs4cknOrKa8aCRRsVCk9Emr30q2yMnTAGlApcdrW52nD3VLD
URp5hSvv6uaWqyaagBKOwPGpu5t2NNRKcq5Thy66vlm7/Hc5xNhnyWDRxph7ztNA
lIuNBV+EQN8iI1PofkY0d8cXwKbAdaH3ZkkA3yejjPVPoLVdHkgFZqNguh6LNKZx
U3wHvoxD4euCXzgfzYSnb7PJZ/8KhiUiVlhwd8b5PSZfr6zr7uHe7moDB4yvniNK
uk7lK0f0hnsMKbI/Sydq6z75/Ja6Ajy1EiTP9wRlYqzXZIHC8ZpDqTym7rF3StyC
/4O+u/kGcHVpj4uXfd1w91MKVG37NHJudHrUGpZ9ilx49YPPAwoX/rUj/hyYuekQ
ZWXAAPaqyAc+jucZIjnJOH0CG9Q92GB2u8iF5lZUnHRGC+iRmeenLQwEECt09eNI
DZ7sJl/Z67ybaMUNM7wrnbtKzJac8KWZ/7vvOGIOJNTf9F9S5kX6yJqNxBwVZ1ou
izwxeyPySqw+5sanXw/ERixcQ7ka68D5XGoo1mUEYnPJdniGYdHcFYRwM84Z80O2
ReGO82X6YdtgHdFlEdp5OqWrnc/hVhAEQ3qceQ8eLV2U9KqYaCXZh9VTtmyzzjaA
Tbq2sky/6TvdxjAd47pKhNThyVVgTwKqr+ge0jOWB46ALSOpZxj8p4dxokKcI0K4
O6oH+3GNLX1bKYSjLMUzO/gSdYt6LPlqACLElHaGP1IAXVQl1lE9sJskIaWNDcrO
85XCe6FB2ZoZWgwhRF4S+A7MgaGu/YPFDFM7W02zArSokECQoMD2sFEs/Ict+WdI
9svjcf5D3bWujJ/0DFdBH3EvH+fAPPRK+9Qbr7HcYrhq3Yyfrw4fv3gruQ3RWT8y
WuVTKJQABERM06e2SYkcUBzOt5sMGoGqqfUaCk2NpLGWnmwCG2Oqs721Q5Ml5HQ4
sdSHZ/8fP/bd457YU6Hs9lc1W0SRC9CxwH9aG97sM1vmXpsv/Oj6HVopD1cPEkx/
wgqUjB/sr3nX38dLC0aHwe2q3rebn1HiDZzDxJltEjOR9ku/YZ4pMY4L9oiz9t6+
i/f+VeXFHGzzQwCy3vEA/9GMJ0ALIFfKzQ20StUbPnfHQZhw4/EILgRomiZRPsfX
onoHB4gEAp2dslyi6k/fv7+1OmWgtHRkoD0owBH+t+rdQOaML7tmBR4GIXUn6mjX
icf4OlX20EfFd+Gv9F+yuqUKTbPvaiiF+tRmUi8VkmyKsA0K8yzMBTV5QKKShPGU
GuyCgwDnUU98JwVjrDSQnpnFjrJpoBzDbbT0H8+w2QTyOpYtvGX7WdHBZVrWS9YD
Ux4AozdawdekcaqFKnkWDEDT1/7ysJHQoPRg22Mun4WgT5UI/2z7nXir+q/omP+X
YVJtXk1U0jCsKak4XtaV2d7l2y/63r7Sds7mY/4kFLrKUXW0ubnTYiBkW02SQ3Bx
o9ffHF+7hsfWZfpemibPTSyp4m7zR+tNrTA4Xnat3cIk/hwHIiGr3wzyLSy0NIKY
TBBIoRvIndprpDpOKl64vOaImLgBJy1/hgE2BsLT8MuPW/nISU1hyhqwIAsb+EuB
i0IrDZK9rBGd/myz7LGMnuO3wJTlc9djHcMiqvhL7IGiOp4hv71Pjuy+HSs6lnUQ
NNUnESfy+1COtfykwFGnW7JeUBy3u6nAWlgzOLJF+dwVOxiheMa8S2o1N1hb2EV6
tQ2gSZqiKiJBidGlv8iZ1/l1dnbCTf+2tnrkvOzSPMgFgImd2uKMTWKN/S9uDMPI
B//CAvK0n1MxMugxwlUafz+9Kz2VMYGnFYX2zEtOkV821rTOXiCX1gdADV2/JdF9
kXYNVcr17mmYlaVbh173Ezd4dEaARYO4LPjoUT7x1gzkdyNxXl7/KPhyc0EySGY1
7T2wBwHmkgRapIkYI2gXi5PItKDgpo5nUkNrU0pYvbkECxaV/fksunxGTp9ZCFGN
+pzI0t9WtGqqscfTHuNCc6K7yOYePiOoJcsvXDq4/tFY+TJsyXI+ONjMn/jTmhBq
VuRuqorKHZ5tDOBODv7p73xVNFP3aIiDq6C4f/XijpVBgJ1jksLMrMzsQt8G5hYj
hQOUqen/7tZYtpm7tko3nuW7Iu0mJv2Z1cAJJS9xwLTeTo6cA9KiCcHWVdO1ZRGs
Ik22NEZaCN1yiBuwPNV5Oaaho6q91fOQKpTUQe2JZMABZrisyWnms3xgc9DhaYTc
mJKq9DO9j9iVT9CvUNMReOtUrjaujzAPI3kyO7BklSoPBTAk6eUddbpW92s9VRqT
4hV0sVTRMqMRyaBZdd2/YKR5EEX4Q236l9Add8AjUZVdf096uX7B7AAuzqn8I7tZ
aOLDDYzS9VxVorH3di8YEYS2naMTslbZNM6Y4FZUJwnpQ+tZZZgbFkLDn0kaETHE
Htj8/rlvtMeHESMTneN0r6uxspqP9lQiJsLhj/u7A8BJMV2demPUl7WrSGerpq1Z
eg0mQD8alGsP4GaqSw7wAr8egzAxHR11RZamVF4fZwUnkjrzTt8/z7txOeNOe8u3
hPCHQckN6XxT9vn9fYf5Jxjs39OshoXTyLZjUI0Axqd9fZCnoiuu3LIeWueRpYhf
si7HBw+bqW/RZnMvFRk+UUTVzSDdudiHeJg4pMYimYXl0Hmr0Sb0tPzJdkOrAarX
CCJRWcrUiL7ctGg8pRjVkU1J9ic2v6HZv02QU01BBKsqTNsSqjBFHyycqhOpzrjM
SXsWBT1vgAnmyvEKz2g6jeU9og2uxFmAgq8uJ7gwu1xbTu7SqRRFqgmf4HDDceWA
aKo5CYmXMxP8qkJnLVSbRx/uP3D1flpIagYL1weJGQBLElOKoEua04NT3Iv80g8Z
ipEtYnoOqEKZxylARfLPiICCcSpIwyWA3sASUdfwQv60gqpNiXkZNe65XJlvfy4w
evAVjb06pN7BHuA4qjDIUiYRtwZ3dVbKlDgXiNGeyHn/1Hng/vsoHSHBmj4ErpEW
9MZajymR6DCJDSRqIf3qAw==
`protect end_protected