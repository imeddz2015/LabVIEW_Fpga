`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 10112 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/59UwEX+aE7FohaWu0/8IpTj7mav863zUNIsgIH2BWb
Abd9opeuBjbGF/waQMI2vMJTwD1ie1YueHc3nSNpEh4OXp8P5ybZFY89uyGz3ztU
W1EsuUnchJoQgbHZ/sLbgtGRgsrAFn+ZoIeGN1d6RAF2wAESJmYP8zw+p00RvjZ5
cIKFp5nAtYJJL/0ymHGZSJPSlvzY1aEMaBUpk63EzhQZkGJgfNAq6nNFa0QduNV3
2EbXGck4YROZODPMSQi4XKtTgmG9oHBAZIZNoH3ARcQuxsMcXeu+05rVZvu0BUx5
EgQ9srXzreoQGJ35fIkRtK/Lzd1ahYb1t2O6UXgxHYDyFq6yYfopDdLOVAyvo5X3
oWtNhIJeYNE2YNh6LDrXa1kvfYnqg0LVlSOcUpYQnIVsjCQbZ26LtUSB1f56sAGH
Cr4rJ2SFcz6MQeW+3t2ujCQLewPS0SEXgbRMoRs0qsZeZRFtioxWnmKKtgSxV5fT
P5rxWfw+o3yBcE6Vzmvmi5ehqIV1oZbRAACPtPIgeAM88Lehc6vpzZgvrKn+m6YC
4SrPUJbN/K31YQm+Sk1LZLB6kDVzjwYV6m8kr4VMjMVNWhC8mQx23vKZmbmRil/+
0qKYU5OncmBnTvNBiVF9lQFrn+C5bOTh0dAPuml/Le3DT/Z2F2vwlGUNQzWBOBt9
FNYeHgr8agKRM+Bmo5EFhxEP+X7d6P3x3Tc4gjIiKtHUY7eQhe4huvela6PuX3o1
BhRH1vR/puBADfnAhSrnLpNjANa4LLlXhaUUe7eng8wIiG9l9wgwSRchuv02uLSW
Ixee6GgmYRNr4wL/vYmipVX8aPZIZ68vyQhZ6aKFvZ7sEeTVwUOBxKbOKsOmxi8B
2KZfrFSQABaultglTvHVzPsJut5tRxWAgx+mS3yr19Y6S3GB4makqmM/RMKxXKbG
mVZUYoGLLVsP72QQ8MrYyusftM25ZI+BAlCv3E/iTQ8VKbA5LvPofat6fU1qwxk1
KYZu9WSZw4bKldiNNh32i5H/d8N2bF5PIQ9aov7Ps8L25QqVBYvV8Gg93dnOzOPh
iA3Rqa3/1OAeXo+Iwhhm3Kwd4B0B0Ea2R7VjpjrDTpkG95a7Mx0GEnAWySnowsPY
H79tOzUAe5rD6OPVbeujkLGTlQOFex3HDlR2YohR27kDJpxnG2Op1mBi9fQPc6I9
fAYhoQmhJjdjDPnHsfgVaP35QgYOEN4+IBg4SKI8rYPGitz8Gcn5MkFDEyBVBPwI
niPuF9NpU4wVevPxHXz6Nhv4eDu/iPIEBohhi13Y16gAN3Xi0rEUMCUgZX4niZH9
kA3SZ0LQd5G3rORzHB0e5iktldVMeJaZVsp4Gby6Z5LL0+lPjs/P8hshU83bjhDA
FSiaD3e1sAttRCQN0v8usrvwg6wzZ/Eq6QzHFKMhkD9Hzbfp/oC7shAayEgnoE30
+kMv/skT9oLp8KApzOYZzvaNoxxP1gA7cDbhu0NgbumrfJB3myxP/q+MQmRMAuH0
VculSH4zXGAhkek8Bv0JaOG2JSXo+mkjc5/PXzZu+3CyyrEeY/a4+ATevbQ5tpSM
8/pp3veoRaOyY4bDC4yVp7cgjGjHB2OAssojasUwCIr4gwCGCpxAhzQpbRcsjmZO
aOcyE3+9zmt69EEBoutHtbPAR0ugMXJ3xupL+JJ/EQZgKEh9BFcc8RcAcl/CYH/Y
ul5426QH8DZG7J+7ToZBWC31srSUYGR8jZ+ikQTelSP18C9+q/rvoaFyxHbtforp
kK4135vfeo75Hwxv5Y7zv1xWBfz5LZhhx0OUMCSc/OjoEzPbmmc7GvqgcKvTOU7I
Xp3zl/3t9MEB0RH3iSavK8TKvfT/qGKtTPWMB5jIPVTtrcbxW7Iz3j10mx4PNii4
QTlaIejD3pQd9xoeZoF4VFSP2qoEwjIJREFgh33Bj9Vk9h/h2gNPxIieZrLi7ckW
uU89/5yqIybvfw+heSTqv91wDL/+M4XwyXSE9zMrbNgU0tP9yuHO91hPP7ULR/xz
gn9oZ/5smJU3HL1TWbZEMose46wU3kPAke8Zxt0TWwl7VBs9AsN/tQjAgfurX+H9
qUcatngDs+NXxMacKF2qOgV0h31FVmDDlSS27PwAuM7H7ztJakO641+wQqB1izDa
DEWSHcjlyY8ZMWwD8y3XtAy1uccYcqBpVaCl0IoDPWiZfFbdX7PWN7MAKnKKQKuv
R2Eo2PFnN7N+hU0y7qcJANkblmSmneGEpcVYgzf5JDhN9HHDTqQQkndJ+0KKIdXY
ihzvz1urznxqcdHNLzf6NPwSJAK0uM2PcTmzv7YiEivMXp9YYVO0m43Yyzd/w4lC
vydzG6guWneVB2wMYlBYHLbIJSgOzv30PKEXTNNQWiK3letjg/KxjZeV60jouHvs
dExors1KK2dlMVyd743YQp1KM5Bph46RptOmSr6LGaVLirpQ76AA907SWLGopV7l
7yUQfxUZRhgn48YYRo9KX9S04YI14CfeiG3sPMt09eOX9bXt9KTdFqKLPYzogVpk
BjLf8YEWSKDz24TUd9cCEiG6IknLF5+liRT/Gmei55bjdTUuTnE2nwWUYSCycMcn
ncie3rz1mwa/iWzP5A1mjOWu7DC+Gfrsd4xzJMFX4ovdyEidVMPl3tAxgkM7TnIC
DEWR0zXEBnWiqaHO84w3eWzVqxFdAgqAT6xASnayOAZKudFx6WJ4zutTAeO9QB1O
n3Gm4mng+NoQtrfK0L40w8+2b2jXtxZdzDEH1Fuu8wgjX+voyJgxJZqbj8gxZa3n
aiWcA/83REbie4vlA9wKvy/mnuocDncvM6Vpk92Fvi2HmIxS8fMKr1MEncFlY9qU
bKEcmSDenGD01JBI8370OTYScHVRH6Dgx1rbjlMtR9GMcCpNJcnKcpCoRUtxp2ek
fikC2+FxwzBIBmcjBjK+DnSbAzLgDpCfIEff+ONJqBFOxwApnsRJ3D6YZ5p+gI/n
P7GF5fsYuzdWUdThAtyKNRiCrhvpcfMFURvW0VCXSB/ll/7OAsdz4DBwOLOmiuOc
2CyGo2iYlAPN2+EOBfP8ODqUgCYR7rQib04sYr8m3vUsZgGCxmLZ/8UPTCqejXUo
WaV7GrPiJ72H8blvSSVjNujM43l6Lz0fw+QCaJH5hTygc9lKJ5TpB9MqdSjhLQ0U
7aETWMQWd177lA176StysXJY9OLueYGNySGWT8Fhk3/bzGSE4r/VMyCq/ncQfQjv
V/CtM2LtAAeTkWTcMMQ4paOCFdtjAgBPC5/25DRphetu937NkJS1Ee8NO5lLy9Lp
RyZqn4swrdrach4WW5Qf+80m5HlqLv1nPD2bAJ1o65pUL8RC4yyVeH4/UOQNRppp
p1T5hMDevPDqqVmi82LR2lmiiGKzGFxe24xtWha2leM+E9jo3Wx7JrhBym4QdRXa
DQqnmVJxzAZ+P9oXhd0rxgxSVc/MoGbbkpXw+PFRiDJGzBBIP7idwwfhrFNFlMdY
g1j4ea+jwBI/opyFZRzq+3BBmjRJJwYWgza4fvu2iQrUmuD9/7pkKaBQDKREF86c
67SZpCQzdF3waPczkNkWS2IC4OZNd/249gnP9J0rfU2pPoNXOMieVAcMAsrSBWYV
MKtY6dtHWI5/Qhx9u0/IhUlwVVbpQp7VdW4xPmhYj0qy8zr5Oqnf+iEfePkFqWVq
yTsvaqLkttzDLaiBYaPvNTuJKXCnS+lRhg+f981S5wW5N7hFpQS4Af0wKec5KFh2
lqIdo8WIWzVs8mD8lW0vvlUkmNMv0OAPTlY8bYJ+1tbV5a0y2Hw7H65ujnaOV99p
rIpKicL7QwVwuZat7g1iZhMQR/yHlzInBvooZw1EcfuOQ8JZoesfkH3ZV5Dh2TR2
qpbVQbiq3B0EMZ3v0zJjpVMZuLq0OWeEkgS4mtSPdPN7GfQVxYGAApmnkrpTVt7A
gaTdqUFawmp7XNMrjkUN+UGiBfPh9yaDaIghhw8Y4FlxMM6hrLE57z+lCQXMckfq
ANNTd4nUIYZVTwKNgAdOoEBkRt53Js3tVdiRooMQSWcTClOED4hI+F/U/h6r52NF
EztvHojtnUieQVCNJUmC+Q7mENex+f4a0P29WiJ9SXStDpcrbP0XkCoVde9ZFkNp
aHSGj7klYSDc88Li5D/IGoeXSdrF4GcmszwoRrjazMxfVIRQ/xXEgRXTtSZHjz+L
+olYAmZ2Wm5qnc4rv9f89ctXosRWrP6ZN3IukzSHkzZX+hss6KpG7/HvINQNjrcE
/GoqcrtzF50H8nZYbYbm6cOmU6xr42soM9hwekJi9mFUEKLZLT+y+0zItcQs0kw7
JXaYhRDVNcW7uq6UBRPTdPfi+5i6HwcaOQPWuKotFS/qfadxHLZAmtLQYcKX5WDn
kxHlBSD/2ds9Orsp5AdlRwB15r5MCYV++gtliCkkFlmMUfjZpTw1qwJC5KqV14x6
kaRh2o+PX6rcQ8+QC+aqoJ05OQijd1yFnFoB5pQcHhGWJae0XNKirohzdz+tLum9
vVIQGPjx66CXZHAMSGvsl9tDrKkoRZRMN6QjQsezRG/Y2YO4APr2E8WMJdvq6CQB
DEzlIwb7qEFGLyrTnQHp+Vdsg9q2uxMLAj7TTazCNoQuYCnINRKmP3MvkPS+Bdtb
5SWry36DiUtT46kmqzPsyeFoxJyYVIe8hLmOo59eH3Sg7xOfm8AQ2qsSPjpQAkTD
XpbS6QUssYX6l2LEUxRL1GYf5ec6d0KfRI7pNBUtfP32NWmfwbNHaFIhEAKnynCa
e6CsMw45RHA/azwVW3DDhtENTQMExIJJYI6af367UI4+LTZatz+oVRCaCiVIOPJG
DXSpoPHR9WYOctMMlJV6Shm/JklzKW8gII67R0NxwrmVMDolddtiIO4gULxuao/C
+UYn73qQGjRieL77Q0HIHoJ2AWI+kZQbcaFVhAeXu4l/+FrWzyHETKsa3r2jMxDN
QGfczwZRi3rB0Ndyp70Oudx65diw943jlisyBtG34J2ZzpnQ42M+8hUVPNvQptwd
j5WY8bSjnnRhlgyB88xfMzTHqeeqAd/3QRWFm2XWHsleH4esCcculQbl0k0HS1nJ
yju1ttT7wWkDuMUtt0bOOaBekhGA1N4jVeM6g1MbA5ZU94fZpix7G4qFeeZ4OCaB
YaduC3JgUYcz0AaU2+ThFkLC0Z3Xjb6NcvFJw4nckck9ubN2CZYeeuvV/eWV7rzA
euHRXkBGVHfyvb94GXcbKMJlJirrT2Qsm2TS+4ZcP3jgcMs2TJ3/jfNpn27as0b1
unqfceQVwdZ7DASTRn2QxZnguKoAga03UbUpMuIBDaWy2VzzTfMllZ7DTcsTV8X1
hfFXQGEmOJsfrExE4jUFQfn5XMO201nsEEvkXCP/HLyfiD/S8BI9laeg0EIYJkpo
gUcmNKuXlewRRv2CEnuGKVRBvH5f6s7PIzp07fzCM7tpSSoyNhrKezyMjllJ2YrJ
uMmJM2NYcs/HDpyCqRJHg6aFGsSoI79yD5M0/P9I9KK0WrmlFIwX26OrEL27F5dE
6KiIJ4o3LyUgh1cfnrm4uPUtqDNDqCVxvL538WSseIKeoav1LabxCL/Jysory91U
62aDPFRPfngMCKgVVypckth7svdX2o4TzgONyRFulu9H1c3Urkzv+vCX0SJ4PgdT
4XdYVwV2NWiIt5p7k/pl2gtUED9OhA1SHSxzjvHq4oewGngBI+7WpE1fsaBmPurG
eP6HCGYq87JpCtzWghe+V6f+WAnjtP7wTVSIDM2QMp9PisYrWuIcbyeIQKkyhQqT
2sYCD+aSeRmDR8Od7bhkJpTLQGBDjSvu0S4umqV7cMqA20+vqX/4BZKhCbFCYTf6
l7zgNPNZPcTgv4tau9ZcehGHfRb34difDSeAmsB3uizbh3+xQ8LdsqvfPOU6JbHa
AXVrfShf0uT8JEgNWoBh+1KFdiw6fEZUDZb92xVdJ7FLxNRfmonnDfYMyHUbRilA
H7U999bta2okPUJ1Nm+SafKRmilRrlpyVLdVLjY4+GR6v+A11CXQiMvyRkEk2DsC
1Z4KzYjkQe7LEEDeMLv0o0u/ZTqjifnOgXG+XvHVsNfKHqdHxTF5CZIWctF/bmtu
poHmNet6qcVWV4U9Pfm8qVHN7jPM5j271GhfEe9WsRA78PkgvdH2RW6KffWJ+Vkl
vgvsJYeqVM6Yte7E7kXY2IHShyfO95gLQYeKzqYi8PijB/W1E+aSrko1Ov3GVd/S
TKEbcFUl/YhK55JYFzGQrsLrXy5csabENcCrxqqtH6/u+hOt1DtmnkGESkmIX8fX
lNjyiYxYUIfbRCpT3e7wTBsX8M9DMF2H+qiAp2hhHjc8NoA+lMmGwjVfw5zzZ09a
ZSNDRcQAGjttJP6VfJHwoMJgBiTHR9tzQl8Vxxp2NDZfz9aiJXXtskxxAFyhLYQb
m2rAgmsF7fWGk50XIV6zA9prEEvAiv3j1SwXUhL+ND/z1nge59IYdUc6QI/TyC6o
DmwwN0CNknT9QMWfG2Cm/0Oq6OmF7s3g0w4KdRnnkuTg2LgcQVoqB9KIsKd7ki7i
87+m+g8LPgx8l4CsRhWCvKU70MC1Y8OnVogUXvIJaE41wY544kJIvb/B4M6KySoZ
dwQpk5ATCTL4pY+lkUGIeLmIPlkQ5Q7wMez43mA+knKIl3DwVL1UVC7hcddo5hKv
9fhS5kh+6KxSp7br4c9lDYHzj7vLACOzu1zTauKc9W6OwNruf7LTOAQZtJyHzwGz
+lCt3gS3cQt7OadfKnRe2FSOg3meVImRBRzbExN7S3ui6+w7TOETwSM009cC9au6
m6Xvax/fWU6DSfb2WRn33JW3dOylVDj4/CooelgETLkToZUU+BtAVQ4Ec1gXNSfc
l2K5mmBf/UiObJBhDloyBTnHUhlMD7EKxwRMqb0XUnS8zZDj02u0UNAo3RS6E7fq
aG1HFUhBhcY9hMB15d385ym3e/EE50Ou0PnI8DpTcqcb7uNY9+B7tTteQ87xazD/
tTvo9gII0XTocY9l6DGDF4LZm3ld/GpMYH2DMoSLkHcZkSOMKe+JDy9ZwzU3ND6D
3qeDj01zZ8wNYrsSTrrest0aYvu91g5aNZHvV91oxLU4tQ5uTjy2zle2g9/nDP8G
FhjYO5+EFxF6iLCpHTqtshJQ6DMjimazwif0/fMXUdxcgMyd1gqM9USykn55tT6Z
sQj9Nj7pslSoyZSiRJd2XpplLQ8PpVbfgt/T1WB+RCVTsabYuu3hd0p4wb8jeFLk
kIPsDQep9uX5gQ7pbfT3Vo/K17zSe6ztduV3srxNO/aVyW5YvrTmt5OTT68DvYlX
S/4DFHSUdO9/6qFBFqHQrX3vbULTcOO3909MAX7Q/vm9vZiPtUkWy98dpLd45TrT
ocPYavcLUB5OrOQKQLVD0gNcqCNEXcZb33Rh1kfVGyporSKB/KyoDkZDZCB557ue
7j7e5Y4+F/Wii+6L/uV5AhmlqggxpW1ul53mEE2NgR6TlrV5lxiKnWoD2oEL79c8
2oJnELULM8X0ruKB5E8LIArN/v+yrTSd/fzZsyuhpazNenhwpqq8XKcExmYNE1d7
cgdRVkM4wFboCarHYzn68NBm7/ZBz75m6UTpbn5nXbHdZcdIDWKF1cwVxwHxzwv0
T54vP33q1tZIUBkIB5ZtMxkBRW7K9xxs72ZHIDnzRG71WLGaMxAPkvZilEDdng9e
BK51iplUho+B056Fb4M232uNPK6+tYToBfGMwfOqaax4SQ3GrKPxziAvCOw7Xi8m
ynzxHaycMuR+m2NZH0MYA1q7WmCddg99Pcaf1GmmlCbDMxMuFiVPw4f2TjUSdT3V
RSgFuTlbjpdAPMwuSrMZrllIk6B+mTQI1TcUTF6ttKC5g/sFVrOo1XMNntxKiB8C
AiLcxZsHWiE3DN+2jirg38SNjiu5gmfSI6v5gTiKjxXFfDAWPTeSSR1oVO0FjAne
radnEgtAPdjO+lVexPSZxYApLnnjs0VlUyH4A/VPdT1+wnKWYmCHCVOJ0JXdtyZn
kRdaIwFLNIAQIusNJyPZCNKa4tbTvyvByGiXCt7+GXNYLe5LzWhWNNLdgpZbNJbQ
5OZHUJeC8p35cyr9Ucewre+pbSDis9H3jLCNrg+e/wV5Z7AQNV68i7HLvj2hIEWP
H1VFepjTkdMpkdzhwdXSxBW2mLixE+1WXMxEMWMX+XFuQNHFrMaL4tpf4pMUCS09
f1QMDpv98IYM5Ps5TIGbSLBrlDlZJVNBTtZ4DwNNAPn4iePLbVe0ft890Oj1W2zm
SLxXWpGyV0m5XjJc5qrRxA5jnGlCSx/0kpISu3APqJQSn0DjQnb3ju3LLizkwbDW
FDunyW/y0dgaonzbfaameAx/D8noaJWhzzSkV39r/gFGGXdHFU4IS1TN+aUb42yS
fHCssnZ9ZNfkEI6XQ3P17wN4eLv2SSoCr8OIIClRzsdc6AOYSLw3W8Sido4b8P32
iD8Z/4iPFM8px9Jb09WnQ7PkSlmJHIauNdTPVRuZM3rosKbedSiyNCOeZDWvK2Yw
eCegZUwdhsFT0YBsBuNZYmlg/W8Eb2t2W/gSjPA1affleu07dwBBXsOpF7QvmJF7
tskAIhB4kRdvsLC+zVy093abXMO1G73pINpfBDZpy9xYtWhaexYRwi/RWuqnYL+N
VADGc8Ljs/BZB7jvWCEH1BIriHFlxgETpNR/5CAiQBmT+L5XGpjEY4fvSAqOQIU4
YMV4mUQ6UZijXVssbPZpDlzw61uJuea+f14ED7T1FLAt0x5mzcKJZGXva0CPb9F5
uQVmy+Iuyk1jeqxD0QWkUHduL91iGJi3dNdGokM22Y4+GZEKxnz2O/7AjP2nMDU6
Dg2VEieHHZdVQTV0FGF3+KSU3bzZoGpFDNu8Nm/ZMWZXI27bCUy89PjEDTS8Icg+
LmIs7oigcxc4qbi2TWe5/ydPRmc38plmFctO9RSQ7FBU+sdl68kJZ5doM7EQAR/W
Y+xH57BFubTJKxH4yqaZ53CKEYA7JBAVrV+uBdFZO9UgFFmcfUsGbxMIAvRrDHjN
l/2dkGUTmJhaU10Y/dHtVy8MoMTi5xBNuacxrasuVT0GlZXOCFODis2nKRt3pOl9
USXDbgYVZNbqkEyaBoUrhZMH9SYEnO1llB+/3wQj6ZP0/gmRLOpkw+Nej3hApxry
Mq8fsGvr5VTNQEepvggS49ItqSULXvALlGsJXJ05ozANyMgdJE6sINus8lkOwN45
7yzbQEH2/yHoZX7WwygRue+sIzaZeOGRAQG9AbbR3sXEMutEGylZw9j6KzU9eQBM
t+q9vdXI8CdxS2igyUa85tC+7yyJD1eLD0jVUOayJ56tb8xeXJVlq/3zTvoyL58D
ts1FdLA9xk1Qonu8QmR0LEVFv6tHbJll0HfdM4kxDtmcdJkuipDMUN3j9EqACrF5
QyJKpJF85fKYTd/DWYV+tH7mVa3ZKMKK618eWJ9S8HCNjQCrNYjugUsH+/BQYHZ8
NuksjizhWn6MFtB+afgI/wf2k0dT9qJfekxblL/a7gp0YqVVt+ilwRKzKECJAOun
sRFoZM0PzEc+ettQ1puLf6+SAN2kvEzrIcMQwr9/J31uqBaRC+lHTKEzFE4OEkE2
42GnlV54TAzVGEvohuDx5lvJKHe0sYP17+KN7VX7Aru+SozixcTGkHdwpe9BpnKF
6CBQPXB2aJ3XreDLvWq9/oPj2CXChrehy8wtsDjwics00ZhRvft0RZhzjNDvAkYP
f9ENVKsoOJTQndss00ILyFH6yNuQ9HwidZSR/+Oo0sNxXRkbRhvR7GmD+f683hRu
BeyRMbv54K72EcztkkvnVHp4bazMr68kF7fmyAJpMGGZG9eUW9TGPzcavhjAsaRp
zfcFjYz9lD7O7fZWWClQa/HNdScuc5GsfwTcGqF2WVKbPGhT3mOK1SlCfxjVKAwF
qg39vLARrIqnhu2ZNg1YlLmVKEKwu8rbLOWD8emXxZkwnuhci0PMZYSnaATkCQY5
6eePOk8IN/+++0bjKGUATg/AJ/SlaJLSsgQPZlmTk/Izi/3AEBI7bZNWGrlRTRsD
bQza6jvLwgEoUQA5YB/Wi6N9Zg4ZBT80oFkvoKFPkzapJdt+n6nKXcOnqcO8K8CN
fjlXX1z5iTbrZWohbNIomaX4ADVipxtT19y8GhzXhgwZYDbDoCiFjDgzLZWLAJUn
NOjyFjx1mVACDLC5uuxzDa+T4aosmAKalBCXlGmJIdPfhEiSOB91CmSgz5mWJxlV
9n21GY24WgbGivNyRdWQPraHMPL/ezxHTMoxC/n38zMNS+4C5ZD36R/zHJjFpvzb
/l9HEY6bjHc8pkkJLtSDK0xF6FGDOAiv95SqE7sBxueV2LJMC+nYY8osAsRl4QtH
ylkQAHOXpqLZSZYgomqCL36i7qifjLDq8BWXPLJScB4ChIiwszmEwpUeen4Fxycj
fqaAWp8YOGh+jEfQhkSlogJ2uDiDcTR+E57mXVt+EtTDghEvpHLFvkeVMwUe/xcH
KLqfe2gX40q8gGz2N9oHU43M2eDLXQI/rBrDAzHpMJ4JL8Wc9Eu+gUMIQ/F6nscR
JgDY2hfiglCGl9sAteYP+gHRfymkxJCDEXM6axcUcadaucFonmlPzeR9GGvlVc11
Qm+0Oux8IS2BiGE2NPdAxCMC/0USWhn827hZrCXBLw4Z+mBWf4Fq22Vyv0D+r9t/
yRZCLOQNCmjOEVpKrk3TyeIA3OUm4EOg9bjEuBlq3ytyTkAxXWEKFtJeR4y57tpO
D7hiyYgdS9TuxQ63X2uaNXIuUaoax0+v0fGz3m+MLxcfhDZFM0nEO2XmTht92Vq6
gyahi2Dx29eUnxx0VHzSH5JBA4xcoejSVjnvJuoU5iR7O099cJVOn/UZExK1Fihs
kqzk0blgIs42tq39X+G/b3fu0eSSbCXmu0FRNZLGiZFL1DxTs75fa02GdWO8lxzP
tGxQl3bGwhHVxif8fLNHf32i67/TZMKYlfvfqx1BluujoIDPBYQU7VprwiHj+EV2
ILgspP1ghiMRvxoZoDKQ3saWNI7FSwAPebOn+4gVZpHHlAKKHWSre+Kvr2rBEuO1
BaqL2fzrapEyx8gEZnXGIuM2TMaTHtFe4+GbB4AruvfYb6fFYQbrQBlCZjC8yNad
C4TUgZoulUcljhssbftVS/kbRr4I2esAjaGcJ/s48JnzEC9pmkDEy7bt/pJhYsjK
9wHWCnD04zitfMTzW6ZW/+pM+DOd/YqhQzo0DADyVWyIyLQUnWyyovaLk8SGuY/H
1tCXX3FhF7G8s5LdUvGiscdzHd+Bm38mS+C50xZM5BDe8wGMxqmQrYCneLILOung
O1tsqq6y7O4xojPlFb3QL2n7YTOsjJqBRMIIxe862GooPMcEaN7FMm7WBXzG/imu
GFa0z+wsMe7/Y0sCwNTj39mv9iILEwuJZ9Gm2CiiP6VeimjuMESN9+2PcsQA8fcL
pQONfuj8A3B/r5e5D6nePsmS9bnnB68cIVzBO9YLCQ5d9VMgLtO2Q02S0gRoDSVj
6VFP1uU+t9goh3HU77JCaxOd0RjCMh/t5/vbSAnHu24F6TEf0aV41oe7Cm2UooQc
9sYCf1sVdWGaVDi9qipLmmM+JkGs2i7sWl/zrwr/uB8x4PIl5h/Nc87AXFp3/CEv
2Otz6UI38lqNGO9yVfvybn77yCeXW113ABcrzx/KcWcyyXefijWnxBxwd4iWWSDx
cIq22GeWj7K7gWBU4Nw0L7gxzM1YinWuE1JgjQaX1YuSUrXlI593A439iDcAtRRk
IVy85BkZDO0BooeZHl5tNC4mUYoR5k2ShTRZvwX1Fat5qDDe6FsYBMh6t6/IKWb4
WfuCpcMKiUfBZQGVdl+T1doJwzrz/O/9KM6/Rhrqp2RZCbzlISlw0gGZSZOSqqCs
8VdS0bpU2WzZbteeHlKdUN2LtW9gar3rrVIBKx3ytt/kUa2ncoXmYM+0bRb2HcN2
6Ypuk1aNBqAnynVq5ja39xopWk4CJf6p1eB8TmVZ/l5Scolmv6MnNdAscyXvrU/+
oeC4NeeCZOtRElMVnFNYOs6CV/K6T2qJcFAgYVB6xO8f4T2PJXUjhzVPCmaNalgw
lievow3LV3VAacpzHTl3b51P/3hJ66WbgdzzbJ2VkYwnc7x0QEFYdhIgKWofoV6/
2B8RFvlSmonIBk2Pnwp+7Q8aJj5uBleH8ELv4K4s3Ly0HOeoVdgfPZ+XxNL0+hZE
Z9p4uacvXV+jLdirossShZFT1Txy+Wb7tDVQiwEx7Q+zPeJUW7j2kiIJfc0unW+M
v9WzZp2+qlrDy+VER/FeUuky/y5FwsDF3pfW+dGw/ujS0Kje3/8lLt+bmY+IQnOB
vnhC45uhrzin2WIBhJgYOKMLxBEThRxxiBaTsu/6xhHBdEWJzdL5JPRPOVw4emVt
udrvitcNMBilyEYy+Wy30/zsIpyvVtXkf8O31cocFyXgujPd2fVF0imGMMOpETBj
JOckE9/wkS42r4vtFib5Y1+e7Klccef+t8B8HLcvcgv8HFsFKENSVi6nk/JEoziv
N3nqp8s5dj0EdZcD3pchZMgKNCWMbqR4VQqjrFsFBeu/PpKXqaarBTktkb2DUykW
9cvg2R0jxJXy4H8StwlqaqKCUI88kMCAw6kyUv+D4K//iqMJdOxx2a90/mng+U49
FooIIAAdGI9Bp3qbsbao3Flh3w9xl8mIDMXOqKh+wqn9x1EAJcx0xVaB9p4pIt1V
TWVUrsTenW1nMZXN8jDYIYXXRoy5btaTbgM9qiqct9rfVsYC0dSEO1sP0lPJtWay
PoCk69a2eCm2OcPWNL5L9Jp+fLA9NmohIXzumkrHWHMie7UKpqAXiYCRPh4CuoGh
6MZDPY1R+XsnuY8fBHKKu88pg2iCh+k4k5zIeALBn4dtxlFrqT5+cTq2yzbIBt1e
ezmideUvyN3qTJKaPPDZNrmuptwghRlKd08ONTQrDiztttbzPMN+UJCVnruLcjH5
fohJq2bMQDzBpdLLA1DwfXky3w1PVqYqU66ceG7JNQVNS4MFhhnNqhoBF9XDBtcn
OkNYDnhzQ/d9gbNVfIV4u60F0gzzifPNU0aVJt4L1bNKKb6LVhVif+tQWTeZGR+2
2ZaU/zXEtrSIfUC/xlTXc8x7Mn/6grVCCwAJwWDO8kiZKrbikOMXuJLoBHUvn4+v
9F+5wCe+q1MQamPYp+XhOcwhxhF6+uTvpJuMjHJ+u6ZgOO5LMwn1apzCtAObREfz
gepODNtGpcJfR6NM638qEHXGXy6jMK1IZr8LUu83nIRtCPS9/jEj7tVaSEdgMnaT
9VZWjOu6LrS7rSZIawiSZmfhcmaMfU7IP0V/JmRaKZ5SsJDTBZ4g6Svd+6bPvoWQ
MnaJN8CyInXbfop66HJrPfbSSz0rupCPXVc5TaIlljU=
`protect end_protected