`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 18496 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/9huKRhRMtvnNqb3Z+UU7TahEoHV+T8U3P3ufru7l1O
3DlgtZzb9QxCbOjthp9+wDkjygH0eUfDrEl1ovhZG629lG5sTX0R4F+QPmxXcLFU
UJ+GckzRFU5vJTnsic8aviKz0fWCrcGC5y7pur+66FyLM4qFHUo73MIh7T14zc40
0pSEB2lz+b1G/iBRZcPf0DQbQhv7ZeTGvX5JIR/wSN2EnjLb9bghRnfYyxOyCMcx
FvdXT2CZQMmdy4g7Q8/QJon1mwgyKgwD1Tnk/mnBRRsfawFx3R4BiCXgBuVyxdKD
qin2ceC37QF694Wl52QA3dtRboLzJqeFbZrEXFOT+DTXJ6zlLXASay28AKMUCRX5
ZelL0/9Av94WjQwaoyAAxP4SfPyTVkRgEWDWDuRTxvInUtzyWkE5yiRCIU+gaQe6
1h68aBVo8gnse1RFoy6xANg5hCfMGq3JCgR8I0yAxgB5GGk5kk1WMWaxnyNdoc5J
BlMLnTlOv2P2CjRumly6DFe5ZgE2JSgixIgvzqRPrVAxr5eyUoBdSE2RTN0papzt
gCb1JnUDNE7ownXfCmUpLr63+mL2oD2sPsuKnMJwWGgjJMElsIQbbWXeM3KPVDk0
IZYiIqVU7ftxCdTbCFx2K4tL/Ylno1Uc62beTb4iH3DyGemxdnC3isG3+QJasuvT
2b9+MxgQ6xWuIXbD2EwifbmfKWDgynYo9pdAkgy8iURkM7pdTTYphIvRBLl9Xg47
Ko+XMI/ISqCjB9rQksNBLVQi1TRHSw/rEAOOAgzcNO/+XUetQXaG5KmIgLE8A0jp
TfBERob8jUuLE8847fAVRf4HlDCaNGKKCn5edj0nnvV/QQWz0waTPTl242LUuyRM
CxipyzU3mNnX1nxq2vls079S/6Qs1GcsE0ylY/uirjXGAX1x70k9/vck29JX6wLg
5gGInyQ/kQ2JAex8uGK3XNXm5WMGOe5T3+69XbLoXBdnAgRDePOupkHqa/lvJfVI
dU168YXwoXsuB64dw58WlihlwNe/JQ4DDL5colG1NNkeEwm10129ABN2sinQ1qHn
/aB06bdM1F5CUuhsM+VzycUfFHBj2jzWj4PGn8gbs4EVyd/2lymWgDJql9jYqSUI
YXif05WTlzD6oUIIE7Q5RaAH4wIPCWbJhxjYcrSBLnjMB4U85OYB/UpwEu4djeCC
z8nNyA88EE3hYcbBf9yO+v55G65NMoTBLzZJzwqux5hxz+2c9RKiBgxE0B4VUdzc
OBUNoNLr/R9c8Yaxpkb6I46uZQnO/z2HRh3hY+JuLpmdV4ymvzjeq75ljm4XnkwN
4ubzyUcWoJbx5Ue7H+7JvfkgmGOI6Q75TKdx00vF3ZnMgtWs2E0dZ3dXI8MB2LuL
S1qMa6jY8ICQM8SpS5b6OI3uhrUyM7eOnWi2esVT6Qjvfr3Lb7zmpkpK1Id69A40
+wgQEfe9o2XicjofUaSGU4jPHw8QKJMgu7goTBvhHSqtHp23VqNQYPFgGGcRTw0A
TnaTGguEvA7wOAtxixWc3iKkqIArYJZTIZLRcKMV29N4Hreyax+N+1y7qeot4xCi
n74YYBRt+cfleXdhSLi3KgA1acRwmAdRwbsc61dUHnaP7pL7wTWtL1qR+D0Z7y1W
Q82yuz+h5Rwz2KqPUa8BObGKcBhh9YiYXDHn4u0hDMPmHYHOb2olCv7xi8evV8u7
XT3PjcthCUaLPLoAWwbxIS+1uWlZcbnyYCOKqwwkg41fhwf+zlVoKv7zroqVeHTW
Nd6uFBv+YcgGfENJzPsZ6Q7WIIXFH/Zg2l0KasKrVQnWOVWeS7GBgbYArUqs6Xd7
rBBX6/avMzzt3Dxn/nONCAs5+BnR24zNlkA//Man9WgcnlpC5Rl6p7Di2r2b600L
NUFEL0mbpc1hidsu7QTBFv5r3CE1Yc+CQMqy5+SW/y+hsElqzCNrPyTVoddeJEtu
VBvNSLVcjTxXBJPlXC4sE/g5l7yB0sdOcynw4dXSMA1n/PKpHcfjJeAF6dAwV+fK
IaIJCAEOgjERmePxbBFdeLy9lLcGNoZ8aULHcWrh7A/OGPf/efKuhXYpDGH5sm5y
iUn8e8KRhnkntjE1y1EoGKfWIvWfUc/t61asAGIwkXqxQOAtzxAtCGT79rHOeliR
8fc9bFcXSw8rilo8oKfS7CXDeyifcEoUj8Cb3iB0Ig1Dkn0UNwUOTopkpxpx48Fb
oldBrCjkA0TyArl/M93UVHtt3CU9QF6wwCeVAfGSbeVULpr2l43yxBabHmpeQbpO
x6RrD6wjunhQo9Js8g5du5XNFTy7E8HuYbZBsz6zUCPFB0nm3gVjg32atzywcDag
DMPAwciI3Y1Me3FnvDC3P+ptAIYHalzLYTCHqw3WQNZX3GsGn0oLAjHyuHcM7uYL
mOA78GjkGP8d3vdaFQSZ173Al9Zovfae2x6Hjy4bKSE3WOzV5ARsZJpoRJO1y9RZ
XLy8v2nIKqZt4s4WDuHrccHXP5H52/4/YK0aG4P5C317BbDrNxEw1EAA6V98rlRW
+k6v1fhhqBmvwey0N2SiVpQCMHPceXcTPy4wcbH93YPEiwQUrHXtlEhDM8Y8h7Sf
ATRyB/JMaRuSxxTBYdGB4y8rrb6fr629jnLEDYz9xoonfpXvqML4D4htflV5pvbq
AKvtf0xmHc4iD+oX+MFpKyHo8jqRZNd5s+/yRf4a3QLaDR9SQ2NdHIn7wyQujcVY
39KtJFSnOdKlGgpmFfmH/aoPBEh+/4a/mmOzhEkPXx3VefXLNfwHpQtYmB18FMQT
sGcH/tLY3ds3WpjiqA2/JWv+0A+uFe7D+OVZYVmPkmZY8F2bKluMid1w0Zr1ctbf
c2/Aa7JAokTLIiVYp/KkEwpeJdi7DQACVmeP3Rzqd88hnf52UQ8a0yRjvVDzNPiv
UPzHhbQwb5LtnT2XeN3mFgA4l7mbBTXAfVnkLgN6ClYwWk/esGDWRULdjigmth9N
iYnyfbGjzrd1ghj6Ag6SV8D1cVSSsb5Wdy2AW7w3Ctu8C5uXIZylyfYswvsRcYdm
TQSVFNipruPMxOoqYOfkVsqLvT8DYIHJb/XMKMybdta+HPBc3XdN9BVoNnt5M/q5
Bsz0pfSVfp7PiGC2fqpKfcDJtWDD0d2UNpbXr/9xRq8qrKVSMCJh+Azgny5Hp3JQ
2g6kN+wQV9EqGvK9IF68N8tWp8bE5AdN9Z/Br9REexiRhGRHTig5LHVFjU1CwrP1
HnXUH7UngnmJ5jEvYnbY0WEbsybLM1bgXLCBXFuthqSlkrxNUBV+RL8vugVLeal1
Cqc2n03z4LOKGhjIELEqqGf5I3P91u8KiCD23Rj6ld7PgPwDoIEP9d7YrZQquv08
uaaOHgrMTmdmhew/oouoD0uFjuOpOJtYh1CB3bQpHQyi2eBeuNjlaOFdRn1VVIdI
TQxTbl+2NoWwC3KDLpmzY6Rx1DbVMWRRDymvuQM75/IpbkMggqSJrYhHci/sEtA1
9YlRKsjB9cQFQcsBch69SxpiAv9vHEk91rVG+tQhspZJs15w4IAlIhjHDHbfZn9j
RPsv5D/OelvxdanRNcX2glM5hdmsquhuT76Y0SkYs+I8aGUiK9flPdWDKzDYo0Cc
SSq8u9Gyu8oAsBBdWz/1NCNzOFKN+HeAo7SuLdaQIhsEYnYc0cGEcxgoXU3h0Ofl
1Za3O0mJZk6GguIUiBnHrgqfoKKWSvxp4gEKuDQBnvi6SJ2FfYUzezqj95zk8Ou2
SVcN/KnJKOzi9seWB9eTq0RyNbQo3w1QOIa61IRGpZzLOoSFVTQPqNdtmkggNXUA
JtJagNTtOzmJN/pPAnSTkO5kLYDxVfs8WDTh9jm+oQGSeF+VQmp90RiHb9+eKrdG
4/M/ZppHwMhzcP/vwQc25Y9gWdAu9dAYZRQaUZjjj53KdeBfRENUm4mU6yPBRayd
e3PwbDMl5maQg+xIBlgE62SovYtwce+nFy4V9ZTpE4TJgnMhCZx4lWd1jemUDC30
QzLiqZxLr0QCPx3cUfMfnoLt33XqzggXzrS6UpjsI//nsL2iaQADZpGXGo8KSCWa
l8x47eMxy7UG3+Zf06rHIB/Mfvn97keT4BHVbhLrL0AB4nt0KzAmrOxxSC4GuNYZ
yqOyi7wAVOxde56iyZl/T3kNjtxMkMifuygST4UDbsPs2vAMuz0mxYQHLQgF10kZ
3bK/OAjUqyv3VS71AKnLub26JFM0K21JbA6ImqlDEuna9JJNgDbrDEnTyQZZr55P
dkxgtqzx4GSVUryhG3/r536gwK4stmh9ixDwMM5x2s/rgT8VkkAtwrVUQBCll/rB
Tj5/1Ytm8ShZKcjdP1yBk36Hj8dc3zPW8fhnZhrqn3ExNzVN71+4QW6pEg0C7dz4
xs8JwnajlOccD68Byvh4K0bTRZDnux/YVSvf1TNCZ/6VdcV02+u23BnP622hnzA3
b7+tUaILOh0Jsd1ZRh4oJHWzL3pnImoE5yXYY3YGKULOeXY3mGqGpowV7wkEiTz1
tmY9kxeNgq9awqg1BMkvdk1KBmsQZAgWa9JANc7KYyDxuPtc3EUb57u9/7SzJt8+
hllqCCk5lyg+7JWjt9vQKFjMSHfAGS+Dj5ZwbYtPa3WJREQYXB0G+HWauLYj2tap
eABBGwPofJfH0yhkSDT+j+rLsckKUQ6KNpTQ4fUzJj0PRLYmmpLFNY/tdzWQj8N8
bwgJHzKwYhk0UA+adQxAG5N/gCOnsydREqvW0pRcUJKpZJB0uRIMmTDckedKMEh5
aK6H4kEx24A51ioOaKuTSqYvVX+TaAA/s8jVNts8E7V8TBUflxqx1WfRpDz/l45H
+Z0MehMTKt3/iY2HdbIwWUKn6np5/qj1uhJv8ZuDP5J56ixFNdAouutH/o+sAoXf
M6Xujl04BfKfYgXgg5n7B+qOwizofYK4KEePP+1/kKj0An34un+pxnNyEVyvGmID
dQWyYwcgRFCLMSRUj4GqpmEqTh8ZMQdteCNxeYTXeta5SG59t4MYDTYkdSpoFeRi
7CW16C8OqSXHCA2TLmJCvZ6r2K7eQ8AlNnwlhFvloCxyqS6CJTCUqeNXfpwm8RTt
a0a9J17wLfwf42xAnA/pXdCCsdcj1L1WJc2J8jDazoWezPULiCJcB2TcVoPM3WDF
N7YBGCat9gR6US4yLooPXcNo4oQ5+GUUALwIOTDL26k3yl070hD3u1hdxnwEBx/q
2g2lTZ9ZdNQ9/MZg9vgCHmljW/iY4iikPAYgSwFLgmzNe4lGcVLh1mnuCbG2XY5X
TUngk3WB9F1G3+9FEAd3JdH65J98bYgkdLAG4SbRWwd55W6676II7220cDTkW3W8
0wSpraBbE9fcvLUIrSQOdBiGAmzlYfy5bOncQUpaYfyJ+pSZdX/ijU2Pu8Jk6O9h
ffxvvm/93FoXMMIrKAQLtMrCa+k5gmpErq9+tYAMadvkyUFvyLX3mdGo+BAQfV3i
w2Y2BVN5AMEszD7/AIanr3IpfMRf8juqWpgyPH5VgQYaFKmQ7/lqZO7Ma8rdZgzI
9xk1nXdrwCwpW2uPGeODY38Lbets3j1yoagQquV5jQCJEkd+dUZcW6NEIMjhyUIO
pyXZNOIc4VNaRihHazcGmBdot1XWaeGBwgUvLWrp0TE/XD5EOVTZz4nM3VZzGJrD
Uo970x84vobmN0qMRkjdL4UBA3QZBO0Rioyy1x4uX180A9NIp7ddPM9FOFe5jkvA
MWcq78lTUOgsyRqt38aiUy0SaXeg/mLQURtPe/a8fcDi+aibOZykmah9wrm3JRKz
dUjIqxNuqQ2WAGNr94vErBOkfV7FDQATHvpRj7CuOQJxrmETCVAfJO26GTcyiajJ
R5KbnZInBExRyDmIUsxy+pd6Bx51KR5zrVAyI+Gx3kqpFugHrWERHjDfOWZxwFFy
FgKt2h/PQ/dAbt/b/nApdVdcoqkz19LhmY1Vj9A9sqTLDOUMtPwQoYocOmd2u7ij
YFNRAqPfsKdnI8cGj/BUM9NqFmeVOHdY9AGxepa0xtaYyEltfgnwapwwT9NyYorJ
lnIHQK1bFK9PNxWFbNIC791bTJ3NDlZ6CDvUmifQwMU4GXKt6JINw++GGqNxYQ1T
M6Himnp14h43d6a4bUyA9UYwlBiIqL+K1LNrzW/uGr2EAi5OM6RbGS0kICTQLQ4l
UouMh4eVQo/rKOoaSA8Ag6bFOX8knIr4E66hJ6TUQZSsMb6wHXVBw5oXgHMtWaRA
J9YaOfabIVR3sl/yFrY8YHl5GJDi2lldIi8Lhj/XCEHRC3hGVOwNCgwto+zgHbSr
fURuCWV7qpvcsHkkk09+GedQZe19FxrDyoQwPZWyVFb97noHezN+5L9Fe38TZdKy
Q48eRg2nm/C9e256Ds9dyqxT3ff9U1rx5gtgJZY2IK6ZjmozRTpNarI2ZomtvMmb
GwwmezsEObUdwgY0mVsn7cEfYm7G/iunrczz+WtLnrlWvPlrYR/+8LiDYDUsa9gS
YnCAAzHcQU8hB4oktE1B7JCEKQnJo7mZFCTwl8Qg4H0G8Dyd66e/Sn3EEUWdNwEI
zUT0p8C89quN8iJlr46MgSzHnDv9C3eIk7hHLhNjwZAgcm+CxyK4t3h4xnoY1sMw
huZPX/QK1U9E9ri0K8fm/lsPs1CW/nuqK5FfQKedO8o6hbsZw1akG1g1ZpoFBzVT
PdQj1PBrVIRrNcqD031Qf/6Om7QXVx8Nu7NzP+QDJS2wkPkNmGswOBqn14oa5XZT
NfgVi609Acy4kropndkrU63dtwCu5/wIaDTtoVUIHXpvikq/S51h69ogXjLGti1s
V3iTmpyjH8OA4AgnRgK0zDRdpEROzA1lh+dENoOzx+oY/zNTKCRTaqGv4Qhyl78Y
jAcI7gqzhiBcQkUad3w0alnMh3F/PeVLnGV7tESONBIk8KFQC2ruDRKC1INSE+uw
y0iAPsnz8a0Ynsbexrdyu0mqPTA69QoCtKIbWwr3fupGknfFarDRUuJTjH1+fGDV
NsccJrS6A8HFdih5RYcg1BZ271JCkJBsbWZhgvNOGeX0AxfgfsFujbq4IDQ8EN8A
J7pX2CsOWtwgi0sbG5Atu9AoPzV9TFJU1qIqEFlSdN/b1iB8/LgPI2g35rNWlUGH
RBIeksVTW95pp6V+B4TDl6gjyD81EMPgPTSCYpsQWkNxVDHbFuvfRqK8vxCziVHT
ircjJgEf5/B9LTok18G6329qXPS9o7l6nlIh6JK24AxKyTTWIRBl/A5pgj1BSXBe
tUFUy/0M8X8EINLHpE5pwTwVdjXc3tB81QVR4ulfacAyIGapiNnW9vhhSWRGKPFd
RuplX63VdcSnTVrwC5B8iuDW9DnYyL8yIJuLcN5jnh98IzmGxbsY71ZTdwPFjcMd
uiTFb+1M7NceNRadGSwKpTHpl311YfVuNM1yuWMbl2oazBDmYa/k6G7gfCHz2xAw
ZySr51S3ojxScjQcYnkreHJXaVTF5WJSNt/A4uOhPmCEcl8GOGIcviUYSu5tiK2J
ReKoGQCR3mtoBN/NBD5kLwR1mX6vuH48pxVPxFThsTG3JAMfKK5BLnn004t+IU4C
4MPCeZCQrNv+P3qoh1pwq0BslYCxpefB3sojLg9QtgY3BhfyI8G+RijTycWBaJej
fo823dZQsZYwP+WLNcHJCPtGm8r6Mce7c9H3JMZ7qhTNFntF7FYvsxb+6Mhq7gHU
AHFjAC7vVAKfYMFxe4ATWzZOhP49JUmkCcrpWe/z5Gw5cR+m8NB9yIblmlPAqFH+
iN53vINPDhf9OqJhah3HGvH3DazvHGbEI8OTRK0e2CW/gzFdhAokG3J97tW0+PWO
UHhMS2SX7tFRXYeaXoYTjwHdiaFLv3a6REve6CwbdC9fKgT7MIPNyNQSkTXKXd7u
qnSZd2gIaVO35ykhSNwaiGpSZMVRptlm5JwbTqI1XgS3m8pd7tSGmOOeVJsQYc2U
0AHMYjdAypePDVgEIikVej2wUitBPnmZDUurQjX+5drDucNYMjPGO8xk78Fg6+gU
cb0zvSkpr45FHCBoOBSbe+aikTpKcPCTuOcaM+zzD04bi9HvQizTuo74nNTEV01F
OoIRQAbpso0WiRK57KIBxGJ+YGeDZrInTLeLNPCRzLuoL40NPWn2GRrsnOPGXSCM
FFXgJZhWGVO5L9heRu+bJbQagFboilKE+4iwyBj4ahs0zZHjHXymeZQuunNMSAQd
5KHijZSNygB8zXDkeVXvQPRtxnNTSnRAPMPa83PFzbgtOKRFxrXGZnsKUGnp8vi5
/6IFqll9PJSoGQY/11jvIWIBTDIpKMqw95FwUFJKuesM54zK+JBBoBPLmbAhXwKz
fxGA/9G+0jFpHbCAE8j+ElaATKifTYE35eK6NpvLR7IB3BBx2N07d/igRrKPQEaS
4d0ZlugOB/sd8SYBUs0ubdhcp2eyZxoPEKRMqNqDzjRY6RzgiQqq4duIXcJLR35f
+aMSksovBj2AYxc3gddhInxd1SANN/j8AalH7eGG2V4z/zXSmJB5Ah1+ni36V1xg
iHT5PQZT/IUU9XJi/S2LcuG6xxvZ0Ag4O+AKRZpuJSORAruu2thZe2yTvE+o2VfE
vg76mj2UKwkdgl2xNXWMnxQkQIFgo9KZKIGciPMQx4btNeR6K5AnRTl+WcSUR9ns
gK3RsPwkg6gL29TfcDObmbQBrusUVo25a50e7eAeH9DLJ5o55QNc6AA4BNZYoU0+
x9rcaktp+vzFsgLs0kp106GcfJJ/n5mPyVxMtfHuCOsHbnffThZM6bWkX34F1QWM
2eF0Q76J8kanaXTMxeLom/eO7D6EbIekl0aVK9X/YovBFoajSRpQN5XL7W9HaDeL
ZCDxxSlI63IfNzeiHjq8Y16auStspomMMV1bwmx/sxNJoS3naePjvh9+pKyipyR1
ZnCpUy/XTX37k0n1WYi5A01WNUsv4PfjVrbKjvanzp65g2n0qoM3Wkic+2XFKUXY
+S0mNJBtEiKoV5aHoTY1bbNRsqZj6BjV43XC1/f9aEcn4Qf6PeG7Cg2th7Vd3QST
i2+qaJsgC4He6n4Qs0J3HEfol+4LhYHTtCLlrB9CbyQWHwC+3IMmEeFkcdQe1QP5
R+xL0dXJ8SGF87leDFMNoXOnw0r4ks8avykDSlbrOCEzS8hULIBemW8YSdagK9Qq
8bPJs1IAK2GoWVpxVqyebyf7YftABRfppJ4FGMVTw61FkJa2pywleZSpWH3ssSnE
7sSbHqF9Q7GMj+Bp7IWHH1c6/OwMHg2t740eUxBXNmzj4hVY/wbeWQ3aEU38bfjm
sbrcHMwduxfcQwuxdfz9kxG0Vy5zNYG0VS5TXCjczSAbkZ8NMM1svw70n65hQh3w
JjuDvtrtKiCsUZwU+tdvd8cyqDNuRRTPr/lyOIvWSTrNaAtnbGsaHhA24UnRyIKq
+xqQBtJUuf0CLLrKwSa0sUQ+WrEKzKUARw6qJP+D0M1sg2FbpRjKycahIjGSmQKj
rKVXsJ35ngE0EzNqSQZsX2EXP2VvXpkuCeoyS3dYqz+GI/0rwsuF6kqediRKuN8O
r8Vbk9gAonBQDbgWV1SN/ld8jAxOXB7MlsODxceNArWMiYvvKCjbRCmko910FDB6
a1lVLSjOzxB+xcI0jUBM6MQV3tSmpMk/o6wrvv/AgD6x1nBqrfYQK8p6DPZbmpQO
uHAYT7saj2rf6t8F6qTnU85o+KXYb5J8TeZ/dpd+ZNu/6f7Gt0f7XfKQtrpg2kvU
+8wVukeIGcFGUJ+6yie8ylDfwORDIPsTFQXzzBM3qOmls3h7z9Ue2iGnK8N5gMSg
t2AobmqsIMHlHsO0n0I1nWbCpLj1Q1f5O/DdEotBWUS6Wty9vScCJuk6gEdWb4lI
ftOyOxIjbBhfzH3QWwdH8lCOI2l2M4nmBiGAVT3gl13BWKnFprOn11k+jhugHTKb
HK9YzY4+qKnEFewTUazEwZEeIMDRaP/QTaVf8np9WeLDL8YTWAJ9VKQej4K/2PCd
3zA6MjEk0F+Xe+Wisw0S9MW2T32W2/uM7IXig+vei95xubLCYmV9iwmgCyV7bE+k
gw5l58hDDKRkidUBXYR6e8anoqbDx3P1c+pcW6dp7rWsRUlQqgSBQKUwPnunhw6v
ufNoPLCJg5TiyJlqiuwI1o01QPZTtWkgqvpB+zEaXV/fQbJm7SlfAlI8ZA2uFr83
MGVClIe/8sHiGEfxDwwkyfzc7x9KqVZGGOPvgybB11NVkquPy2QIZHkPvAkZYz05
Scjll0l1qD+7akIbwB7VPiVvwjG16yPSF6qOYbWhGNXDYNOZ1xH5DvFSwedAfXx+
3H0JV7trHfBPyNMPiKb+4RjNSXPOZHEY38R2/naqBRMIA8B+EQc0BEOjuP3vd/KS
BkCI5zFAksM7qd2h4lqJX++pX9uJ4OQ4V6pC6b8etsEx4pJeCaXkqR37tx1dMONf
To9QklL9LN08w6t3Cuwg3Cc4JzNRA8MnsjN9xxOer/dM6a4MIUUr5qqEbxYTBNdK
5TakAoO0B6VHOXhPz7/sRUo/4qr5z1pMhnEuDliwDWfiW9aKX6ORcWzZbvepcjH9
hSjiEOhxzd8Em0ZPWnBw/TTeifFN2i8CddYTy7oNRS3xhdL9YOk7zSe44d36O/7M
PgqLCGJNcg1yn+rLeg3LOwh4Q1sftVY53AqwjlfMyQQ+KPUG9BBY5C9n7l94ASeM
9q1EUBjMJ88WF9o6UM7kvLuAzjPUgcBZcLhQQV6oxVlT69QYKqwZT2eepuZ5euSS
umcpI/kbW2K8BroBEOJuX6BNjfLdtR0+kWaTmwQ0r021UDJX39EsWh6ZG0daPRet
YQNjIyolun77UwOQtck3xkba2YVvnJQzfUMHqDu/WmH9YZ3/1E6Yif/7muhUQQ40
c8aICGkIeD6Cqt5J89xHXkLuZgZEm/cWeoQp4wm3Xw6upDZR9xyC+VTjRopsMGbM
1OHA5g6ikQGe6DG7vCuZTnw5BBtRnLvibbCikcH4DKx3tUSYEwx3HcrwBNslarSX
pv8ZxZ2jD5xKFb3jOZSDL5fY1muVBPiBKcXksdF78ECd0lYQUW+5XY6BRWEL81cc
jRFWuQYuZGRYTXHhPR5JWbMy3eB1ydlhX7akEVRYm06RVdPpWtqlFHLhOUOOv6q+
crY1eT9N+ivBV4AN2/r7Jpt1Wc5Co0I24xXI7Whkk0OkgucZD8GrC3ofh3ZvJEx8
iIox9HN7Kt6faV+cBYT5yQSK3XYcSTs0t8Rp2Qeza+EpQlByfobSV3aPtOUwV37O
h2nNKZZ+sCEBBIzM5JN89PV8lt0s1aicEUBzpUNwBFUbzRRdg1XjhZWDIRb0B5IH
46DnVY1DDEmeAbL68ibQDTKdwRiSeI5Crsdxfg9zJVIT8U98Jyg+sHQhBL+pefZS
UT7Gv6PZSBQH+cLd0MJMjKLGl8JLu+o6r7sNTI/1KqNDis7C60bamb2ODH5xe5zL
K8sN1ft7e4guhJolNZ1r/pahdhMrDTKzlebFcxwZp0qUWu8a1Ro6WlGLD45+WuxV
iEF7zXaiuo4fkr1rt/3q36W8NQ8E+fCWCaiNfYjrUZSff59RysLpuEXmQfkOhupD
I04tDo/YG5RN6k/gJW8kBG+2sVazOfPUwvk/G+TO0baMYUCys8SeUqLR9biRmDhS
058Yb5KoKiGmuNdnZ6HtEBp67koQ82+IN5ElFk5Yl4+KqXrxxvKCkEwFR6OstZCx
IzNFS+a6620VZxYwgpBofPorQ/v5LM2nxOvFvLTKuIuMRJA8l8WlGVAM4Z55Y6ay
A/qejD2Ce6SYruQN6CEACRzErQxJT8kUaD615xXUjiHTybsKl/hJCs8NvbULCwRL
zOoRJkBQhwSBFwFd7qtPd6qDYOnnF3hs8z5oDfOHgMmA/oC6KHF6MZ5GWfO+Es14
jB4B+gIDQJA5jyMLeoibPLsk5O1T5Tv/kObn3D4NY+Acza+ZBLNmZocOJOJouITN
+rUeaXSZahWKoX/G5rs8yIJXXsSgy+cGsTfvlHhOdjraiL0usAczbrbRLzxQTB7/
3YypHri1wP93lEEPi/jcZzGPYl4NacmfGEaIOlK0YfOk5OoGqL8cT5HC+MQ9oQ8e
Ae3x+Oql+kJMErbmY5YoSMNEI4XSvis7rBfIHr4OH09kRoz37rUsIsLN30mY8l3p
lLBnP1KwQHZG/pIkYQkFIEWZlOJIe5dV7FgsV2U6yLwelKLNADD0sDJ0TXcZtrgX
uo4/Vg3cG0RoaH6zAIMDjBC+fNAvMiGkCRWi6DgZev/2aeC96fOB9Vn9rXNJFsYu
muk0YQFdb3sc6eSQsZaKP0pTSBnjGDugzRul79JE30rM4iDKIDS2At56wprG3Scw
wLPidknzF2ZaQxcSOxxxo3tnC5LaJTQbwC+FI3slmPbGBdUZir0rc3aOaBbIThvs
JQqKjr8fvCJjbzdAA/sCLKDx6CQC4uhpTmPR+/D2vjzjct9afo3uoteRAe7tsfUK
aBoC7uCzDA6lawQ+rmqTDg+TQM86W/XmGJNZgvy8xykPgVdE4cVZwfp1J59PHqt7
X4zL4m+CHLhhaAwM3+KEcQ6/zrzPPwUKvLiKzmTEXHNPE2YWmPyMg853cBM0LEQi
Z3QZugNq6/Tfv7JNnVvT7+AkdJN7UE68Xc7lJLIzjLcb6C+VGKBGdKhkDBMTjmdR
doTbEDcEHTN015+O33xdIJC3xbwRV7lHM9vzuNFDjIyHxKFfFx7aMMbhY1okTV3p
c6P0s8tl8GCDVgkQVqiLQFDbf2WYUfqKp0Uw8KZm9FqUd6dtsgWQgmmcTU6lU3sF
+P3Mf4SwOAbk2jAeL+pjxAngUp9MDaISxIgsQ6tn/qypTZQc5c1qf+4A+OCJ+5zj
bg00K9uPY9vyspNvDfZYLzxPRV/JC2SwHHv7MthcofVXvJWCUMMgJDTHxmumWWWq
LqzaU4NPUB7EDfc3HhEjOyCfOkLrh/d3Riy2opH0kCAzUsPYJE6CkUGlqU2VCvua
kj5GZJMU/mAGvB7E7RGwReOOR2KOhipCwEtZzUwPRItvk+g1TvbJtwPgkio4fKFQ
Q+ZbD1v3ZZyZPdp+r3eHv21bUmhQd//KBHrycgzQcvj32+FXLhdOoAxa0gIWu91C
vsJzY1s/IRpD0+ACS4y+a+mzfBlvUDYi7Yse6Jj1Ri8M/DY+VSE9NQKV8fajiy/C
LVK29Jj/FY5oBOv4TmLt5YhyoomjO5nJI7HHVqAX7+OMQrklUgPnlYeXuWXuF6X/
jScNOGpAXJ41IxviMF4WOoJiWjoAgRPoyEMOouYZi5EJgl+N/DahiUlBS53XG00i
JH/KveM9Ys4k3wP3j/ipn96xdViFapPeYCUmD1vd5fdc3uisoVT/VJtfVqup7ZO4
xttJsoDx3B0SoKQsgnKqQrcx759m1r8HZi3tCDgh4q1UnvxrTbkecK2Ogsgj99nX
B6FvhXLd2gQIgJ053nZDOr2eLkYey1nqnvXEgVGn8WHG+fHvT3NSC4c5CGDsENZs
a1jEIK7tKQNVpgeSvL4C2hXHmbs63id8BLMXpcbYMjiTOF6kvGZrFh192abEw5Cs
9BRsynS616uN0r7SJ0jTQ6cbOJLgFMRd9Sz/hStEDfhncSNBk4FylVdgLPYn1Bn4
IH80d0o1E/sc69E3jd2YomMYiJ4BMzVhKk6veA7jb+tRxryh/opcWVvH0raFWQd6
cxg+TvterbSosGlhJ9E/3Wg9Pyd2XnQNnZ0TewDjo0mcXAOBrvbedJlm+tgqraSx
QzwS+a6HAZnmN09eBVwm+zMOTUsiLbtB0pWX7WtbMRTd/TEmE5Nf9t1UFWsJ/Oc6
WazzOcb6ehMJF6nRuTVF7cEgWcjawrXFT/FmZ8mN/UUr/CAXj9cLvKbnw75TiBsX
CkyBo1BdAl/PjdHG+CimdOHKrBgufGF7CkAsEtgJadTX+/SDNlhe4eakl0yIf7Ym
EzekG/1OLkuBCRlJA3r0UJlfxzx2pZbincPprUdyZcITTbDgazH6nuTFavfBcGv1
5TZpVgFAKuOPMfrtVSVGPXA5QiFP7MgbNix3dUTKQFoIP0EdvDeGWD3PGRTc6tS7
flp5xEj0lXPMigywLxKTgnVLqqSTbzNQli2zn+owjDuduBIhUDQpUb9upZRoh7IO
x4JKBkt3KmBr8LbX3yiCRrAJLcNEN43sXvE/fDpPduKtnAjGdUlaE4obaiSqz54i
bKw6Apgj0z8quoGtmkZ8ndFOzY8FmI3122sUemNIHkAhVpgIHeWqbOiu/3rXt/QI
JAHOkPk3pYBuWL6aacWlmSH4f3De4q9T8rKhds8iEwYOTByNz8I+RtpsSu3OMKnE
imszUHf0Ozubf/sqSPvkFjass2uZEATguigi7vr01PbHnUq2dh0QcVGtxGkbuMdF
vIlL4+EQhJynTWNY1oyQ+WRxJLKtg6UejeJHtUp1xCTVReq9Sx4Rrzr7zP9YtxN0
YI3TWiyI0SLBncMlmMdt+I6kvQf5ExdfIhJ/2MOXkUOyNyRyTyB5hFBX9uERzC9i
Moy3q6RF5HYkhGiLjbPKYGNoi6VN31L6zCYMRsJQIoDueT4JXne8EEe7nbsga8KJ
sYTJQHUdkSp1etbxvXJUFDM+J+Sct4F4rrrnjkjnbuamoMnbmEqC7gdc7RzUD8EJ
XvxuMTeygSU7IYcZIZajIWIZMtvMeIgFYE7CUTIxyoAumsQTLxW3Ix4p/R1XdgRt
cQGRvuz5rJVudknJYHFrRfYVJ2WZ2oFFRYiJpN50cKj2ZxcSzpsjdSxy6vFU0gTH
088xDIpss3FNKdRxtYWHoVNFiQ/vLpCN/y9h5og0Q9s2QfcPw/W2D3Av3tz4Xjs4
tcBGP3s1Q5oA3wxEZ6CBB/vzDOoDeQtaAgvxn/KUKgXJm7/eUIFwAd5W6YtkrWxi
wN11cIFVcDskkF17933yMcAu5KEnBrpXvKB0BueYGDXKbC6zPsM7j2cuYWp2ZrbO
/IrAgEnCjGrA2s1brRkWntdvIKsO82STa03+SRg52W2RViaqn5MopLMJMbLwzN0h
I5uJ84z88/2PXTv7rCGDGzExv09G0jenxrQ9IN3/f7mcYFtCriJy7ivEODvyT9E/
oJT1Z5gKnQG4TObyhH2EFC26HuKpXdpuZxhpgEdagr23H4hZWc/bOq5xOznNSbFv
6XCQiEhpMwDdfOq8wOC5X9EDA7zXw0MY+UqfV6Egphm2mTw8i/7lUxGinTRjpP9j
kh8zGvuB/wlxuX1OG9T3X++mTyMCIkNlAt4pWdUj9CHa4AoaYtwlG6b8ylFqXySj
kUWpMGR7zpDbFcaU+IJSQBlwfdQFejRbbws3h7MAYsCO5px41Oblqu6K4/Q5pCXn
htLUjRYvH5eOyFnPMFr5tFOmfqN1q3jj1P2Mn1qxaJn6Q4mdSWAoVe+LjCrjOeH8
ZNjQv5EsipghMMW6wuyE8W1zPthBKP77PCo9PjKUZOdFOzFyc3rxRS56kgxNH8yb
0rmurXcgrdR7HZdgbf1fHs2cBDAFVETCM7UNKJ8qxZZsaLwPbEsfhriYQjxXNJC5
EMrLMq7f1i4HT3U3rZj3BhoY2iOulnEqUiAP1xvPmgYDesArJxhjaZYocXqpaUuX
Cr8opJrFV4RvlLXqsH/X7arUCUgA7tlddHN/HsKann7Y78WsCpFbm36/R8qmWNgL
YV/p33S7vwddmYprhFahMrQv1kK152L/laAOz6THewpstUt4+Q9yWrbT3I6yP4jN
YKcqL7zGFU/jJOOh5CwwTqGlqbf73uDhG/VgYlfyHqE2maf3HwpuSwAbVe/DGdwo
EOVqz8mARCsSxngUZ5jD/CK3Gi1UwJJTw6/bD1HiI9H6EOs6doFTgjYBJmvtey8j
yBgG0VBC3vWZfaOPE6y7ll/t9xaAFPcTwo5LxNaCRPUOG6dKvJZfrujCw2H4TONS
mKiKhBp1515S1tvm31oYF8+j5ayIjNPJPtkEblyHoHB5X9aGoLbqE/IJSvAVVDWa
++YYbEFXVyrJVS8p2CqSPJmzZTzDHlTVvj+ob/pW0kKNtWz+khL/oZfsdayuHbDz
iU+RiNV2lXdl8/6n83yAxOoYddPKhQqJgV8ioQ1fryQr4yT5U3dQ1582ckj6oXhH
MmpRqVYJ+6jlcgOu88W+L8o1/OIQH/dI0B5QII6LZdYHnY4fGeCXNi6FRWrnEP6r
xClJFBpDzdnlptvqSzUiVFnDUJeh4w8GWkO7FDmvonsxKR6jFjFuHNnA52ldpFmM
hs6en3DMz+H98jrVu2ed5EmH244bipWbFsqUxJTrPQ5klJn6sXNMCHKDihtmEn4r
svJCdjPznQP+5AL7c+nEdg/e2vBOSAc7Vdb3IDcl2HZlxhW6R9lDix+ZwDUG+6PB
0xJqf6KwfRHhn64CGIZy7b13/8vOVwwPOJsKnbZo+dyy1yCgYpvTwEe82FSwWozd
lMMquu1jLJM9ZdAmV5L6Qr4zKSNeFhaI4gZR8e0fORTncVPLAuRIsm0fXJBEoPq0
iTxn6nCO4c//zfhbcTwIcOiX65WJU/AmWp2NXsO8h+w9CqPtUJzgDNKTaKCBnsX1
MLqINhx//UuN9w+Vk4dc5qYbWKQz+2qzkS0YoxJNIBN9qdnUcnJVGIdTV6mL8J+k
y23Nk59MyoCQbMFIW6tR3Pew0cZRwYGKgZyb/6AGBUwde/fmB1NI3up55FOtLKKI
3TAmRm40IRT7x4DutN4o5czV67tEF/8upcJAfE9SWro0WSmQz9XxfEPcAHHTT1ca
GUGRJdDiPrcu7WNSIWf5LaMeKDU2/pyv9j8QSc+CPT4ooc0OemruLIKQt8Ejik7c
4JT1RvdujTe7IYgOGSchuUKYa1DskKSIWgqOOyQuNxi97FkCHWbKod7gZ4zc+JJO
+CMWNcMo3J8lFrG1LixcUU9AgXOJFTJMOC5E35GseNL3oXw0WZ+3RgqoVY43n8oV
xa+yYbMlqA07uDUT1dmHAgbtiZC/P6zZjw+HLzLHGUKeTg0iEnSxiCY2FonahuXh
siWZslXT8+KeZhk97lpRBsiupSmQ0TC1YNN0EIbgRe5b1YFhlYdxrY4zR6vlb3wl
iKU2/cNE06QGkPbB9sBsqRPdXAdy5bzyUMUH3pYPkhqaP2crkg9dyfgLhXnZC5RQ
tZGtx6qTICvtxdy11OaCn/icjk139O4c7zxU0YuUHOhno15TAKNpH4C7REeDyzX6
KZZpsPj5WGN1ud3h7430EMg9tP6+/Ts/mkgyKmpxl0zcqqH1nuH9jpkvqqdcp4ad
sIaXDcXWsh4LWKAdCiKLy79INufO+o27fa6fcI2/Wj1jf8/BFDuOn3r+llMSyHW4
H9RiYH7YiMLuUqODp4wr00KhQejZT7f7JxNjQwx+j9JvffoqeiiJkvUFvd4S/Gxa
0vQ6b8vzDikLsSKpWMDiRGKf+1NBrfCOIRQkMiPPBVDoLDs9qHxzOpoy1LSAX+WM
t1azTgFiFsk3HQ6upIPOplteobLE70IG1Nevt2CbZtNv5tWMHZm+84m0eVqBq4Yb
JqGReRvUZQTBHQIpZgdy/tZM+cF8RUcvtdBKFJZ4lt6/X6Uov/Wj6V9sLw+NWgD+
4qHSKIzOfxzJCsnYmxBvTr455V2dvQG5199wYBEoBnj4XzzbVJuMkrhFjju/0nGd
nvFPaiyPibYGODg6kDYQbJM91ITcAxpJJqpc/60gQCr35INya9misFa2aGmJjF7m
7RZUW4I3Hx5gdJMe74oHPQ/B0irF7sTAyFfef2oN2mJj4j5GgU+pEg/l7hoJwvw4
sY7NMhCgBCCR4Dt08jyh7boeajyqW7dEv9nayYKurs3MfkSjxSPl5uJ0m9/fEgy5
Mkz2hO51ouuno9Il7NheEbWr7NreoSwUEC21O6RI6eTBtHTDU9oo8VFCbk++h227
xvaq5XNIQZ1suHQeZ/1EhhVstz2+BYUUxTmJy1T5RGmV015j+aguQetWDTtBW079
HLDQpHYZAuyA1N60nR84owqAsA5YXtSSBXekj1dB/c8BgBcPOV8tdCX+hrmMa8Sk
hGJDFwZPF5fynWiiylRUpfhFAgtQ+L3K2TGFS/VF1/Qud/SMaF9z7HaZkTM2YoT/
vwmp/Nm7z4GEIvddXGhJOor/R5Y8C7d8NYy8Kb4OVMzE7A2+cF+FPtpirKo79c5q
K9P+a7TXhHLsHlAo2XIt5VK5ChPrLZFT3zueo4HRk/n6NfXK0QzrH9lsTYQqhdb6
x4Vc8d3dXChbpx3MGZ9YcVzxk5VkyiSEzg/wlu/jpOMfqD2hQ8Q0Nzpd67QbJTeG
LrjyveD0boWewRjaKPDdftUYKtMBvup62AbC8cH/egzY29zkm+wIEkG9gzsAgQNL
u64Z+sUFfua2ZW7GtX1d40BsieFPjooScTuISeZtRpW0g3nJ50iYtkbrSqm2angC
N6rsygOd9kdrJ1lqR1EM0k5qZH5aMN7SRPOyzCSFKdT82VCwEISqQax24+IppWxk
hZ5NfszRcmF1TtquirP/0R+S1/Vj2ANSXzfedytZr5x1lOWywRGqHGKw1+k0gGU2
qgJyTE0XFVrDz938TaxXA73WG5zydKjszRBfd5ihl5+auLi0dcn3ceUVy302w+pQ
71TnxbKinyWSMDoyQANNX/xdbNkRtmsj796vxbXovIiK5Ayha1LoFNc0DJCI9yDH
HtXhenvmIdMaPXW53/HcqYpMX6yncSgv6M1Yn7x4KZKYAofjqCluBct4JcylZ8Qv
4C1zykOmwA8ldlXXq1QLww/S5ObCtzQC7FTtjkGPfILXvdmWYUJ/AAbpico8TGx9
738aZoxHdK24jLH8CrvM/nnxKZ4NPdgSXWAiMnlPGLrfPGdAYNDNm00PSJUbfSdC
JBcIQTNHSpODDkU0Bg7enaOHH2AQFclA9CwZpYjOBqm3UnE8uzzf2SR1VhRo9Sut
YfruM+HJkSZrTRbGTaS0AEoSiYR6/uyIsFkDWLsaG1ToKdOlRPyPHI1kosC1OcqL
UnQBytQ9QnBjKOwUT/sGpJVWQrrDF0SUjZsDVmdTj3tt30VQYaoMfv7UvkFmY7+5
T5iUyGVPkPHVh8gUaI/HwbVqw8x75MV8RA3dVKFOYuXlhfRKbr6mCEdwh1pLXd3J
n/ap8gtcf4vz1gauOZW0Of/Aju4lXHXwHRNucZ11CHD8QaMi0E7cnQ1eFYqW5fZO
WoUmliUygnBUa+i0T3twmYDgoN/cMWoC2t02KbFW/qU2JsaPLgQP19R1UkBa222L
DVf1pZCp28FiONq9c41gdoA/1RXj39bgF7rtJvAqR3/5mFQy4Z6XeVDuYp9HlIlR
6tpfX1LbL9Hbudgicp0vhnnmVDejUWLlblqTpijJQXDL/2Tae3sSKm9XZzPiSOsi
KTxcDPorbYNydIfnul7SfIZsu1Kxu7w4mXif3r+kSq9975U+dfP8dtO1uX+b6w/c
22c2n0vXCrPZRCSSld2YKZ5ifnUst6vDNFrwU4mHSRBfpis7GXSlx7XUOYEOwWGK
2VyiQjKyQxIz974rSG1h2EdSyG5kfRn4f7Jdc8VIdAH9zRslYCPhuwsSCSzrYvQU
WqtyG/7VruCve/xDXMaixwQf1JH7DN7fDBrBJvMxxdFqYcF2PVYJBa91xVHNw3VE
a89bAAAdkUkmExGKmVScpvrrSJSRiFm7ebNm5aQJrnmtqBH9fds1Ls178y3fLi4o
dkER6UJYn8lcI5kiLdQNh4i7yd/IDWTNgAaZp84axtID6ifAzwxHP+/hxd1IVTP6
KDIhCWTIjpaVu04hKOCtVdJVFhRUnqHYNQ9ACWtJI3jSk/K4JBmVGpldkfou2VIl
dLQEvAZIYMS4WOZdsZP60uZ38uvVTJc9J+RiZOfdupi/vQK6zknAt6IUMBCUYgif
34tFMBoyxnyfK7NOrSDHzRBn4+9Dis9qKy4c8vmBVT0a+Y5OGoNFUINVg9nANDz+
h2/ZYym07wyItLE7UXWdK/+VTuAe6ZeZXFOnGMQgtk6+bM6bVrvi6mcIkwNkCSa3
YRLjW7T6T/le5dxVqRRAZ3Y5ODneAyqh3aGzLhY1lZqoamNee/3W0uOhNLB26oIO
lQa4NVeqjeDSh/agw8TtUYqkYdDK1TzrRm8hLn7DWk36qRJ0W0kpQV4c3AitUYVX
QUgo03/YxosX1A1eph8lNR9b6mnoFORt3nFC1XVH1pu4ZlkvFBQaRUi0yD31ANCx
chMNimSCfzMGxqpr9SSh4z5hRKmQW1u3pqzOh+oR5SPKXtO8LSC+cTwupAn05UpO
wmjOXNfV6xeVLQv+hGC+dSrzqux7KRDoCSa8Yb1xT3qE0bz3ADEYJ4tY9rmfaEJM
v7GnOj9OuHmwwY1BTP7PouAz80TZO2tYru3BVbiYB/UdWrwpbmsK5/CahT6SaDWI
9RrwmKa8k3I5hpsY2jWi6oxD9J8gIp/+9chHUKOFRBtMj43RYQOVZOfU1sgGrkZZ
5VUNRMtERYjJ8Z/vDnlw3KYkyGQ9EK7AWb5Bs9bNQaYcBwEbuu50k88fSz3xM0/9
5i19eFfbEph5EK/LDbgLGpQrRmt5KNM0kzLM+99cJYdwZdQGOLuKyGa1/zVSrYGu
Qcn8iNpdgDJJIp8suyfeH/M99985ETtu77XEyOyZaeqTP6bVAMlpXcZ0dT1LRHsq
D3iRlvc8nufvn74ps/wEbQaIKhw2wHL6Gp0uzeEQMN19JFSerbH47csYA2+yKriF
CkFsCixAcE5EiLEw3wzkyir4L8sk5s+2L3PhW+6T9/98VPA3pnBD6Nt4B/qLqWbA
Efc2yHrSpSwS/XqxeSYw8lTxLtWS72FDAIxVxG4qzFT+it+CbW5aggJPL2pqA/2k
WHzZbiqY5p0AJVnNifWycBObNgn6ErLBm5JFmuLsOL97A9769m4tKHaMSRzs6gcm
KKH7sBJFYnrqCxZUIBEL4CnMrFyXijTTba9EEq4i8Cqp/hUmXBlQ2XrRRBO+G7+X
6tHsBJNeeDKwY0xgCbMH/xAy3qQ6Cqontd7wx+9ZUa2MnYE243vsF7IKC2IDaBkK
B5LefEoXb0P4yNPKpIpeJDUOXYPitvv2jC0cO47kU9VFjnc4Ph31J+OSZOyiCEvl
O+uDCMxeP+0euG9bzEf/i77t9YygBRjaD4iPi3oz4OtIjfeZxlCoG4+Gd6n00keC
1zZY9x35yLMzOtQBvBWsjybBrrQSqZWnmtehu4P6je9jmJHeZot5cvr6dUqFi81E
RiDjoUWIoGOn0zJQrzIn8pY+AcgbFWodAjIzeKCgrsUeDkDet8Bx6liJ0AnKYKLY
nWAM4H5ciyVyR0gqX7b+eDyFX28686/OKr9qwQt0pDnL+d5m/5M2+1nG3o+vHWoV
/oApjqnqR33kA28OESl3igTsFaoDHuCXfOCebynnW0Tb+ZEf4pJVXsCqTPvNW+vv
dMp5ox5U07DJ4F3705u7Jqjzf5ld8ipCjcKyiIGV9VbzlCg5mlJfuVM8viC2qSwV
oDTS6fEgCMNGPbse73p1Lci51FC2tSw1mQygDcyiupMmmczOsd8h3pj5/XryoXx/
OlICURG/RW7igWqLg5uGZvD4UXdrlibAhdLrVL2WqgA1EvRDidv8DUZadB9WW2Yx
XcByBUeiZr1xDWgS41tGmW/yXt8cTdZidSIGVLeEkCn2i9HIUoY9ugJRUkeHkaOQ
ObvvinltCRJix7Bgo9XHTAQXq81u+cBjZODcRKWxBqGmwzInA9A21RWP/ZFYZDNg
fBepqXks0GZuCC09mijHIRFhvY5o8XlaQyMsk8IJwoqCDMk2yVBr9l8oOOmsxTLP
axB5SkBzgTxZXwRWXuoyy4nzxkOV6zRHI7TqVu/Itr1CMvPCcIGJi6CC5REKf9QK
h1WvBFiF+mUc6QhccGJ6f1Bgf4KO6ZFY9H0dhZgU5xAZsMVaLCPVk3pLiMNfiu+F
ohNjCsl23vmfl/jgYXk5cEtohna56+4v7qGFmSqzgW7cBC3+EJqWYhK/KPCZacFz
Iw+iD10Y3bUE/vS6qHEDlU7WyC7MYW2XIXtJBwkaQXH+5BK0IbxkFlHEVnUh4Jxu
G38BASOviL1Cwi9UmnISsYdo4McW2L5EqElCndkJJZLDaTlEnT5zUfeDNLARTYPd
rZkP2KvvJc+JXzXea9soCruhSGzrU4uYwjziS3PkmiDUnlEtZkDfrI3bDgyAmo3U
UvaTnKKNkLA8gQnk4pLrOeSOtHWxXDC8BayjkXtkKgLIPCUu2Ro+b898MoO90GIO
91BEMV/DB34AS/pNX0xlyZfkWO5TvJ8aAFEH162hGgZ0/WMeDYCTiI1LqGEph3iE
EgcUvLSDLCLj1XubkxeXpPG/NlwuMPzvBVwQt/uuofQmJiZXqD0YxbiadhMRvE8W
GF2gLRwQLHm/QKUCR/432LNfo8yKiONeuataUFcNdHJAySTgOf21IF9VyicLkWbz
3gHl3TwXKMhq3lhzLDS8xRWUjYPinO93VuZMlbRcqYV8mkwTXIPYm+gkbUyLUQii
v46X6PERb/kQEKrdQs8bnVOW8icJ/x/cerpvOYicIfg0lzGmEDwgY8LzFug00cW4
IAaBaKNMR664E5Zoa8IEWR72GDRSHI5Zucy4RK7UqvKLjAvxEcPJ3qyY9tHwKjuX
2pwgGVWDSmGttGtexFFcZfq6sy1gVG+yFzSLGalwFoyHSkLBnyYE4XFk7V8CPzgP
uvYLH7datURLc1Wi62HlCjIbankKrPvjPUzp8uA43+0l2LjrMNaa5kl+KBNHC0tB
N1RrSqygjI2pwOerQHRoEUlhOEFFPwYigLu5I+Hom2YAPR/uB00dN0mEp/F28u+a
Sopr91brVWAL7UWgiKMEetOOdAxrvdhkjeoDlL9AY4W2P9LfGFZNOdBAN+TrEZ4k
rMAS87XF9InissFvbbhAVISDCRlanNLnao07gtuofTMfrFaVCHwd2QfcY6046L4V
vrlCTl3hAMMY/76BBWOukJ2j6pIYp/rxqls8f8zXkFGX+Pm/LqyjCaQHy02hbJnA
RdYXkpHBbWk3YRIYl67spzK8aXds7MULnNPcdIQdotVwg0FE3oCAkN1pVeIR4sYP
tWFmrKlN+efj/Ltrm4KRerTjcuoi0ZkVq2mBt63cokF5/NuryxEJooqe2yd07Z7I
Sbs0gKN5w3jk5a8rxJvWx8BWMZif/RCykorbFo3DHjbqhlVKLADpgv1S4ekRbtP3
GekNEZQZsHDRalmzRyLN1a36ZNpqqOO+K0h3LbiET1QpCtAFX6Zwh39yWaq/1lEm
HdrI84L4SvYFRjg8ZmLWwuJ765FwVcs7npnc3V5a2I7GWQTXUD4d1vYm3DUM2T6C
ucuDT8S1PmUToaXY0je7lTWQqRJRHPQCfwMKh4UG1D+jh/GLpuyqtRPJa1YOV2xq
81eLf7U7IBm+xmDuyyNiF3ifq3TC7LBczfblYRCYs2PV/658ZcYCiOhQ5PydD1Yb
pQKrvAVZErnCdKatGIU3RS8YwsycOCWOuueP3soMmU1sLVr9d4P/gWJeHn3BAs1I
7ssYpdQ0Y3dNsN2FSuMbysk5t92cPvRPWSf/qvhPiutuEC+mJz2FmH/nrnhiZ+Of
qp4duuyuy16mrj1VXh6rmNXWGph2dyMHIM7VlKXErj0ShgPJbpB4hA6ZcDhmEg+1
sEhAmwteeB4I3zmG3VhHts1IFRNQLwUs0aLKcCrLqXGSeyGPy2BC3k2n22qZ3Rw+
le4abhq0tkJz8M5xqIx9cV+2Awf/3W9Isw6LgAensOcKMiRTeOG3kYSFyydCreUO
czPp14Qn866DC3bLxtktQbzCi2GehTgMTVGDmpjGbwIZ+UAZSvwyJN3JU8YDtGPH
n1x4dyaviyMMR6RRSjVoAieYtTThlHTlL+J2+HJJa08KF9ziaOt1cnArF39wFqZl
J6yeNnslHKKGeKBEiQiWvas8IJIGBvr1pEP8SBOKAspKOSfWJ/BCiCgyOH0vhb2g
oBdWonW1sRh7bRg9++qLSBRKeaC4nx4l3mixTGEWkkCl/IAEA0Yz0a3kHY3Ei694
5YcaqTzCu6vwRQQU9fAtcWwUMa+C00keM1Sm+cv2SKKsK3tmKvH7MMSPYPrg51eu
d0go0AwlFX4nedRiKR3PFGtQxEJ2d0az3LQxsoOI6BqX1J3vNSE+YU1UsJat2PlP
KdFt2+SxF9roISbZL6hClyH8tQM+nEq0teefSfzUeHPhPy14yhQnXa+8cpM0ewam
vjKXoK0NMcM1a490kuWngyBVLawKTNWMHN8mUYnZESIX3k+3b1igcrhqzwV+Wz3K
kVTKwX/yMntJx4r+iFJCLAtpY03Pgn0yxmW5MAXVSQyHCwMJlQlDmhjN66ise7+j
6W5Oq8eDpQ9xckc3TniaPVupznoJaCP8fdg0o9WQPvkut7YQKTlkIAL8JJzXl6Et
VfKy4eG9JHG0PKfgcvdl4qH8GrxCMrt/Vni8EzlfABPigrpE/Rm1PLVMNjqHY6Cn
c3TDa5NHa6V1P8Cr2Z2U6yEzxh60gk+O9wHsoyeqAYIhtOpEGxmFV0D09E/CLqGh
ub9bMT1zIYiWgdK4UB08/g==
`protect end_protected