`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 3984 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/59UwEX+aE7FohaWu0/8IpTj7mav863zUNIsgIH2BWb
Abd9opeuBjbGF/waQMI2vMJTwD1ie1YueHc3nSNpEh4OXp8P5ybZFY89uyGz3ztU
W1EsuUnchJoQgbHZ/sLbgtGRgsrAFn+ZoIeGN1d6RAF2wAESJmYP8zw+p00RvjZ5
pBGEHX7wooDexzkaqKS5GyydNoJwsMhyVLIIOuwrtp6N64vnovhXbCPrA7yFqJ71
Wj/CTCAh5E0PJ+L1QZEgXoRUsOANGjbVJezcgslN//qoxN6Ntrb+dx3voDGE5vHd
ZPpeJGsBXf8hZJa9D3nMLzUOmwFiyRQJJPId7Secq/CCiYfYcKkGLjncfcOCGxH+
c94dUN4KbsjgSY68TQ3jHS0eUVJ8zCnFWXHLoz/npSDU1PnjAtges1wqrXmLMyEL
tIrVdWzsA7i0yUodUjBGU/VPiPybzOWuAWFsMWlcFZ/rZfmbxs23BdWLbxSW4JpO
XqCTLjtu3D/UOg5QzrTMIqNn+yzCKuJDZA4IJ39zgwsBcGwU6tZRSAdI3s3VnZiV
LPzMa2GwkJu8vYfNEEmwlEGkgBVxfx2RvcgkSF5nb8Jj0ajXk/QE9zbYGrMlnzpv
7BzamBcrfyyQsTWcuGpFV1PJVMBDJP6jvDchNXM4UKgPvqWtPPpdwY4lY/xb4pCH
8oCv377nqiQrvQiHqcc28OT5kQKSKVIkN57JUKBZwpVfW48CX6RWIwmf/O0sn8Kk
6IEF3aPf5P5EMxRKSop8UjH8XxXo1a9AIGTTEFulSlXko17h9nx9ez+bzg0eg0Za
zqqEwR94fiRxChbyuKWkTsWBQvRFwq/PVUDZQo6RSRAwuFGrsvrrjfzF99MHHN5U
cklnvPP4wglRHnU4o3C4UCyONd78b9tflxYp0ANxHvSczDxR2bEB2dS3vPiGVtWP
8eRC8iKkq2TUMwlnYFLn8IbkzIQ8M5Vzj7PHihz57/eBhCZN7f0U9SR/zMApAGm5
RUWSQnkoSU+HvyTzJLakKkD92DCmQqgSeUAmGFwmnkJOmvLCGcX/MI4ET3g1+gxc
WTksRJ8J7Fnnq77yu72we59+DXExlk894pZWWSOLqW5Lxt0PryMruyDfGo1+nCGX
UpaCR0glPHmOFuT2nMs5CwLAKajfamRzzsVJ5IT+IVdt2HAvcH7W5XQkqg+t6JC5
z8WjB/dEogk6SYr2FM1igzpOYA0u16sR3QEE7IMPGRlUwT3zntrA57JNWIHvmnSp
AmLZLTHUZEUJDNc+wdNVa8sWcAFCqsE0Yf2chZhQPyRvaiaHBG8gor9EZ8ORBwov
aCa/PDv9XUvXPMEee55rZtyvOrNiwWjv82ybTj6v4F/2n8bCDLz8r9OtSMDv0Xmz
TcJx1C6vCLbjE8Xo3NvFqN0TY/zb4NgZTcVdmM79MFXnDow5+hJiBVqN3ct5Tg3o
itXsS8ijoq1Tbx25hgxQuoeSy5cAnSj8+R8K+zybPziKYTsrEyWwPf0VAQlSL725
EXq6FfJi4zmavMQQPbcIwDShwlN8mJ0wOC7kZs64iResJRleMBaZb9MNX+VjFJ8W
SULOvQaCtp4Tr/yciihBpw5h3UgATcmupa6Y0xXblsmL4mLaEgOCjJFcZUfKWIVw
ylWoTzo8m1B2WpCZPEtZOOnl3svOWdaUTPxkaeRocfzbEVMYEsBe63HPR6Bkksc4
L9W7RJUZmvpDxWaUQ8iDHG3vYdPuaUoF8poFurnoatcmNd7lEqG2tYqi8RrXqZnl
+xq4Mdx0QNNdIFnAPrl2seNGBQ28+d0N2bWckQQHk4FQ1hbv+A8oGNkk8wyvUnvP
HQgQcXnSfZn28i5P6+ZsSyYmI+ePJyBkC1xrduOvtKDfg+G6wUB4vCiogq466zGh
vFfNmjrXXBJYSjLsVkn9QDt9D/2gn4LVsD91gYT9kXzuE2opSIR8QeZTy3Ib1hIm
caElju5sfjahCMpjDSJUDsvFciLj8aJVXQmUb5cv6irM4W3hFo2IO4l3VAe11GDc
EzqVNA27i2S35VFd4hjHyIciyZ6gxqQk9wk8/sHrrminu7k7ClHNnYv4qUJv7jzz
gMh3sdol7O9puDMiap52ptMNiiOlacFfJOzzwMgK8xH9ajX3snJaW6zhIrcfG/ot
yg5EyvMLXQ8WiuL3wYVPPr6i3oYjBSTsvsUdj6CugGv6iDWH9mHtoW0D6vSl8RKl
0l2KYVBa+0x3g2IPxTxBmC0L2CCtg1iFpDT9G5pkyMVCH8dcr+waDvskEWvMtikE
yHwyqwsE73gpjDs4BsDDzszP8ZbU9Dynwye1il55+U9wHeVZ0fmjFcc7GqmKoPt1
6gpW25zanYIWM5D2GokLUjYWtUv7PAcwLHGbB97pz39MgMo4lwyJXMtO+M6CZ/Wr
70cnEz9UM9xuu3s5QuvHTIvPa6cC8HyE6anWS8NsH4e90WZx/9VDk9D0bM/rlehs
d0+i+N/5c7q9OUd4jEwUKzVx3Ay9hrLkpIN47goSamGqDFCUt5KDQOWMwC6THg51
JzkMYe5VZAWwkgzd/LBCDYSMkFP3wKFDMDSI7zRGkEeJyYWpq+dNTxKyf/KM7Utm
n8gyk0fqjs4Yr+TuNWofJ/qrV98idHi/rik/3JSyP5z+DkcrpPpXiN1D8B5VbgTm
sIOYlrPEIPJAgY1Nm400IdMb7bpYQ+rrF/+xPxjvDT45RrtW032zv26aDM1wm+UQ
vFCl9VLo+PR3TLLf8TXpePSnHH7UF9huZ6kdvHARznOp+fgzWOV2BKFM9aDMH9RA
oiZSjwxbBhcudjpPHXhZFAv6nQXvc9PRZA3WT9nfH27fhOtPWl672oa3Kmda02g5
e5wvfQgFN9knuqie0J5R3RDP33Arx91GtbGDYhiOvle5QoJzyB2yYYmWSaykHlIM
FS2EJrkJ8m6ypqWGcrrqj0xixARGOmnZyUzd1gNu2VoD7tO5PDO3mgPiVrjxS/j0
d3Fm6CcvdBaUY/d4V7Frecq7M3qD6NcRl0qNSMJz84KTO7f8yPBiiHKWlkLncRpM
UOLvJAd0I/g3ZaKN22mPu3WAmmkVvR62tRbS5SpPhW6rstTRxAvXzr3h4phsIW8m
4uacga6l8412ZaT5/Cn3JSv9YYYcH+Nezy/q77DCxTAzu8E/4Nxh/q0LYaMnjhYI
aBaucfn2s9PVRw4+skdYmM39iVuDNkLRqoMVYgH3jMBUODQBVY7lWZTJHKFOsbat
K0tjMYu55DVCQFenqsLBXcQ6N4KcGg4xdxAcu9qBbkwLAgdG4V80ExxNZ2Kyhy+5
dT+VFPekUUp3KlVWxsL8EesQCfF3fSPaigaxBrOVfB3pKzuuKqzcKAYoHnI+hrlf
czrUGtraONC4RSu+3TTW27623OYYK+NUmzaPVTHxMPj+6gmWN+/7nngcfexR1XlN
P97h544LuogSYEG4QR+A8dEOZczeOrQoF46KkrySm5mJbqxgRx7/JPutH+Hoa8y7
0hfJ/KL/r9NBvbhzTMLQNhFS+S53bqkyTuz/ZkyTMXLYlAcvSWObJBtCNQOSpY4q
FzNjfF6R8VgT76201pXPfZR84WNuMJ9hqg6E+UsvsKB18qF+rrMmQlAg0WpD8Bgr
KeRYGKAvcoGaYmqExvMgjnlwHHspU2U5KgCMBgKfmVlxfBs4My5+r1+L2ZnSWin5
TS+wDGuNlnhIa4lATS/xZLSpXkEESB0bP8zdDSJBlIS54duQmfMLfbERDmGLkR/b
Q9/tRgWBlQrBqO1sGzQCPkhbL8pGBsNiXJvjDj0fk6ebbtPvF8gqMQum3fu2eUNz
Qg0mV1p03emDPe8ImFelda4fXUZz92/zVIp2p+EwROtH34NrAQNf88JkJvNmynqv
vI0KSwTtKgEb72E3CbMbudj0vwV20uUrBbfecDBWgIAvF/2xAqNO25eP4sR2QziM
LMt0DArGdJmx9P8IgMfKipcBw+sS0sbFDsX0PypSVrcnEj+wnSLtUtMq+ueh3VCv
NGZkYn/n2lB1alNlEj8mvSJleRLP33BUdFKluAew+8HEc+W2tXSiqcsezKSZRJbC
9Q3MRoHrmTRO9DjjSg5quL1snk+hd1hKbVnIoruhJ2tR5DFMpOsduvMU2mNi7duM
SzTaxtRIM6bz/wQ/UTH/0zwER+Ojq58tZAfBycoJ/Pq4Bx8nymRxW71gHtxQqDb2
GYk6Q5axZeWv5NM6sdumcOA+uDQBAoe6H9c7fYCYIOYrT0YHNa2FdI6wGaLraxas
EgZVm1aqNVCK8SE3Ao5nmIKZjALckdUV3/fmnxhqHyAHDp1QgbyEkQPCyOtJDrSq
lCtyLKvwHPsq1tGQ6kA39MBQ5z3scjKV6RxPgu3sGLdcHZFsmiThX0ovxPG41guK
BQH7ICd+hMa/rL0jcyyxyW3NksFoYNfFyWNO6+S7KA+bBPCZCryB5t/90seDHD4c
SrvnrBb9a1HmOiciOzG21rHb4jx87lLExgStgufx3FciJwe6tKHRgr3HK7lC7U3Q
BQgO3znyM9qxijmn/dGRDmDNp1gtlBJyF97R2TiTMMH6X7z8et1bqHu+KAMraA71
yAi8coDM/jneqjlXU4XmLc3FwAZzzdvG+nkDaYQKOKo1GhX1mW2FzqQ7w0r+h4Tb
Oi+tsfdCM+lLFfIxalrqg6XNRgeoVxg+wGW5TxPUIBNmKIQX4shY5GD/y8lBwemf
ysMcjaQm1u2ZWXbvP9quOR6/m1d2TxQrDP4JGe0Fe41A7b15kwozdYWeHxmUsmkS
W4Ao68BVB5628z8d2bWggwqkOceQvOYNzb9cXtB9/xePOEwAiJeZh026KVQgkBvD
4Mj/ggYrB3opCuF/SGaeDf+zxChJcK6eVCSQPuYtbh6l5RFVq7BP/Qu/+96G82r6
NbEp/KEJjpoGm5Z1a5/kdpSWyj4ETuqTRm4gjSXevFuZ5yNODy3FP6y3lNF/csV1
Qt09oAFnkBRgpAROxT/n97zlIN8NpKZa1+xNYKkJF6yHR1BESw8MAhIFW2m7CWZn
iPjTwx8Sf4DrGEtITR6DAFs2it9x4EFfXIOOePx7aMhnSFCKAab8kGfJ3D1LThop
GY+oqAGSWrF10FFW+nvwemsoy07ZlIe9uATv+H/Q/Ai31qaJxNIslQsSgg5Bz/vA
BieBQemc/Jf3bx2sSGj13ejXWD/i2le0KiPRcrJJAWYZZKtoIHWrBqjmpdel2Xes
YwMO5l13EDH8QFMkzKloz9oUdJj/Ieaek1Q4SWWytqF6c8qoF9QonvjE3SmASPdd
`protect end_protected