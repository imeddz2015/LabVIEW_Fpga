`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 28960 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/9huKRhRMtvnNqb3Z+UU7TahEoHV+T8U3P3ufru7l1O
3DlgtZzb9QxCbOjthp9+wDkjygH0eUfDrEl1ovhZG62ur8/hAbusuGiiehYDnExb
Snl2WiLGbLj3vE6+kkNqE5MDzEpjGccDYSYhWvMaQloZ/WzFVLFB6NzRynHdJ+Sx
nvr4ZxlJzxMx3YTPFwLBBwZxhfDBk2WpVZKYmXank9agQQVKyTf3T9+1y4zeyWuX
hOCCLzOTvP2Rpun0oDv+XAnYwQfmc+T8uhyzTUb4xozwvuVfv3TC+wZe0vcy7E/D
reeB44TS0cmsYsv7KeRqTPAL29zMsyYCz737hWlANN9HkXBCTujcOiZsecyOh6sG
Go0AdsYkD860dKw5IseONeMsjX2bnxUdeIQ+7Ifjl9iwlcQvzaxaNlBKdW4m92/N
LCypCkKKXs5HrFkCRFri9euXKJ3pfFA6/IPrlxeIM7SFIZtCAMmMP/6KYRKtgcwP
euzR6frH1NKgK4V0tVLBOrWactfmzVtUhV1y0yR+gcGzaXvNS2BH/lKNAhAjPtUH
nTo8dfQOaatg/UeWZ9umTZJpf3U41hgRZc1Dk+GPbiZu0W2guSvhQIonvZIS8lwa
omyEQY9wwekPOoqhJat8xbqTnJNn01HS5lEmGyhn7iTdvrVVi1ihs2katYB2Tt+f
9elAHe+gmY8JZI2Rx8YI3mWwMypiu+DSv1GJZnicjjdsu+KtgsgbmHffncKKHMOK
RWidYVSVpjbW6J2D6qqdpt/a8SmQUnqTXqO+GKLFBMd8rba4K9eOxcnygem7mimN
RMG0rsZvPQu0236t9EGs33PxTflAf3SHn9eZINU4fnO/68HmXl/GgqP0ic6eRYsJ
HEfkH160Iw1OX85XBJxnbS4ME05iRS6KrUh4IhVTKJBSKwnmjEYaTccVHKQgA6iy
jS0mB7DM+EYtayEttZoJDbj09l45fG0XbjGvRCruB5jICcJ1CqytFLQSAGHAF4Oq
t9sISQ0T9eIirONHFL5w0vzgw4kwv7Rq3y0cnFWoVxKzkz1o64M2jdI0SP6E13FW
cOQ6Uf/+ABjcnToEItiRD7xCERPrQJm6EQSbtEYkYpJAOSSkMioVnk1OzKxMMA9G
QhC5GeYva48D8RgcuV5N5ZbDUSqSfJd9F01cFmZwXSQC85P6pXLWO76h/EguGXTL
TvG2rjUxN/XUAsT3v4TxaUZH89wFgWWF9B4hcayzj6mTlCQjjPtoKaY9cx1vhLpP
/GTfXO2ASU18oDHul54R+tPnOqUwhugyEGw2A7+4w3dAqSTQHg17h2LMzxo/bp11
4kbYO2z2oiYjlj9gQqp7WwBDuYXEbk07AAId6V3KmccBLLgKoMjxnxylmOYV7hcn
072aqFehWG9cyDG1nGuyGVrrMsFqn89kANI28pzrKmxKX4SOzvhgfGgjQdYH9u9R
C79niiPI9Whe4q6F82083xWzk14PwAlSopcJYpSMq5ro3Z0uFWPJwWN+ijiGi/Pn
XLOMChfNR1HvgSAZmD+RsPuF+xKdmPhoIgZTTeuyOC6/LST3O5YOST9ye2asBBl1
927MTJHaENpT/hgzi5VfkGNWc7Hq0qIxQdnmM0DEqdLLnnuIw8A0dlll5G+6PgSu
EPaUbPEmVJG1TAhBXJFXOPBtyWWa7SnYO8Aln4lTjc9oO9W1OzjBPYOFRS17AbEN
5dwbRCyI/LsMKLk4AzmeL3DxYwJKjJubY7VcKuHc5LOVYbKGPrP23/OBQ7Naxb1y
AoYEMnLh3u3j7LiuTj9GN84SJElyJNUyfhyDDsaTdg5E7Z4bQm3OQUPj9iNuPuHM
mcX0qDqy9zYWMMARkeolYF3DGlkXfM9z65dyaAm5i8V/roPro7G3PbiYgUU3fuUF
GYF+2xK9doKBGWJWLmg1M7aSQgOLCdUGfxUOlkB+tte7tdUcJW19oGZO6y/dez7H
695hlOkkH56tc7Baa5q9zrfqMEB5e6pihjhsnK/6gjEEwYmY5A6tGf6t9U7OiIbd
0UrI3N9NGrKWUWuCVOEJZdVG0gqVVjIKvI8qPwlIN9i9xbLfE0BKgYw2WXryFnU7
vq+VYeQPDxdKsMKvREcxNbJ1nTBeNc2TYA/U+9ZzTrLewYFUzm8NVqFBR96ViCCL
AGwqwJ+k3+KDjyJN28oLaCQFYYiBw1zp+Md2wOFvurB88jeuqkHgEzDgav7f9JVC
oc9Yq1RiHFuX6D7Uy/7iUPHqFluOStcLCOd4BXIVaU0XZ6UaN1FEk5kMJBI/OqA7
4stUES8R/vZFTXoU7BooGXAo+2ThEh4A7pMPiDrd2JnOzYb5TtsTM8OReCLzt9hm
xKTYrEXp3H0aDwy1s+95M0eNdcx6CoSzFs1dut/xJdKP7QrEuAz8BT3VYDZeKw77
JFG4XJnv33crnrN6f2UGyoPD5MMOfOD2mfEoUH6zgueL6CidGvOI7W8xq2TgBzTO
OKUGCBGibE4sCt/uQnHDbLVfDiQ/d8AoRHKp/qb8ToqtUx+5vGK8HWW72BZQZXU3
aKcs8YdLCbrQeUhRx9riQyPxuVmS3lZ9YVc13NCdbQ/sdndJAN4IDpSyi1GTfh6f
8gPpqRE05l3Bk1UClYXkaP5l6Ayur0G+cEPyentPsUWqIlVjpUf7ridtu6tJ9rzx
4iEHkxBz9uvPbXeBYcISOiQJQiZ6X97qwVymthmX0UXm24JU3Hfq2r5Brs+cNJqj
pE8oRd9X4HKi2vyJj0t4dK4f1ppfyRr9rCAgEhGNQ8nZM4CMe8INxB/QzhLdnLjn
2ADU095QFeUxhjMjrPzCtx5tIqOGvEpJ53P6R+5loiOGX3GWpor9PRsklLx5WQV4
pf0yfP4WMWi3cfF3fiv4klwh7GUuGX7/X3+sCE+CXxo3x/jcE7+9OyYYduL8fADc
/xGgO/UVZCx18qkoxfjzsu/n2gxereEUHYNrdhL3AVQoNGqzWtPA2Wyej3hJkgP3
KFxfNnYxZtoS5rdPG1TJlAWTIT2m/qOsXTv1NOZoeS8JkpzFboNW/Fnjyzu6gKTY
QJr43GLChKF5E/CoBtDSTlzPGUNT28knxDOltC7UUiCYGs2Wi9NWpl9mSaIY/RZG
49DV2uh6umr/5usnooMRkgcN01vCw+QJ3gNqGbdumphO+rQZSrCHxnAsUCJEWxQf
Xea9cQ+hoH88lwDefShiJUCPt03YjXTJjhTDbgmX9mv/IlSKzdbzLJ/IpoDCbhnG
dcBXw1+hM4+O7q4EDioUwBqsCRW0KgqFffZM47OjFx5y6084KHjOtDxaMb/dM8+B
rv/scAYq4QUsT8zu9iNMnhUVehq1f/+OF7mJPJLVbjK/F2cW8s6a4hTWXniV9/wi
ovXDFb8pvk4DAURBW+IINzKE/hLBDkzx6uyQ85PRot20WDUdpSdDNjc+L30WJgQp
8q6q3+FRoLGWQonO5usNXaDiTPf3ObWIQmkUXqqAlCwQ02GpvWK5jG6C8n7mKKcT
q7olKzJSsr57z5WcXhb79eiUL8Amu/qef0yLeIcrnL/SVzWtkgLK0gV7xA2n4WyC
RxewCAnUCJtqzAYe/CTyxcrvJmyxuo7rtAMVA3f8o7x0o7VbJlfUkHJMs+1rrlpb
qaSqlDNi3EbVra6Df8ai0xijPpjP3q9SWRWLpqhtf/PLF64A04XyqFL/QlJ91Z28
kOW/wxfzioJT36mtYITh3YvopnmqHvbvwc1tMGXCKuGe3zXjl6sJsEDz4Wnjo3M7
8C/fM5jjXkcNH70+p0ZSQbscLepMC1bJDCjos8L4KgvW8y/dg1QYI0T/HIMZIO3L
73PHpdngFTBDUF5QwBorXB7Lv5wplZ9tfBkjNSppgohzbprbRMaEv58+0OZr0yWv
WX26/4jatYarwFaMUf5spTGL6rJMXOGoFWT++BksSTaDo+QZUGHsmFIkqUAtipxm
t8+9T7w5lNUWC9xAC/X7Ya1uWcuaTVi0AL+rxcrkUzr7qwwrP+wx8UiGu8NPLReh
9oNclOocTfbV5f9QJfIYHWRNw3tPRzoEfme+NXrTTXHHHJnsIK29EWZYZvd9wYYl
7YJFjy2X2Qmv7Ajet+nCccid8j/fD/M5rBbHj8deaf7LdBT0XI++I1dTU0MuZ7IR
0FBIv4aWvUbuL3Zg1JMTjAfKlF12dzxekoJVtLF+judCi/ZaLbH2fC4BtmKOGdLC
ee7Wm794huez4fv0E6HVQ5PuFBOOOnwoBL4mUaGDVt5iEDau4WgalTIXygJTDDAg
Nw9NSdZKN1fAKNg3qcPDwUfy4dKPQr/8z9QpwicPnV/XpVWEpL8mXB8IRHlot/eB
Aie2i4mirO+/M0UYAhXWLgW3i0eLl5kHevcjB1IiQO3+qYYWKJSKt/PWqpN1T3sS
pYS5tWXxMpeBhftJlG+VnIGbTn7kfa16+YBwOlR+AYPaGkKOd+pzEUr9C+plwlKm
Ge9JinDrAp34v9gvWYpqj13NNQOrDJ7n9+O6XzCUY69U7vp/fO+Hia6F5nAIKHbO
Hrg6qH2KaWyNSOEQWqzB/BL2t4BfTgDtS5W8bheoLIu3CDYP3Id84W/EFRbOs9lw
Pwwpjf0Ipmsu4V6fgTRh7kq9964GKS6Pw8KCJwlk0Webi+NdQerO08POXYB3ecvQ
bqM+fCg+k0yWE7SjVaKCr0GN6A04me7WiqpX/95NkfyLErOJJRB1WVq6rCEF76Gd
LTJOpMx0TdkeUqaRhfieTkfB4p40D8EJmtasadjibyFPqCZYUqdnr0J3GNz5F5R4
RWgwg3TeV0z7RTE+ajiPDETMTGUQVwlfOTnN7PuA5Y3KGGKrD1rP9HXZ3YHW8Mjc
sdPTp5xM8aivVieny1CFvFuRwHBC22q+oFH1tih3tv4U1W+Oqpn5y9kKr9IfTcDG
cwae9pUzxaa+ElwdRYIBKp5G8YAKm3FahKkiHdjRc0sQKhnxi4WWhxiWCL7M+nLS
3XuTTPy2ukbLYgomMYhPCtz6uTkrLL2pPqZKprGEwdwt99jBRF7EOBIDeXwnbEpQ
qIfhJ6LhD9itH1Y4PncWxnzRNv+/geP7T0+d4r39a+v+WosvNUIr47xOa1LlkVBy
GFkm/66g8Y4ebmds4wnEkAb6+mJIxsKaWPUcrY7bLX6fYEfp1bmqUMilpQ9t+Mu+
+r+yORcB/86HRFg47/MwbLLN8GhTLR6mpUGNewsR0MpDonGj6ZhbDXCrEXt/6ZKW
Kv887Trp9btpHES7Rypj5ZiE2hpG+/XAXn0ks9Hu9xbM/La0sVoyKGqgZ6D+iwSR
yukSetLmxRZkAgddMt7XyCRj8X81ovWLP5V7ZJ5tg+hN8uI7ZiGb4cGyBCuTjwm/
SE40VFhblocwspne84vNQ3B0GVpgGaJedor26i+f/yjp93Ldhmk0tS9Fqgy7Q74e
GV7yrdmAUtM3SPjBfW6SW1nMLceQQeDDEhGPymGx6DSeK2R7ZeIllI2lEJpd6Zr1
D0i2TNVsj/3eupNtY07y0CsOEgs5rr7yPC44E5bkD3EdyTCREWmxALamuPx1c9yu
yiiRIWISf4qY1Io+BON/KzzsaCqMckz/EphHmhI/MROQh8jnFiBXf6LqjhxRnQNT
+YqN6ggzN0v4O3i9gfY+WIrasABBvmN9AtZkPBQL5S3XTgxk5y1pqFFTcWmPBcZz
/YCk2/xA53npepkJF6BgoEElCPxuMrfMYC/Lc43N02R3tD9zq8pQ21SeQVEnFH8H
FIMZfbGI89ItVhryE/s/nWGr1AOu0yf9HucuRO/sBypldwonHl9wNptOOcEhRUMc
5Oiz2lCh4mLW7hbKQ1AQsOl14zF1nyfplX12pBenwvdIU5vfn88sSKQQXY0ONuKQ
aEren0Dwo9qIGIZO0XEshsZ5zCkdaN898rOtRunWmPcXZtAvpvhd6maMtdWVcHmC
9YNVyrJApYl7z9zfNLbLk5J3NfHFlDIeN2SggH2QLtIuviMSFrNObaepa7awNt79
rEfAdt5EzywpBx2deTcPwLx6OD2zuus/SCJi81NHd+s1UbQ+DpA3sGS+xHhp0UL9
hDbX/ZKXWg15BlajsrnQ6e4jWysTRnMhQ5Nc7u4jmZfYK98IBXrwdo+2BriB11Xm
2eCYP2H9x0i49q4Z5clPPLCFFAdRyX3Dl6Jz03JsqOBS5xb0ZOLyCp8hQLccXRZc
/x/NPPlUCRMp1Qj1fuYISH1EjtYeYEUVGlkPN7fa+VCOiavxsglXR/RBhlaAgXpM
BW0MAYPOdapXVc/fNAf7mP+9NiWzl0P61cOueeyPfdT6Vlim1YVqKwXLHpFGT7PP
04pPRx4cneT/lnK798JGM4qCX6erCYtAoZkCTFMsneqCN03rL7bhUjQFa+ct+jMn
hBvElvS9oXVfpd9LmjdqFt5xVKp3YoD4dHBwMCfekedVMb6J0oSIpnBsX1s12Iz2
P1uomUSBr674vzujaUqC5NwGHubHROol3E7xkN8ZYy5hFXK9wto1zfMOApP7XIVN
AlzhAKxSFFxHA5vB5jNWvqlzaLGBVG74FVXlSovHHHbIAU2A7ejBBUJTNFkoyR0T
mlKlKVDaDc1J8tFSMgY8FyiF1PVGsxtCknyWMg4lj/RCuPnDhIPyPZAZh/2wbXG3
aqII1zGvMSky0rS9HBJpjISPzaerByFydtt5epHuAj+enwa9INbCTiuh0/SUzhKt
18ApoXMl7FVaQoxfwOaHjxyJCXGBa2gH6Kmz+YIlAL4EGuV85g0wGL4b/ow6NvU0
+kTI7o0qQjExEJ/uLomuA8QheQpe9I4vIsujhrlWNHJDCI1MnkVrqn6LbNpQnk9O
6SMEWrgn3/mN3okwyJssfBDHY+5WklQiwsZ+nV4FXMWIlMd+zBiYwn4DIBYvbuYt
F5et4mzbql/zWqkhqLma2D27aR63e1ZBuOudbRmpZ2hCoCgSiuoy7JEQUUtfsoWd
Rp/XeOR9kxZOQqeL+Wd8K5YcAHZTXcLi31hHFrF9sNUh/ByImtPUeWrkkdCaWG96
mcl3L/DudYtMQqLerGNkRsUp49ZpeUVUmQhHQ9Ud5Nb5vcfW1HdDVphjSX5ljNR9
9J3L8xI/nTEYEHuP7kUr+fscr9fLRXsshu2/tp/dvVrjScf17gB2PsDxB6hqpDYi
RX3XafkTT/dKRVN71w1yPtf5a0JdKyAB3fTJdwcu2H4J7/rmYzMmvS8nCYx6IgT2
2J2LXeFvRG8RvBxRMHpteyEY/tPFvTk8gXpj4IujeQJRuC7lIb/w9G68Vczdnb4L
mIm5KnAWaNEvkqOkXSpcgwL5BTVdtlXW90/dYTvQ8u11kEgIc72DDZ3vaIMtZJr/
UozdggFUOO5buCiv2Ne4JKgMoGzzzsdtuvTtEXAuBPy+ZVxTVeUe7tQWRnz0egDP
UyqNvOFglvfRHhPo0opaHfeRQIQb9dFHpPSCnX4CWJW6F4JIGv7VPLPsKxV2u+j6
XkRKlrCRk2QPK1S8SHnXXn/YlRaon3vhrQRk2EMgo+/V/tWa4qi6iuTG7VSwKWG+
s5SrqwY37JJmmx+YHxOVm4iPdfXiUx+4/pf13vWTf8O4tVALMvI3v+xldTq6ipRC
pPgSet84voNTQBgMHqSFo9cEcM+KvXBxL46URa94S4W5mP/CUNM2Nyhi9DG4Cz79
eLCAliHcOms65iMi5dWkqUE0cKLnLuJ1n9GBpNcWiyAGFhLBM+5fxL7qmj02ZwwZ
VbVhnL8RhR+Ag9z7HbOFQD5XJKx6a/9bw9le2ESZZhcRW8qeuQ+03EcCZsR2P2Wi
530XpucLN9kcBQayjXIhtJhEOgV07Kw0XxotKiQuBtgM8YNlGGzUSMKjV2711m71
SdQ9PahXnTkH2Qt8MIhfZu6bg5Mxb+FmTKneTNL73udNhpV/ejJjx9yvf8UbqyPk
I+gKxVplNrCpOL359u//H+CtML9hGHcv+n9SkaHDgrVNaSWzLJhGF3z3nHwD+hh+
mGyB9gJyItSbk+/xew7KIZyGQU/fAK3ZHUsK3AHxMEj1mMFp3Xh6hkNnKbbOUvy+
f4MufKVvEQCI7ZFboXa79h4BfAp4E8cbryqoRx10ZLUJaP2sMq7GjyvleM+Qw4km
VNvi9hbIlJInBbRSEtYzHDsVkXhjptD+wO+rz3jydlatZbIJtnG3lsYdx7nL8jPY
HyOO99E5Jukb2Dvx0yQLmXpNRyimj+npg4iStbaulmMVx8P+bcw29EF//ZGiKQQt
/ERkQz3XFQ4tV3nPO1RPZQHk4Cinb4gNLEoAXm5jRFiJL11anA2fiMj7OYnSN35Q
lE58759/cMPA3qJsz7vyQZi9BPy7BESRLH/ADbA3VjrCTxHywf1s5PqTKlZnStja
84sS+bvhwhi2RA223nPhtuYuGx/VxnvxNOuTurWMCCZTWSxdfEgJwE5A2a7KNRCv
qcAfgvwGmahnv6VzRQWqyxdP3aKMwZrtoP/RIhQJckmad7bzAB3SK5/KV8Osoykt
7+cskvUF8++Ul2GMw4PWgR/Pmhrvo0nnD0Myv2ktDceQCU1nBJWs4nhHx0roncnT
OBEO6N/68l3oejUL79Q6vqrr9duskaSSVeKfrPS47qpS2mNr9uhIUok7Sk+jVrCF
PwRvijGgie9QeEe09F0rFBdIAElkVMxPBXxYh3X9EZZkGWIK+vMHQDJltt5Wda3f
8x+heXcKEuJGyWqbfpjztLA/xg3FHzMRnGVT4UR3+o3Ydj50ms9S9oCif+mJ6CQ+
WZRWFzXhty9csS+uRhhHaZIbjxbQI6IBsXM7nmC3UTG6OcLAi0ZPsUfCJ6926I6y
eQ/1/roB/kOOZ19VAAeOclwWqHx9D3ZEvCDBfShX7yvIqYVACWZxJ9TpjQv1bLwf
lZRQxeQG3rJpoqVDbvzyaMnDyAwq4CqPsGS7DGEYKF9eMuUmlgHHVbBzv9MSuY0O
vCnZm5D7WUejl8sGS/NYJI9ywbhCzjaVNZL3vtMhLMRxG8RoBX+rlkmbt4zkk/YG
Uw/xcnbfUFac8An5oInjozYNycBkfJ6Jeb/f4WaCOP1Vq+3I6tfcVE+e9ysw09Gx
B7hpKimQfsudGUklxZB8yqt9E81hIoMggjgMvhul1pl0Tf7NZ2tsPHzcOUdK0rHW
JDMISD9nwTZT8LMdpQVNNn5lspRSosmNe7vBCSysYEt/RIcdiBMkIJS2yZImnC0Q
BB5vS3hAkIAKQMG+gsnPbiAsNb3BajHhYQ54g9EZqM7iDBfyt15AzBkEFlOjt+Q3
uZIXZpl3aESVc9rfCAzZ4aofAZm3ehO0C27Qn1uW+87oafmp08eGD35H6KGXSHRA
Gsu5gXRUuQgW7WxE5G8R69WM/993sf4pBVKPf3oiZyWDBR9UoZi26yTyGG4u7gfM
Tk//C8q90Ps4CaBPNUR0AqiEuppykOvD5IyGfw0YtIGBjV4IemJN8+6ZrM8d6uD7
o5FDPWkcSJiuDiv5DXjU7sILsUG1CRb7bRp9FcD4BOelLi+7tXcJHDJjyCZVg3Lz
4bLeqX3lO0ahKWpCKmeENErO5mvLJRffKZSWjYNDEIbtB6H83YMHNJdaxGR93iya
qSGDDIBJKz4rNxvCD4YaRk4Oceeq4M7fycBlOu/NVXyrVm21PMfMB1QzhbB5azMr
n4JleJbUWvnvkLfd9I/lH4YlrzBc3GMUVi8x64X2OymsTXYWZ98PUNTBqIxNCzY1
IHSB63wZlLi48YKye8SUu2x5H+V8uigpo2A4qsglGlz3EhHrZ+PKuOXjEX5aSuLO
jIJPvRgL+YmvzY8kIJkSUqMjMw+PdQzylfUH2+9XPQqlwjcNkb4rubMFBkde5skV
gDGBXUTK1goxQuZEr7YMb6leuPm1Q/JAA86lRml9PWVEUrNWXHtZlwP1x11sSPW1
wOD8SCoDYEMetE2AEmOCtLUZanEvu5+YzxnmLp/SxEvyP3d09vnRal9QSEKu2NVK
yUDtCHsBijG7B7iC0yrdtYqUlUsOZ8lcj9H+vMmhk9di6MqA3cbirA+kiD93APJh
4Xo+9T+OBHVdcEg+iVvgGHcHlfkkome0oI7WFnXiEpiGAGDKYrkhxLhzx4OOGvJp
ECMeLuW0UKACXC0ipf5i8zDY7duAZXnWo32NUxyiU1H9b17I/9hqbxRhUQanNZVN
3WbNFAavf0AE2ALP8GqB9UoFUQ55FMLzVL6ex7/2Lb8wvHnxMQxdKA6MSduqH66z
4Ck+AH8qFKQwIoRZ+k6ogGPbt+7mCao4ZfAqC+D+1CSpMS3y+wrlYl8TXNtRa7eP
pYzNl/i3Am6EAXy2ax6NsReM4QgHkj+2F1ac7kUNT2MrB6pqm30DpPDLlyBb/pME
lw7+UQ8lcRuXIQtzXjZU3HGO5XFWVnBXSIK7D8cfSD7wpd1vxAp3PgbZQ0+AuPZj
PoeJ635ZoLR8loAZn8PZRsB4aAGsNSzbEDjKeiyVVw0iHxVytvl8jCuqugg4D/fb
vO2QN7L9ZTrMc/fvaq9T6Fyzw6+vNnI18C5nGvrHZWVAbh/RdAzWX2Bwxmx32kV8
5uggR8fRE8AM4pWnM+x5ipBkNjjl0rcU5cZ3loW1gijAQKtCh/1wMiGG8h8ZhQ/v
1/QoFjq41LQVXk5ihDvU4oIVh8886xgsB6gn2jt+pweyAaaQIT2+w5XPojz2B5Z5
yubl1uTG20QnMvtiAnIB6ruGr6smP/Dr3E8ifNCQhh/cZo5CYfqCGB6YP8XKZNXL
YTTZTRF24LF6KRgtngTHgo6Y8jBj5yUlR26mK0pSd4oVpcuiyXQ6wn+mORN0eLr7
z3FIUME9hE8dRs66/5yHExOKHZkvYxYslPxFq2c4xTRrpA3TnwoQpk3Pvh8NOfB9
ZAhElkC/e0bbh7iSHTNy8BorK7ouBKKQHkBTurQE79NilZKGyvek8sjkPtwQW8eH
IntWXxDWqk06Uc8x1/tZ+twm9iPMLnZX+ASlc7TdiavkTmTNft64vw7PrhrEuYgY
HpjQwaEo+U856ssB3YeJBAkaMlb5xQGaKHT5wz1b9ILll5/YXoew9lDxfoDkVBqD
fsHxdev1izu4UFKB3+cBwni0G3GGMpWPNCqteNL/MK0ZEM5FTfArIWCiRaAYbzd5
iuQUnWvXKrNQ7/dUCfqJU9Vf0En/QbP5HfIxyTPjWpaZnsWHffi3TckYPMuFJLmo
/o0lIgTh7hslEDEdptp1CVfo0aK8r7DnemzP87AfRSPE6muzy5kFG9ntt4aDZo6Q
HKbHGCUNoCSU68xGlWDaqylK4Cm+Rr+sz4Rj5rIX4g6kj4IZ7mTepdaidYzZHwOJ
AVTfGdBG0JC/LltYHVq+qS98HC9hZB/oulOsbU0BYKyinVrRYMzlGc59OAuEASTj
YqXqPCwLh23Y7U/JvlWEsTUYhA94V46a/Eq+WclimP+QTo0Xh3HL0jMeZ+9R30j1
+ILpCUYcXdUoC1aIyhkMLOXJO+PrmulpwqH5vdmhYWzPkWDMGAdL6IfH4U5rIYQj
VdlvTStDIjShhAbFNYIawDfMyT84EliOQcMMC3g4Ws+hfqkm1yA7NoRPymAGV6nY
++WhNZun65xghlKkaO60gIbEUvEdKJ0Y38082gu2mCNE6ITu0UI1iKrKZRpPamin
fdsEpCGLMd6hQow3DmETvY4OQmJU0w09WGTr7q09Wpq58Xx81JpmpNp6I5kHnenq
M6cCVsqA5kWlBonRwzO66wTpgn9tQKolvva+TlePLOYCErVwHuJJ7Cj1zWQm4E1h
udicoEJ7iafbY7Od91NHzx/JAYrWU4/WfDa217IywquzylqcltAOEKwVM6U2uSMp
5ammJOaqGrIerC1sMVvEUzGaScwojFWpqcJSNnHwOdEmBREN529D9Jkq7vho1lMe
38i3S0Tlpw0xV3dCQbw8Cjw/DerSoZpxkBqxObR4hXk/X5qxejhUT/CsFpJ6PcRF
G185FzXMVLoVP3G+55Ddiyy7I1jyrdgomz/CLJq5j0yA3IYxXcc9nXK1mDzYfg1p
fDgmDyIgnj28ouKNU2n41/+Z2YrnnBXeoTvqqj0LHpBlq0FqCxQuViFMajEUrG7E
Vyp5ozJJ35cxVTt1byo/ItfgsAhvm6New47u3GSPsRgpZ0NtXDs5cw0TKExPhJGr
8C7TBO0C3Ra2w7mFspXIrzKBLuqnY61l+1qGsrG1Hc69H0vAVKBzjUTxwmiXJrgG
2oMiY/BKPU+61mTb8wMimYPNDoXVNW0mfhtXzLVU5alDhc1v/sIk66PtXerdDuCP
B+7p2zuQeG4A3+EUEgZf6gz9QB4yj3SQqxg0f2nm/wIOS/mfy08zOquC7PaoxwOj
tVcovO4NSaSK3yBtAlLAiOxnu76dsr28bn1P1lcqsopA/Jnpig7ieIHEftIVJ53I
Gwozli++/KCRz9qBiesXpZdUqKJFwY6NsnRydUubRXB6JMo1G9I8rl6Hy522Zj0c
STv1Sqe8IrPXiXXE33EFNpouQx3Q4LIzOtdDgRVb0s5RQh7GzVxqsU1mwgr98M4g
1XMAkJU9bCxpe/rjAHdwus0zptEDpAsNiAGYxkpp6CaaSVqWkAeiRTfqot5LIMcG
3J0VyiKcNz7jqHaVpbkKsrWKUhUQQ7hhm+AIkXHjzw/IQRANYUe76zpYTo7DGMqF
5WrkUNzFqTS1v2Od4q4KGLQQzjl8dawAMra325fFS/5J8FGxX1M/zRgDtgR3X1Xx
191tZVCSJeVe6ddihqB8bBzmbVNGUHcOAMRp6GW2j8GNpOLbbfTBe5QupliHU9Ok
mKq8+DO9m8d+lKiYSEzXb15ORqo38hLstsCTBfVZcYvoWDPPGXu/w9j6apa+kJgi
xcDLNWqPTjUzdFDlQBZO78OJrSz6ls4f1pjVI+dLwYlv6kRMeVv2SOH6d74dwqWD
9w6BI5VJAp8ZtAwgLDmy/ATL9KoJNPM6ueHFwEAO1KiDQzKhlPh1OQSW6cBnzuzF
bvdq7ZIJc4/Eh+mYkZ77RxdrrbSL672VWBdO/j+sNng6HOeZmkQzHo2NcUKhiohF
+xh4AI5gKpEZe2ng2SYKrSqUzHSASIdBoahWFA8/1JRKvVc0Sb4J4hfoylJ39T57
0OAYfCbrPpkon+uuw94ZAzRQsKUOH7WEV5h+J973JpwdwfC4fJ894UgOeB5m5wwI
eZlElBIBO3WZNlpuEd8auw+nxbn+OHFu7Leq3mGh4rQo3WgcJrt/GVBXnnQzkE9e
KXEQcdOCdoLFkLTvzNwrgkHrEec2p1oYKy5Bj9ZSgz9fWKOYg+1oyqleiBoSgVVE
fZkmOfJKFfNNltDbpNANrtDzlvwCaXTSJ4G/9ltxbYvsMgOSCzcBevFYW6N6i7LH
UhyVxYpa8LZS43JeQ7pK7lYv8+UWos7cYuJIX5wl7F0dMoQc8CRhoi/Y/bBtCFyg
C3vkoUU9808PrwLbsvvA7WrTxWH06Lc3/oGZpFsUjE3cr4uAIzDVjzZZlboQDdwv
0Owq1E0p6uyABm/wGknduD8aK0qbuJ8UgbL9Q+ES4sGgzN14I9VNNCkufPQ11BtT
gjoKXuwF/JHezhjlBrzB55c0GYvI4tqD/vu6lrqTzn27ARQhJgNGDS/vxm/JO53E
iS7UlrxrOalVdVW6C1N5mKG1Q/07OocBU3Sm4hLa3ObXapEwPxqI2T3wBD3OAyDd
KO6eupWr+jgJYwnw5+UWP8DiLdDwjRqFD6R9bXQDYNL+GpnVG1Raw0EMya/9Wltf
MQZ/mvUubZklj54coyqB6NJDXHZOMvoeHPK94pUkpMLDZGf2ETlSTY35uIHUd/Up
fNxxvmtCEadfcW3U4rsaMY6ZGa9nG19JyQbivETlQqKRlmu2fNeucPe3nGFzPEBl
Pe5Qj/R/lQrTXvMspmB+VMpr7H0g/nwg9EMlJljUDY7+Ehk4PMwc8Vltubkee4OC
HHb6GwtJHNRAcQ4xYTt0jZDzc4Ly+NtrN4iKP1aGaWQP8WDpS23mrV54dlt6qfDL
7xvswHZSNpptyiS1yhFEEktEbpGJg77jV5bQv+GHpxL4lBB2dqU7O5T4HvCfkNkx
HTimdzrXmbCvy9sh6BosjDm1VOA/TvIRNxd6xv0j4uX6rkSOU3S6PM66jdp5WWto
cOc85Wu/A8YvcW8vSUId929jI+wSFCfrJ77PnxoUxhji7BVgeNc9UCV/74EnhlM5
fLdCteyG1sGJMbvpT4P82SHfPWk90LUAgO9Tw3V+f69elXIl9MKuZhfLfRLiCT3b
jPAj4a/SuMnhzFbHtuLt3HBsUv4vCHB/SOswfPaQo71wRhZX4o+26xFsGeSCnulf
Xmp+PgAeupXM+na/l8xmqmBJNC/2HyDSp5TEzVZziHeGeUAN0gNtWzqpIkeDljCH
+U6d8qc8AXHJAGu2WOc+q5jhEp4fVTdyp6YRFuAWHLhQC2faGEWz6W7ET/u8xinx
NX7nRN2U6EeG2rn0uVde3UwBEyruRjKAww4k/xayOzLQMmTqUyqaWGlYtSc7NDEH
iLsR+kd0ngCHukpXstFpOFoJ43BaSQA2cXauqBRwNHS3CSwRnmnl73eMBXz2c3RF
EGvPC46Oz2YaCZRoH44SWpWAGD5LhU0SyNQOAkZT6gJkd6jA59q5V9Bg/21KpZoX
8AWhIpy4NnmZaG8McMISx7y1DFyAvJ0kqYdV08qSAK8933UV/hbFsDojuRTG5O85
ZLBsOO6cPU2HOsy/AppRua/NCmixjrff2w209hqBEpKQMKCoay84zqnTT1g/8Dio
fbCB+nHfvQBGSNsLjm2vdCK7uSQyAxTZmrS9ieX0Gbu2WUuLlvpC0WQZBbBEVNuB
n27nFnBNyTHeks6CN3awfmicCLC7/MUOyipbPYWZquAapVcx8BECM4xg3bGWdWZK
ULm7BfhxiCx7DqVj9lCTloXt0eHSSAA+GSYXoRifDrRa/3FzOoSYaZVmwKtyncIo
fF5+oZIuv0rMNPpVbRM4kOxWoCVUPCnEJBGQbq/1wGrWsMwSokzQZiKqbniRi4OB
EmoCl3ombjOtolQI0ierD3BWx7YtKskeuGrFvBFfElfnrL6ncxDPafI3TkPkNXgI
ZXz2uSO7oyVH2XFpABZyXyuhpjK0V3sJDJkvCEAeFkonB4ODwb9aHN2VNrj1FDDe
UvQMJE1pG1DWQmL1hX9S+01mmmdkT+ObdeAGlwQ6M5WAGtabGXJaSNIiHCTFhCb1
uUwf345aEwYq+cb/8THkwnhtVOX123hKe09M2aBR8KG7W0ps5TE47hly+wovmJZb
wrnlEAN105V+HPHNvfUNX8oVkLngZWKpuggakAnOBJ72x4mHzkxQ950HPiKcmDW4
UVtqD1Gx+SkNMfFbUm0n8G5jZk8pqxB/ONuDcDCz1m9kcZ0Hd1sjI5whM0oe15do
EAqYqEJ4UVTFkm+ZKF2HcRdz2zk/jAZT+kZMh4tsCPlSPLIzXlLPBfyBqiFbbL5W
PNARzfNM09WIF/gEd03t1KwdWmv7xGBOM0Kf139OqFKQl3PT0zH2wsl1Cwwh+sri
awK8uNRyLd/LojkqXqdVMg9Of+Ds9Z5xIXvRg76Xq4RFLFPx36NuQ1cCRvGiPIAH
lGXlMWw4tEuCnPXYJI2GhD1ENFwv+jVKozzIH9zTQ0rBYDvPfGM3FjHERwQCdCwA
S2sAVTbw7KL5ongIeZZAjRwXuPAr+uPl+vRCe2fwTS+yBotTPTSocThqv2mxGKuz
ad4NlUBPiP3dYc9prwT13prRh446qcMtCSVGzZpzmb681GcDob/Va0ZNMJE91dFj
5R0flolCLMIf0e8Vms0Urel2pUHA/ZY2OP9huq34kFUyBRUh/m4a+QVvt9x9hSIV
i2uGPoE/+rs7sKSAx4zLIcVBxP6v1OOMKR4zqv93ML4/Q/ApSVPSVLEkubrUneFR
rgt+z/2E5b7KbMRQlfRfXewKiIKCUk95ftC2gNKwVcM5El82Cd/IUo3dQqKrUD86
pZu3x/8ao996jl0foYk34jNYhksoxOiIm8QYeLnuCm1SJ1q6qTdpWBoiEhLBCKNT
dHNDXcRBFv2ammGp/9miGTzQjHKCfH/i85sLZ1mJtjUmi3sxMA4+Va0A2MOtrUSQ
E8/XGg7J/yTtqKwIqPtX88GfunPp8c1fMPDxh4kH7MKLK4uLwn8LSgbpHgIxk9gt
RqLNM/T9xBkpv1RnGRM9UyoDchXcB7rCTpt/qvHO4LWH8VvDk8CY872ZW1hdZa7R
p5T0fWInV2zzvj4wT0ft6xePvCWSjmS0AaiF4sEgSHxs3qW7e92tJ0XQke96stz0
KvjR3W3bJIhGs9hFTNZ8Llec/tUkVswQ4i8IeOmtvqa508xvWrusmZVTjYAqKb24
HmQrWNltfXwLTXNzNgHZgl9JN1T/AEY9jmJrTyFMM3lJPyyXVyeVNp1Ya5bFNs3j
0C0WHJtRMrJNhgfEZ+qO+FMri7oc9RH1gUIgT/6f1LzwAP9mNp3gTercspB/XoV/
osKvLM8R9XlMVgPkVw3zO5qRwdnKUytdMY2KKYt6817Odlr/o2oJvbGwefR0gaGh
k5r1fVxIW2vdiL2QqutzQKzpNulcATQmzwQ84bWRsTxWCddYVT7REjNk7T0SgD7a
GdQVDGycqPtIZnjW6WeGCe9Z1VjzcQoYspwgY0h1WRKEJ9bQJJY/XuDytmzXLDne
WaUVsl/C7FpbuF0sdBLFpBzMv+4nyfW4UcelSkZCkHBlUQH9lOLhhvKhm/y+4ZkW
inuJbLFI+g6xJbh5dHX1mz/9RNJpXYn/xTTE6Vx2k+b3l1arB4sE07SY61+8P3vB
HEgrWdXjI/SOa6I2zWi7OP3okc98rKgPehZSS85+SziBtR0mwTaZPeT3UYSdmWL8
t3f7Y/Kei7bSfiWO0ToWFnEZzDOQHg5VuJBYFCJ+pQFPupIqVMxSns02fr7RYqk0
UBqj6My24dMo93ERJi7f2S5cX8IJ3t1P9ME6BAg82ilN4YEhSbhYJ/uUnLDd5tvO
eyqwCzb9CZo4FvBTWr0Eo2JdnfoXVSd4sRIvQ+3C0hisEXscBmGitqe7bgvdnaQc
w4ujieX7BRDgk154m+gkbshzm3m9Q9PRut79DVWuKeD/Ed3zFEuQDJkGTUjMPd5Z
pnFZJuaWkj7hr5urt60Te7ju0Tx5CIrg6jkuVy8Bm1GKg3fNptXaobBWAAnzU/Wu
8/NFQwX920zxTC+vSz3D8+BlqtHu/OgP1w3bi0XBVhUGiAKTF1DCW0Gtaag2mB1Q
Ms0WDGbZ2DsmEgDAG+HBioESKxdE3rfY6GWwpbjudOTcwmWYG6X5OgQsTkfkowHx
dQBfWWCnNTv0W82352zEYpvTTSWCIIwhinqOBJnqDFsYlMKfPNSxTQwcUjzLEpSS
0n3J2Jtbs/MMJwLi9QPOJ9Cq9b9MgR4ozXapB97xw7nNNHSxbn+ujlcWSycoeBUF
tYFEVDnJQYQB5SKXVYMeek2o9O0xxRxwYNrhtP+foqq/GiL1xlCF79efXNzSNUrM
HylxWMWy1DZhXe5I7iJGjEBI42r6rGr6YFnL/RniykrV34GSh2zVlgovhv7t2JkA
d0UazBq7jpa6bSEcVBkHDABqNtuq4NPYKhsXNeuNNlweLpjytMi4Hy5qDZEPfmp5
0ep4fd5If8lC91QiAIvt+I85jecoxptwFm7a0okMRwXrDpBYcNc++ZDpbaAwyYaH
GT3HTwqLX7Cyp03iugwbuzZXBk9xR5BI2s9kt78yry6xhBLGBdnFJ/ScPVfA96s0
Jk3C7Go2m3IGIIXjxapfu7YPiCKh6BfB4LhepeqVSURzWo0p5xyviQNc8Kbqb+/g
oHDG+x+NoGcKM9rOUp/K9Hjyuj17zlkFOt0Y+o3JL7zKcSa05M7BcxNy40mWcztU
bZV7OzDBf4RqWpj/RPYVCWPLpgusXqi/aQIZ/wa9HFFyCIMkf2KYyNHZ9/Cq+EMj
OmKzYZETBuhb4k+wHJ4HE54/dttzc/TzOFuC4Rxqi4Wb0zb7xokU90hMEkATxYmq
/SlWDEnb27yM+0eLu7rNmA24SWJvAO7Hf3ek0CXszwSoHOoqqXg9e/MkaQ+KgREK
U+xu1HIimuqgCk4ley/yYDT6/58/3Gd+5kZHnIbVs7sVGnfCrrMLQ7IxYZucZm/3
6X1Eyh0Kbna0do9pvJM4Qd5WrB6FAQaGRw23TwbA2I6SIycxhXvvSyID9I0EjfjY
scQzqyRgqD/LrYOkKOYTIU8mqcuugCmzOf+2HIg4E2QwYrSY9U+0cWu730CY2RMy
jvuKGljzxqcyz+Ov7iLmfTcETEAucszPLZBqkSXVLu5MZso8awpmFu3ovASpjThe
0Irs6ammvLbmfnbUd5cq4qOSX6AzN1bZFaZ82kVPEjkVIkjb7LxKAif2nENbRJmi
DJASdtEzuryyv2cFIPxf1Ztgk44spmW7+GkPVlLy9P0U4+4gKOIEPxvtlcD3QCG+
/9H4/pUUpNk1j7rhdS/NFzv4VdsVIMNSPzuiXMLfE9Gs+R0+8xyQaqzgTgP0ilLP
FH6A6zCogzc6SS4Po21MKo2iLam1wH/KQ1iUvLVfI5GYayi4VIuBkS8sW6tU/kOb
TOeCb6/t8hqJU13TVQXpKXPiydxkkQWs1z9CvEwAGcieAKKtZAIkngun8StyVG4C
8HJ4gadc5w1X+k1ePRWu9pXckx0KSKZbmbIT8x1TsSKNQvu7LcEyvFLYO45XIP7Q
qa8G5x6PMRn1uFZ5IpkpBKBuw3SPmOrQLjhGMt34Dca/sJeayzCeaF6Jxdu51t6S
reyr7PJEPIkih8K3yS7ds4T+oZiC1WqmbVeLvhxRiQYHRSSnhXKBSEBnbLdPFpF5
k6r7Up6xt6/yfaASDGa8gpHD8cvvllNOq+ws5nbE1ucE29/3VM6Dn3FtuORMkbLb
JQpMNUDjOHV2HImxJvcBb6ooxhpjHQb/5x/2UPElB+KTDznLzCa+duGXxjl8cwfp
zSStW3b/3vEhhxaQTj5/XalmFTADn/VVk4fPwdHh+t880pFinz0pjq1gV2w02txE
KoZ3cmH2EOEDhNbRPBfVaDItYqIUdYbTfGuO2B0TmHR/oP7xiGnLHI5PHZcMCOQL
CTemE+vRIbP2ngrFF6Qw2wzEuF92OZ5GbgTkOXf+ERr453hFYx6xmt1iGXMcnVDC
eo91rM2CMjVkq2Paz+2eIhveex3KNpYUi/vQzswqV3noKTNGQndS6L8fEXmnAnib
EL6sT08ECjBUIk3a69Re5xJXC3HDGdSpDSMKCXFO2vr2c95YIIYderu/E7fC2Udl
RRM1JhHivMKQLY1YMhF7xhX4JGhmJGpHSiRvPYgaqiMKrYCDTcla4xzN6sDRTt9g
jKOs8/Hto6C2G23WDUyVRk5etsxqFKgBRkMmxzFqs4SB78Ns25nQ6Qvteh0qHYbX
cb/0/lSjP+glpFcZK26HYXu6XeCo5EQdTq7dwKq+QP3IUjW1l9WJFwmSB1bV4Eda
VZlFaDuAZ7fjv3iO36+OmGOoTnRsOtrtikdWtWDzeemmQ6deD45oliAIJ8oUszAS
AMCa6/FrAq0VI/VuASemyRiTNELjhq0yyxSp4JvKq0UzUWe1P4KiXflRPvC7SrGo
ybpBxSH/QsUYZSDdQAx1FK2Vdor03WXRHyh11R8txwBdNm4yjC37pqbxpuzTCMCb
bPfQgqg4uKYWO0r6qGfX2KX+Diqpxv9nBwFnxI2qq5gHd7pf5EiscFbgMhVDeKpU
vjPqi3ukYGqx20qBfMrOvyC1hBsNY0zPRswP0/b0t000iXyxyBd3RHYtTJ/P5yMp
tIq/9nSEOmfnj90J4yUJ6KKp0KuFaTTVN1i0iSXOXUqkabdCj15iLX3YrF9DX9Xt
DtQ6QhrDD28ylgiH7G3gogVIeIUPuBEHUcJEPeQVGIFMSZO6dl4MHmm2OFYhHJhG
xYcELco7aTT7ga3AQ5l5aCm1ySpRIwe3EFHriti53S3u3jJXQXvII/CN+Gus3/ek
qR5WbZAXU+jqmpApY18hPfM8mRkvwLwLU1btyQkXVKUq1BDxE34FY9p3+j/WEcpk
Ak3wrJzOISlOwluGgVjajDZm8c9ek+8n2IPHAGAcHHkkUMIVw8ihXE8sGdTnI1MZ
x1RYiOK7q26vAWqNOhO7SHmSmkVbFexzOMyKBEfencFPcMDtBdnhKDCuYZvr68Uv
B0cKSStx34UkNd0EB3yK3lKHym+bTP2/ByGAMWqEK2eepmSy0WjGu4tIE4fpW1XC
2tujoEmBTTC5/+LouFsNkRoxUAH+t03OV62Azk+AVo3q9H6QjtoxI1RW4GfRp8uv
Y9tdQbPsfIRQ9OzYnGs3wFmtayy+DdDAGALqkwasXbQ8XL7xHlvG2DbZ1uRXMmw0
SrsGg+uwsXlBgVZSV8eILDzWckvIriI+VVDA4BTNiJ8NRTXVmzNEBOAorwnyRHHA
8tPvGBeyx6hnDzs6o5Ed/FlcnytO8ixHFv2iYUFvq03lZPu8GXqdW5aV9N/mnij3
Gl4q9EDm+E6hJsXsZvTDTfPZwShJBi6JGZIbBUibuWlVZQ5HwVOqMCoaFRdXU5ic
6fnsl31TdKs+xUqgGaLasavfRvPMBNnnnGZE8OBalF5ir2b5HDb3q+jCWx5o0chB
9Z3HzmxotEkZ2KkjlmJOqOgHweCMgd9wocmXLIlmr1uswGGN9+YP92IGL/52qee8
1I1eD7tfhDn0tENJQBMEiKPkvMfA1LQm18d1UvJzMXsL8SSevPu+8tMtJ41v3sRJ
o7ZyLm9HALAGwlKP5LYECs+RaEVz6oTvnEGsw2+EMiWlsaFMdHOjEx9OU5Rq84/r
Y8/HdtZ1kYPcfucxCnNf07RYP8Q5PZuqK10PNd5AO9i7maZfxT0V+CoV4Xo6nBFj
U7r/WDuKRYMpDQ1bq36kW2lYJLvM3PszW/YPPrws65CAD5gV0KKGK+j82W0FkMZP
YlTTKSJSfF9Vd7f3Og0TcD3MnEBZylHTK2G1Fpn7q3cCkf8nY2MgWDCR7d8/dk4v
fZpHfeZrf+4eQH2MgVWEmhpzthxW5hYXlVboJLONwEHeYM2DbTDaVODtdiVZS4pK
mHzkcydQN72rum0l3A1xfbsLtnQ1CaXM6p64yr04F0s/Z61NRm+NqMRFhRHwVXaK
0wTNtN9ad74UgZfdgTzWq8sqgxK+ieB+/Ixxo+Wka91ZqnOGB03P3AmVJUPlcE32
01RCKX+0awC6lL13Z4TYjNLh/SrRHlUftZO8jnx9OtmGek3x7Uyw8xQZWtM3qiD3
A5Lj2S7SIsaFEmsl+dR8hN4eG4thC4RNsK9Yo+HB664SmHfjhZ297FTfJOCuQp7B
I2Sn9/3S7Tgm295jMfk6NL/i21mxZezGXBYtVc8IdbtAD6uhnn0ojNuY5VQj1nRH
IStl3S9X+S0WZMOoVxhSidImp6aw7yYEiKgFdGbuxSZURn1FmvPVnzDo38aSbYzB
S8Iet5Oy2sFgnjXcX3iJFodtW0bsXSHXhxvQVgqock8VK/wcwBDLp2haom7xUVnB
RjrwmJ0gLimhH26VeP3vhdEXX0N6votSdfZJAoKC2Mq+YvU6gcWMkPx2pmrgJrFW
UPssaQKvHt+zPe91MEq5O9lKyfokr4/ptJeGIG5j5y+6HmQgmvrTsbhGXk19AdFo
uswxGvMl2Cipk5fUgHqL5sBcvy4d8fT+mc4Im5+Ojjvq5YQnSfUDIAjARvzy/Cdn
Hi2vrVCS7EECC3XBcaEBC2Cm0EVQocEsPZey50FbHSlskt7jnYMkWqGFt2Qbw2Oz
I1THsyHVDPkQjKCc8cTtzHj6NkhhB1nVriUeN/lcaKADYjSGpnp38z7mYnrED3ij
CZyaDClpG3AOi3EtHmoWp45/jjh4U1udNdXvPrEwR4FC5mqDlcXeC6nDAwVCxFZa
HsUw6C8cLDiG9m2dFlWZr9BJn8TJBnpCXF3XfUUvxZe8pXVR0h7s9Dl5BdiyyXaR
hzDPxf37ZYD4Qdv2hQvyzXfF6V7MQtKQ7kLZMggl+08mtFkmn7fUr24xYueyyPAD
Vot21Pbgo1j8lhVydox3gO1vNSzI+DJ471ijtBXqlCH3Fv2/PXxcexBV3WpvCl34
H9b5gIgWEfNNDcdC2PACUWWnHCGDpshIqh1fpy6atNy1wi6GhN+FIodhedZ5BS1Q
60nh3DNsRIZCcu6cviTo0yJdvNn8jWBG/FMtXcU+COetMYQ8N6XdtvswxYfr3GqS
E/n7z2TqTR+BhR9ilO6/pAUtYMuNQnyQzRu53bKvU70H3gP2QlyHLlRBscemNrRg
QBm19U/hZ+bTBP+gpEH12E5ufGAqbEKAnDrsbye/wCb2Vi9PSKyn6rDVrjbCO+ue
8oPcO/i2lR+sEdDGmcmU7J3wCKW9pWQ/90LkcXdEys5aZRdoL1AJRVTzNEk0mnkK
tbAFRWf5Mhhj2aU6x14TtCO+BGo3EuIZyNylJTqOcO5yoRXExoP9uBS39gBogxvG
dU9t4MQ/Q6MH0gn3FeNU8kJDL4VVDtiNT6CzP4XyqbgZg6csCMHfEBdyZOPxSV/9
EegTp+yjnRiCf2rkDRA1NgD0gJJjSzBp3emLr1QDJJFwRQyh5ghOkuHA64uPwY5l
ES+xy9ebUK6Wpi57AyFuPlqTH7bieCOej85wKkTB7ZNuEO5eb3P4ZsZqfmVa8A17
1KYIsbRpJEoaBVo+BAaF+zUN5GKGhqe+A/Rp5ODc57O//lnxK2HrfYzTBkBAJmsc
DDPTKCCcykQgDNbukb7gpw0vd/5TZyoRTmp1SQP8EC1NGUjvII1sxXPxt3bIYf3/
x4wPGfVYZYdsPfHmOj7eDopkINDBV6TL/m4wqCm83PjFjl7vLncN43qmEM3rW7qX
rG9swNAx9bxAG5sqTGgUl3eSbXU24RpU7fkk82b40dYV5dAaZO7ZMJbbZ9PhwBsa
zpqdjeiS4AH1Zei4RniUheEqfsUxe4qF1shjjEgRWCm+CDKgbynvAy9DKDA827qX
FeoyxlJMhZj3RJ5RQvIA/oyncwZGApRM5CNwC8V/QioIY48JZGPyl1/M82etugQv
4BDDop9N4gfSLee9fOCSZPCzqHQgvdlW4puF6CU1S20Je+VnIY27UwscG1f+HjIZ
jB6bP3CF9y0fZKjG9D5MmTULqvm/w6sKw7wDYkzC8o4y6Vvb2jNk36Yxv2rr8eSN
qJq6zV/uKBK9CGKA0YdPUrZSeQxAqAWD0gDZy8Wp9Z0EZxMGD0TPcLfAKY0jkIPY
z4f4YJ62nhy7jNf6eVbFqRtCiMOKtuSCQpB/85b7/uxUvq/6gTwuwoONKtKHgDZy
pkx9qfVSX6g9s4Cg8ZHJ9EwkiWStmehSCuK4SDbBrKxzCzw2DixjKqxsMeC3otBV
dYf2M21ggxSUQsAVBJNTlmyUOc4+XIyH5qbouVNMebA00ovxFtrZjNuCOidby2pO
rylL6ofMWPrm1eSW83fZ1jFztoQBlo1x6fkW4iI4jzlXnTkACN7N20RP/TYZZskw
NuTX5PJJuaSqZUL8f2wr9411Uw+DI8G4Ls/XsocYjWAbhQXwrTe0qh2HeVoHHprj
mVHWEX3hxxTI0fHdVkDfTa7PzPLFI5Req+L2EW/YaZoqX3c83cmInGJN4zu4AZSM
aK7LmlIhzgP0a07E0eU/KLCMR3r3T0ZQ5LW4Ww23TcmFdPs0sHGsvu0V03Zelk3Y
5wDEkA7yO0reTci387CZCG1TcLPNYK+FyDPq424RVT1L+RbMHEgkF+JKXdjDAEiP
tYqf0RcXJ7fIJSVFuU2HmB9/PZeJpnW6X3hQGcu+my8/kAhrEfjL84ru6Vnxy4UN
mh1dUbdPX9gLZvvr4sIHnLILxzb1itsHN5geEjUxIFxbBnmCDgNCb8DTl8ssRh6h
kxcXF2KW4fxGU6WDgpG1AFBhT0B1nRpWReSz3EXLD1oovCnUib+Gja147mkWuGkc
wtwX4QcQICZGeatNqkonfYFr/HuIOGgzaQ0L+maWQjcjYmSnUKF5vZo8LbDDFzzx
OGeBhWxQSq5eNEeXONCRHIG3jnXFOVfCu5aJpPk20FYBFSz5kZUf3hkK663rCCAE
YVHejso6zrlP3nFjvcmJF64H7sgqzRYHO89TcxOX+QtKnrNC2Xsl2zyyPg899uGD
K6iPuORu7kEQCSxyiYPlq742Ps7S76qxa5wTHfQg1VeqoTyxi2PQ6YafXlbw+QQq
jBwGzF2qHBWm68sqiW+nlvyCPooBvnX1ViOCwkfNMEk27zmFttXauzvmLwkx3yPd
mezaHWTMSHnQxvPrY2ZCfcwLJB60UJY8dosxWXpfjoUBEdg1sj9HhGKBlszbJ4Ho
SRUGfisk72IqtQpMvIx0p9t3R2F2bRKNjS1h8kkwqMivEgdsY2K5+pyg5x6l8mn5
Rx8WzSD8V6T59OiU9WpRifQXUwIxP7psBMFW1c9QsVAAE0mOqZ5YIgVn9yS+K8Mb
AJaXWWLp7OjQAjcnoFADbfkRJlHcRc3s/zz5I/rQhEUf8zvXoPbPMvOdAgxOjoTQ
5BmgLuWDNQkxDtgaIewnaBn7HONh40ycRkYpix+3fqLUyWWIM2DmZaVzMoYpaFoc
1XYIgmdN+Xi9wbiuwlDJz1440lLcYi697UXHSWjhz02zJvfBUw/RowG6IOyn6BCX
rcoWAYeAEQGiSmC5KDzkX0FCXoF1a+bHgT086odGT2bi6aAMbBYuJNDdTmpM2RTO
uXImx6TVHLqvNjvvqIN+7nXdoh8VXssDbOWcAQ896d+Zvwik3qgSqVNZbgaiDhQp
pYFE89MYcydCJ3M5CykGxNk7DY3YVNZ4jI/6VF9ovtMbtCwoCnvCCCWeonM2HHGj
CJeiH0VpsPYpSSWCdU92vI2/61qIgLb5VEc6V/T+GhrkYWrRHQHfh42wyEA5cWkZ
ahalpquiaJFN6rdKh+p55VZ5/cxpR8KqdiVnsYk8C7vXmjVcep7/3fjKr+YgHs0R
47GAuOZtsnlxm+4bBO5nfoPbXTJ5lhrT/fTSI1VsiPmTXInDf4346rjWDnAUC00S
D/3RWCWnyFMxfYBQCpttyRfcUG+tpUuX90TEbONDFLA/UED9ZQyJwTHYgS56TFql
G5IjNYRDTVjvrX7mraYvtGXkjv+ZHqt6f5gwNPSwLH0wms8d5xNgTAjLqzKB2o4U
7gVDLHXXFHqybMDvWtuPKuwmewWWS/xuaAjEuWD8Amd8ASPM4I7JuSykkZxelKVq
VbMmhRgHK3aol3kc9xqotT/TMG3t6t4A+nkXvBfyc+23b8zWCJ3y0e9OXpBk9j5O
gOnnITuuEjaaSobw+oY+lTcJ1dFW3HrP9BlV99u9JIYfrlrDpeHcsQGo1F45gzB9
v+J2IwXvFj8fz9XYdQjkaWIvI7VMmdMBFAWyJqhQpmSGupwztFa1ckmOUx8Ai8SW
KD2o7cj7aPwTqnrQONSRURlwDVXrvdrJWhHyz9zREhaMrvzmkWEi9ue6CQnCbBSI
Gf25CNk/x30zogX7wd2paacz7N0gcEW9f/Q2N8GI1plpJMRbhidNSDBlN2TULBgs
nuMgbEcUMRkDZh5A++D7niFdaoB/r0wQzVzFyWcwOIxU22ZZZl++nGHgdx0rAreg
bBlnBHdBE/qtTA307WWgHBGKUb/xmC1OsRcsfwisHDjHZbmYpa5ZvjatzduLftfN
b7RvXJBRqUDkmJG8aXXZVNQ42rbSmhMIt9P1N8vRU6KVA6clcOnd9v5A6qTCKAfV
uUikzNWnP1A7k0kAzZWbhA0E9jRjKXJbcgp9LEBhm96TV74tDnkiHbmYH2CEUC4Y
lxdaGZFMNCXRT6+/cdRGg/4UbJcUUUImnQjELAzZ83glACLi3Wg7jBUlrHI6kK1l
aC3eIPdkTBCgsXuZpEUJ/CDF7hU9N00XwuHpkDX0Dpo6rfX0+B1E+sujwJqr0iPr
Rw5ZA/kv9WTGxHqGw2opjSqO+RLXxm+6+VgTO1U5CdQIUUGmESZRZYiC66zUoF/Y
gX18UFUsJ5NDHpJxAmI8UldN/BPYyks0pMWEkbr2wgjfxqE+GJUG85Q9fj4eGthn
l2K2fI+wbD1xvOI9y2khbjky+jbFdc4a5uq/2wC8RTldMrkCJBzoH3kV2zhBzWpD
NFL4a9n47qwO/1rnE4QKO+UMGgkcx6uta9jlEXRyo4RHufvzFY/sQV9EUwsQ7cqo
ciVvSGWVza9mTB0cXmLVky9T/XDO0wuDoXPUTNkkQjh06+30BDrVzK3gxM9oVP8g
1C183tRCI52aX8AKhLRZD/W0V/XUM9bQW9IPZ7XX/xwHDHHhXmqCIKBqxlKrg02+
8oVLTxTPTCF+HXui5aHS73R89Wj12M/QIVuMd/yAtXUSugWo+IRRYQ0uOfcqMwh6
+tiS90siFCRTfflRWK/o8v34FSsijzPrvNUuNKxRDSYiLek62FGw9uYyOoUNE1wY
bq9moPmjt8CX4z99AjyXmvZl7db8jnYyBbUQ0qh6BeXVkDMGHODODotgRATQfpyK
OJUNaDjs47XO9J8DFBh1Xt2JJkWeK+LFOzxEZB71IEl152o8fsIdifadPRo9o0uf
VC9EkB/fULq2uEf+ClRE3CVti4Pwfifr5/kwKrhbDFc+oRH9mlUDI/vCA2Q2mJFT
yWVlcpG5UcMexrfFLIyYgo7G0AJHWpr4DGza30IViv4/OIj3Uy/WJgRrTHgRTmXe
SwIFe+rzp8igcfWMUO/ZVRGNdQKUjc4WW0hMT9eZXMuYl8X1TEkCX+LOMxlnJAJb
x2TLE7In1z+UjjNOOclRTWTkRINJ9QYdtaKiiiBR/uxaf26ia4ZI5m/mNZtWJSYs
/nsXS3TiQjIqkx+Lfo0EtxSj7RoCeQ9ULWvUAMsBHfr7P1jVUQP3iaEGxroqvdt6
sia8x1NwJ/TDV6qZY7EiRYLWJ+G8N8sUSh1NF1LXOsjLHNsda0hfrLJyee/5iW2Q
T+SY4AKOG5FEY1A64aJMpAYhdiqBCd0duYva6XEKOnlUGB2U0feZkRRxzpkP00Iz
jocyWP2W5bJhUV1yjemB2VX4QATPC2wyNvQmNAkMk5pwyhzPaewsMzOaZmzFy79H
kdWawoqmJd1D8XZyXpEYP7AZsbriulXEqchLFcVfQiSWbAj6oEc1OBbS1/WgyR42
L2yAwMPZ30iwFdYYH69TlhOeBqTWGGeHzWBmGDNPp1EuP5Ko2WhKUgq/oFUJWUk2
DNnijFQEqCf1mq0+c7ZuRsvNm0f48QNZWf6y5LKMDwdId3usSw4uDTP4PC/Vig+Z
Pz325ZuqH3X4BK+TS8lUw+yYp3YaR8z4kdS1aRd7E5nTEiVpxh/Sgs6wnipTNy1z
HQUmmRFmeJNYPMy3dnYaz927yL7xfYhzKh0rAhVMzGD9Cr25J7BYImoOMXLd035Q
EYZMo7FYiyAPeSc7hZ9ZzlhALE0C+dXugrfG42EassOzehFxZggNPQuZjww/SpFY
a1h8otqXepi5zmodfXZ0ebyhAZlRcdm506YgE3jwoYc6j2Ezb8NZtTjzo0JRbjBz
kfjQbrIQ5AwpC0wZ8PxRTnrxEw554W+axsZB4kZsg/aDPDP70YMTVVHlO8HaM6w+
RyIhvS291DhUiZl8d3ohgquKR0Y52DnbneUr/bnkl4d3rrOv0RqSGiNqG2Bk14le
XTg206yMRNShhN1hpb8agMkLarNNqSHokX9fAKwuVsST3VWIFj0njkinjshvfPk0
4C9+HmtZSY4P0DyxEp4zgTQ/J9871zhmPSt8se623nCgeGx7u8asGEZqOhBZjoUM
cnhqOz5Je5CTvO4YKoCpAnE2WM1+SavEqCmxAEnoWJEVVwhbZwm3iIxWpHSbBqP6
0E0RKvhIz4ShUhehjwOzbzRRXLHo5qDNP2YcQNh1SJUpP64ImWxysLud0efcfuAm
cjXRHu8yvt5JG0We/PTuPbz4tOYrINlfrNl92br4BSS0Nqqo5cOR22GU3ugssyYd
rk21J2ETBpRholpyEmtOcnRdhyXMU9NK+WHP1nzXxGtMBtA69WymAvH9WmtvH2BV
aXsOwrlYfJBpJYoFH8OIWFXcSvoqPCQA4ucv9P5lT8TnoGcKkPqDFVo6ZP3wm+D8
uCrfYJxBe8MYe2eBpCBtK2B11KKxleQ0NbPszLkmnKXCQNe3dr7p8zdO9AZCy+kJ
JGafl3eojGRyMNe9c++lxykrbYd/Mpe5oBwPkTKlD6IrZkSZfxPcNQlGhlx/Ygbr
geGzFjxWTYzkqYxPzTR9PDban48SnDM1W8gF3637OmxvvyFmrkgWXogN3OsmQ8GL
jt5OiK/OgC/3HuYqgbvE7sO6B4n7Kygh8NOAVkaaHF4N8jrLZlRh2xwR+zKbN0RW
89Vc2kKWk1rhZLJ9SL6Neoa3TILMBoJEdSmZKP1/exlJhPICLIo0BJtHdTUDaAaz
bweoQH8cg2Ofed4D1O/kZnXqfaG7TYNi5nZdjN7thJhLd3fFsA8h2tLEob4jYUoy
JGNO6ATFzchw0YoyqbF+srVXLNSGnazqyrtfBN32Ji8PHHxW1DwTBJr5nhwjmdZg
9/swlI/dtuVA08EZZ7HJeiYfLzPuJT61ieedHUSpuppHInbnfHZb5mK+oJE2Y1EH
95Oh9LaUpfd2GL3yk8bK85oqj3ImDdqh3I5p6D4O38C/fpHvSEAR1ZSXxaiYGcVL
2HW3OAsiSWw/i4eztWAc5/2GRkAc1g2lSxEoBIZf0MO4xlZCKZJvTgiNGQjxBKu1
45hYLt4e4IxEWyp/TrmAUYR7U6N4J0+/DzXMwIWvqsq/IhMkyF36yedRwrsWv9qw
Uxqv4Wh7Nf93xfGNI+pWnYXN3yDmsgKGaDewDm+zb7uVrwakdVImX2oviUN+LMAX
prGeDOShvgptN0gRGPLdyAEkq4b1g5HClUZ2S0FHOOeqej2g5qfyHoTeaZJpO5ra
HPOE6VWs/AMiUDEeMz+l4ciP/+rkXmpfQrfbLTS4eQwPCxxIoxb1RGV5kK2Wpcor
oKDjCboencxKM/aLRHjz04ipVX+hVMeidZH8590k98cpeOL2fdYkG4c7hWMm8lwH
buyIjIUvVRwNP3JnAnZLnvRHfqlP5PyupXFpJY8xZqFD0l3WJ5hY6QmaR4VqP/uj
ZoApe7ibfP2rQp02IoF1Fves6zrkgzXkLx9hn+e/XAS3f4YJMHrJXNF2Wd2qMFPe
+QkT9hAMUJk1uvZSZvPUEVSXheqRZ2ny8D2NiDpm90GvZKDPQ/zXKSCRqo0xa48b
rkeM+WEb9UcxbjGXgbZF4SuJ/INT5QNk/0vtAG47lWOluvA48MHRQzQKxK0NCuMO
PsRocoL03kQaKbpfAkd778B+8j7Uz4sU/G4GuqypV04M1tsH41e0CZQFYexR70TA
s3nBgQ6blkeAYaAGXwJMsc8SWYJ1EEmF8NJwee943BHAr1jmIJSPCeYX8FQZ99An
Vvau8MQEkWyfZ/FCTZ6n0tTwNyugI5D1xzxE/ykrzB44jujKtAbd1J98hpD8vLQh
mpFgQSMV2zN0WXNxsKOC+uADuPG1UyYaz3I28AzfftY8IwZ96R0aLfpEqH04IJbw
IaBjr5h6sbx6Ik4VL7+Mr6ZD2vp/qXN04G8SfG8tuvgwX5viUvzhXbikxIMC6Som
23Ar05HnLRYNAxJrpTfsRagSuK+vKRvhdLhxlSjcmKpeiiYkMhGMwiRtgYC+XTWO
4FVcjUcH3u0icIXYJ/zlLBF9cQb8TSEZ9OwxJbnBQXb0xot9mTMghYGONDapVU8F
akWVwLY++oWMP95IgxebyndbNnswYC6HjTUmJGN85OqG3hmcQbctP3NHkkcFVTML
Sf6CYgdesmgEwEGx7bXplVFsYRs0YRIDwCOGyR/uR01Fu4fr9M7F7rMk6+kwILn3
SmovWi15+m//wmm+87JJ4VkO5sOd2F5QS3jRetqzIqdiovSKuqg4cWH44eVRVHwM
Ipnd5WEaOtG34DRWddZoC6obMRqcuprM8qZzvXD7YWaCbB6hf7hO1QKcJWotptVp
4/V7LiOroIA4h6MiFsIW0iJAJpyrJ13dO6cl0oUxtEa2K6spz/Ifq9Wjg7wn+Xbp
AKj7fMmBda1BgXmbqE+7ok0nzHT5v+AIVdUcP8v/QXFobc25XHmPMIQ+5FeBruiz
M3jnJwFup2wqYbAJ8Hzh/9pI39GrPNVyAN27x+wojCrUpM/gUh7kKR0bjCvs1+sL
IH3ehmU4+jXYeGlZKEUW5Ub5r5PTiDLWKrJ64YYb2CCrBdjZgx+cup4FNn38cpuX
BopmMdd0GdHUVQxbDLmDujGzSyyp5sPtd5cEMqDLxlcV0+NfLlTU7yWtuGVAvBaV
nm48i7OBwzK1+6EmGfmtdoI1gyIeC2iIQ/oiXoLxt1wKlfjlSn1s+ebmYDT7pYRg
qyUJ7f3ukuRi8xVAsERSGKdnTekq3F2Q4t+WOxUJgO/UDrkwqsyVsc15+x9ClrCQ
OnHmYs3q9r4k2gnAWm8jfKTCuFY8h6d2+N/tlbFbEsorPBGlTCDhd5nZeogWPTbS
I5kJRS+sGZbSKkwT7yL0YryAEbv0ztW5yWwW1wqvPDt1XJmGlInSstzlwZLe0p+z
1ooWfsHe5h1OvjUm5r2AiNujpZpkC008sBSPPspJ1JmVQ+DUxQtYFH/PcVs8kpI8
yyDs2v3ceN9p3eGUHBcFfR5ESVCT5Qbgjl+2jkzAexdpkWf+YE2Ac9y6VFpbns3M
Hu+M6DVC2IAc5IpAmsOEDKvwhMFVuHQUuS9ScHqU+ite1HU2y1O7KZTm524ITc63
BhyNU4sWoM3DQOlh1pyH5qq4M7QJ79vyn6PXKjnfqYZ9v0Mgqaml7JJX9GZlhYVf
Tv5kR0u9xkZq7nwpl60H7fWsFUWUAZ336TpS7g0v/T0lwq9j9OL7+akXWDCK5HXv
QXDE5qvMghPrP9BmTmoO1Knr7hROHy4edi2bI4mWHPT5hxWrVJZZ7JtH9YzfNgNT
wPxF0hy3r4AUJpvm0wQkZ7fmmK5s6zRBBWxQGhRrIUTj4XognsFV5N5RQQ9Pjq8N
BDvkXCOVZLirt80MhWIPFfbFakDxgcQSoUd4nMrpX9noVC86CoEtLdWOyMPp2eH1
d1Uei68WBpOP2R3hDlyPZwczKrOhVLaN9SUNeD+8SOoB6cjQ8x7VD7gMo7SzBb5S
6YJofnc2eMTkuJ3mOk5yw07wHZmUlAujwGYQGh8bECl6dClKVo6WravBCw9QCuSS
O5GSV4QhMV17naaeaOElaXZfWOo/jRLIv1aw4rzXTdOgEoDH66HBEQRUrJEsd8U8
N9CggD2vu4WM0gtlPRFQ7OSRD39G34HGprUwN2r4LuFMZBYOik7vzNLmyn29CU2Z
Z4W8V36T2F5S1LLnjdBpYMtpxgFlKG4RHPGSi/NN9PwLwet7FjnvISkWg6rznr1P
gCducZY073SVA6XTFyAHBwmRB2M4V+djsMS951V8vVhN55SB3A3eHV3lPIWoPs5u
up3SFbfNn58I4n45qj8RYfIC0DxX/6B93EuHlHV6gAOHVSXcQ57nw7ByWeGzoPWs
dKlz6LzfTHoWNhops8b3pOFxyXyfQXQT5+B0a0Dzj2pvlqpBsZDAVGJYgOYfvh40
5P+AcZPVldV/zfiCWjCiwaAtAkK5s/1ZhLIY95t1kNwHKq8QS+UpR70W/w1AO+Xv
OUBH8914c+2z9EE4CbTmldCiG9NEAJKFImL+l5LYzxpDLx0rfTe/EJ+Yc82uEUwE
yqubxZxQvK8d4aZuV0jRu4lOag+9xFnv3lwlGzeZ3oHvi0CvC9XzLepBn6k6FSLk
RDhBTgEprWZj1U/CESR4yHmxqHnWBOId4qnRm5efuckPShJvN2qbsr3Q733nda5F
ojtZ1pKG7b7DpAcn0sDjBgdjHgC7BetSRAucIceimk5MVjgdtaivab98WBMcdCkN
hJ2YK2jaTnmXFgzv5eFYse2roQF9VU0M7qqq8xSyX9XZApGjIkQjjk2T7lJuhYGU
j7G12IrlJkzVSC1bnvoN8goIsiNCR0zUHhA7lTxYhWEPRGE2KuQ7xHaNTsAguZA3
WG3S6SU98dc03HiHNQBaPE+kdUXO30vqQEwOMiMYzoKqmAiiccx0giIWKX4Up4gG
YrqGekM6DsuusMQJX+Z6U1qio1H++mQmx7Y9LIInuJ1t1HwI1bM+eVyPesV4sArR
WO0uXyl4bOYVf/Vi/Y5bC3g6/ekasaUwv12CSFAO0vyviViioRlWsDlC/sTFgiv1
Riam3CUYI9O9ECx8fnPTmO6QdA7YxVegEp4GEdu7905FD5gWeeZjbb7gBwW/kWXc
E1V8RuX5ctkYBFf2WQ0kic8ORDRLKmniDkdBc3rRMo2PmSQIhycaaEoEw/wpJTnc
+v0FOGe3rl4aeShAlqgUNesyffsi5vJWGqTw8ZctNr89A3a1wgQ1QjyYi84U2q16
Oad3noTwYC8y7zmH8kYcUZ11c6pRjcVUgrwp29hSCngovEQJyDf3M/+7lqmIJVYj
cP2+qdjKDawFIMk7IFYt734grG18ygR5x9x0wn+Ax9vRexYBcx4W3TI4zXBmmKgc
Ap3ZPHwM/sWIJ0gyqXV9kKSChY9Xx99P/VjLlZn0d5CWtn6N4KMf1nvIynDHUn7C
fWB6/eucMR3b+Ab/GERGnYqJNYfd8LfmxYPdTfPmV+3Q0vOYj9OEIBrTxbmcXtAw
KFarX642Ew8SdS3m3PlPvAMC4N/LHx9SajdSwOCAensLyjXc1SWdNWv2Th+2F5WE
7T/YqSZtEVrjnPCVjyS3+O5KkB1ewZnl4+YK/CixrsZmY3GDYzBmpjlveUIUZnXM
AMi8VcDzJh1hwvVjE+edWm1ugKxGmqX44DYpe8Yq4ocWjmEpFJmER2sPj9YKyC7j
iFApZnXVMU+qqa6GYkEXCM9cXTi5n7KhM710nI0bgCBrPCqsxWjMxDrb/VKNgvp3
Wqx7xQM+uhw4SytdOsPR4qz55ulO5mnMxVmNvJLBmUpq+7c38h1rtZWdGTUzEVXz
IaHCpPXd0xwjXZajDfUrTaxcxxY7xUuhqQAbJhklQRxpsHzc2LAkezxhg+ovEDwe
lYbkx7DWswB9AMO7sH5YBwFzYNIqN5iDTtA0bPJvP2o3AEOIqyjA/6a4+EnjOqKX
QM2JsMpbWwFKgkf7uth7Y8CUm3ogkcL3P9ZaoWVu7+cFubmGbvk17aedfUN8aJTB
ePw/oioYLh6oDjinAxWHBexrj+fteyBVgFAabjELphckiSQOLg1tGgZD7vAGOH9L
pXSBM02QXGsN+np6+QRAipDHLhbYv+x1L3fQc93Qwzvsiex/qYHd4dvg7/ovRg+5
VUZeTvQ+KDeLvfjc6yVcrVfcakiNeFozMDeYz4qC8JF/2aFW2jrzsGsYIgqxwgll
8pjfmmbOBWIBDrA9QQNS7XhezR2LoIq21cO+7am3kywjeRBs8X0bmBbgcd7OGHLc
BEZ9x4PUoBcbfugV+kNmOUEb2jAnMSMs9u/UzByWRy3jJyRo3uRlu9Vf1siy9OBs
sSihZZcL9l/rvHsXwNVrfqp1Wo+MTVyomWB7qi1AopGraVMCCPc//pXqIBXkrS5g
lkPjaYJFxfI54GC39PifyfbT1h5RHYpY6DshC+CKP+MoShYDhOTUN3RV1dFqW2+l
FRrGmQ7parIPdQ7L+pGFQ6H6ppHCtVi3YPktJs3za1WZzTkJA5pC4nKxL6rRN7k+
j78emkHW9ShZ9bO7JY1CULCcjPcauQibvkZ9rpEMwpS3cCaW8dDhuaV6aR+ziO5X
Jt0lrGYxzp7R690VQ03rV8Je/vw8ArQQ2V7zApXdYDcNTZXtsa06+5TxJM87z5b2
h2Pav/h/2kc9E9/Eoe1K1orXLZOx2BpMKlWt4gy66l7HS5I+/WXHRHUY+R7xdqog
B+1DW8JROIaAkJscoSw8jwzsOqiIhghkYQy8RrgLqzi9vk5rTg0abWsUtGveSrpu
GY6K/R6WHLknxbNUL10okz5Z/lHvcvQJafaqKBSAgCjqfJhDdrblxcqTGTj4TiL3
pGffddU2DLW3q2+Wf3Zu2GbTzhcY2u5kFsGNybKL8ywph0JvC4XjrBIeEbQRDz0q
49Uq0iTFlwbWHBxEq8eJ7zqLndKyf1yF2LFIWueXCzRB77X+yElrL31ZAoF935r5
64zUW+nr3qXLi2pbnwtsaH3gR4OH/MJm3+Tr1nquXvMsbo8NKwMFYeymLzjbudy+
zIZq8TrAnlrc7fGhbQWJVGZxgQNEjWyLBb7cwUYFkOiLYzZiBfdTPrYI7wbHEi+D
/3YPMeAY6d4JwYIXlaoTHq0rfbqFY3z384IXL3APEV8Rpo7p6e1dtjpYjijREgzT
nXnP4vNQBFj1lh82OO5TJPJqyDxSSLtsT1rwJeenGCbyaP8KPPBS4vFK31GTjHkk
zR0frhntIDqbxW4dTPbwjxBt2daT+y62fJBwMwKQoToHppxP0y/mGVZjlyylg2wv
dDuPipc8gTFVFk63pPMp/wW/ytn8gTE9xObVWFevJ2OXpoGWm70WG7p555Q8rOoz
UhxnmdvhUYU+wUW89dCHroUk8mUoj6ooyjc5AMI8+BxOiVCEXFibakf5ls3+bDF1
0WY/4ag31B9XrsZ4xjbaAgROQCOy7P6Olet+hfC4omspWvE7IiAivAVfAsPJxOJP
XdGznPgIMdAED70wrRLK8SVYGjA/NMTTYJECfPG2sagk10CxtUvDbgCIbV2hCbrt
foiTNp/lQaVljuXuHQ1Ez0KmZ6ZsW4n2yLyTAgw4Z/IcV2WHVhMmIZAYn4qSkIuV
Lwx6jFSaWpMD9TP8sWjLYFFq1lvf4HbbaDv3nJ0E5lhlTHGjQI/m7PaTI5Lmtibl
1/MP/qRb/5CZhTIdL0uW4Tb2aSnHpsUGdbOjgqivBM2BBW2YXsJvxaRdtunB9tVf
qsmi/bmZkBcvDN8y6ioAvcBhQj0x2VRdFgtPXbs0T35RSVUueRhy5qJIOGwYgNKh
0/X9gjKC9CBPKiz01v1YTPXEGljMR6c2DXYveDKQellwtu9ELx3KBXrNCw3pems+
4aJnHfW6LdGqIvRfkDDtf66IvHadNnmOPh+jEfdjT7TC9Geae19231sadWvGoob6
Pf84RvJ7MZwOJivcZpOg8CIc7ixmv2P0M/C/mq3JF2E5+cWtrxGBmb880jhzFGtg
h6p4mQITjCsQtEHKJ4mRnXfEK31qAbV/RkIVK01OJBYNjPxyM208eZaRyEEqZi7C
Hhz5WBpHq8G9FH2KLEAO+6iNMuydX/yGD54hTZ9W0dYaKInbYUZQTzWg2OTaBRaq
rc/EQQ2fVmWEUeZIZPK71eY1Cw/oa6YaYjzqqA7pMmqgbghe/9iihMM1xQlTBHLS
Q3Rc+v/iUm98XGHQY87f4ydqDrG1XQrE424FeKKehwxyk+f0liNldiTAeoU2brN9
S5kgLYvqGh+gKv9pZhEzAO9BEhJi0HEODFXyXpE39w73zmqQEVvLq2R1omYld/tR
yN3uV+KeMSeUhMjx4cSeASdD40a1q0jx2Dn7eTLkjtZQxEUP69ZFjLWH9qWij6MS
Ssmap1vy7iDUpEqVje2tqSztKsV9bshi20+E6fzYzoyyZs+nDd4IEozy85vKt7L6
fXKuOcGHM2vDq3Uu19NOyHrcY713+l8RK4Y2Sys4zJ3Ypn20VHO2yx4erKTJHXF2
mgYp6k4yZ6nBQoce0stbWuHyZlxxvp8veY1H2o1DzkMAVk5MknGjOaXoSf8urDry
8NbrNS/Ee9myDckWCVSh7DGojN5hzpSk1XwwXdYRhqD5SHUXGMEYDRGdRZuzYtY0
7HTk21INRcT1bU5dT6M/mfot7ctkX+2Kygno89QKu6NfwFzMQxwmyn3h85UeUKju
d/f0UcxsC4ZMjxvh+647QIfCQ0SLiVp7R+q0CzeHysp5cA8AsFbrqJoeavyTcorq
gRR3ZH5+yud874QLJcQlHStAvDKBbgENskENnA3EADzc+NchTzlsYmSvbZQub8O8
MoIh+dj8k+XPC35u61gQtd7zQHedNl3ETMzVNo3jXFqbe5uH/YM36EKzjw9VTNbf
J46fSgn3ojZOBM7DO6F7U5gRm2W5YFiYK96xpkH52t7JRipIgZ/8NI3J97oF7La3
6VyKJYuuyf5xITdTsYoAuJIx6pavNcWccmQ3W3s9ahZpcmQGMv2DiflvF0WFuYXJ
qLUPE3VDj0ikaUQMMrgVCL1xt52RPqa8KBLq8v4WzkDyrD3/MgJRxiWqCSkRsGNV
G4Fig3q5kYffjw5YJ4NhF/DxUhB6JLkg7KLuspzo+NcJgH0Tbvy3wqadZP9Led7k
g+FqB4runkISyIC/cLIhyndN7+CTCOZheJa1T7BLlGbOsw1gYtW/qm8W4Uld8sA4
3ob0swBAI6vzxbXMdK3FKHhhn0FaqUZHVxpbyKfJMTKDZoOgZcMmDodxp24EiOiR
9Nmxw+YU3HZaOtvBGbyn4yP6ZGPzCHYOOMsl+QpmdiVGHp2jD2LEkMsDN5zVq4Xl
XV0UwN87A9uAsE4VaXkPjE/UTQwa0VTHKEoIRBufrdgIaBhA5MWO/MIvKYV2DQv5
azxQ4fHcBoyCFSN3xlWutlJInBjrfq5JcdprLkz6TeVJq1hNqR8vAfVXTtdcUi4l
JxyYJFUW0KqkLw6tt2A5YSxjJfOekpFiaYMUMNVHLrpGw7xx1v5a+Y/a5ltctu3i
OCQop39v69ufBgXhWwJ9dSJb+4WvIRbWbmeRLSXjb0IxyltYL10U7lqfbNkEWaCY
0D5q90EQyB0pLsKhadto5ir4M9xRaPYacDMNuMcTmQ0NDlGtYbnKOlZXqnkM6yLt
eawe8VW4f1780i7oB6z6uNqfl4h+OB58xiAbryH6SbiAAg1hV+HK37l2+9PODyqG
WUDa+mRAhf6INCFtKjjgDc3v9f3pD/WLzfN8Ltb1qwnGUtq4thv8vQPt6jVBIipY
SmsguantitUfSgoDav8Q+s1Q7hGhPIcsRl7jjavY9g2AYYnu3laLx8vISC2Ar1CP
nTLd32p93ekr0Dad98K836F/kHPshV5wEcsnmJmtRjtWSwLSYkptG8cKcSx5QMGJ
SQqldMDe9hHJLzYiGh7/LcYBjDiWgmv4r1BpBvRQ6FuwPgHPk6qGppTZfqGdD0TQ
dYxhaQysBtcE5rjnhevmcPJRy+3qLledINKUd6hfFWP4hSNgupk1pa0v4UqxFFYB
EuFh82z9TBDQO5LL+vBSk/lBLPG2alEzF8xIosWAZ44VZdw/NHDiwQGwwOobGIPX
rZTufD03CQcbCF+qZGqVBoq4Za52YylxDNfUJCcMfLEZmhlAxVIL/PgPFCz4LiUB
5tEUJWoGjUi8EFd2yM5PQKQuUiLuXH4WmCweJxFkBxwpwo6C+4CxyKd7VcxO/zJ6
pOyyHp2Rgq04Tvq19ZBA2qyzgh/Vvd3Ln67jhbQWaUdkKAhqklnZtSiR9qGfYmty
LuR/Nd+LtTKhBqjDT7I1FyaU91kJV+2dC5PgFzpuyaPu+vNgzlA2Zzcily0YWSj6
kUTOojFbZH7IttvYfrkmjvo+rtA+Ru7iVPkqxgNYXHN2Nof2qJp4o/TpiNGRSJ1H
1h2BdDTgGPsr64VOMzSYrWF/8QtvJHKHOoV6KbRpgY2LPpzSNQXZDOz8xPMsx6tC
UtGgSZXhcm9DGLj07KVtD8xQDH3ymSswqDL0lAbydVSx4XHtxZA1l7lzVjhWziI7
xl/buTFQSOJAFuyXlqDlK+d8EvG++/pDv/702b3TwVwCRY4ZY49BORbECHshKrS8
aMm3JpD/uOaK74BQnYukyfamTvCr/AL4b3uOPVcpkOiwt8P1DpUdwsriXLiqR5Ke
5QhLbqUF7A26hocrFwBt1PP7ZsR6OFhtKiK8MkDqz89MriDRgLVlFm02i6wQkeUh
JJiwjIQJZuaM5gIf+xbL71p1EnL/O3zhzOagkERw36qLY8EJlRx8HZ1DkuOMLkVC
n1K6y0Q4YLPDwNT97Krx3EdtB7N+ryWbmICRUJtP0v5Sl/r2xmgENYm18UnOeuLY
7lTaIGLdFpdJzGGHmD6jlUSpyiDMfQ3ioahTXGXaaK0HVtpR4HC4Rc2j93RQQPbD
YFptBtap/f+AiRNAtolqlE7O6nGqTnj/n+aCGL1Jaov1bPYB3H5uDj4j5rZlUVLk
uLp5uhkInXNbP4lJ06fyctHu/l4mPlue49/kysVddmshIGAV72yR+xSgNu9UMlo1
XKyhlUVav/VwWpPNsAd3rDnZHEhBL3BVDur5FEgTESVeJYRINAxieGflVoes7cVI
ppwNcRsONiMWIO06Yk1RqnzYQN85wSvBKuDuk29fi7V4x6FVD2dFv3+19fRrjvnp
jpXfTIqrjfITYg/s+S8AqqUlHijCgGJsYC6grRqhGWA8TZKQ0s1kF55Iqq6EKwDC
ExMZ3Gi52aiLGMj08bF58Wt4PMR8vPBC87FirwJag309k0quqw4lOETg80vQC78H
dRS5yUlB4EPYWlHG9cF//g==
`protect end_protected