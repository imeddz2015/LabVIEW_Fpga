`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 62656 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/59UwEX+aE7FohaWu0/8IpTj7mav863zUNIsgIH2BWb
UbfsOuHiq8mfytoAtAkoScwHVXfnjV2F3HSui1CFatJEIrJuf58vHXQDUFCcgxl1
FCLoMYyb6NJsW3/hjbMvAnU7PGbvT/1+D5VrFazCFJ8MieA2LKVVZN5vVNyxzOQE
Qd9mvYROJUaB97u9rqtKpiDzhibz0+egN/mD/1cKR+koVpRdftkpZB07WKJzuJW7
8ZsDrDPHnRT4BD/0OlW70aS4Iuf5h+wYWfUeEKcNYLdHfAAy1Vr62aaSLwUun7s6
cG0LYNmXe6xfdSx8B0GgkWeu+7ip90HolWVygBytt/82FHI3xo+zmsfBEpGO6Ne+
JpNiowVvETgr9yfGepKob+xKbuwvU3jpq7ZdrB/TE4DiJ8i6ueYUAo07wAPh5Wh2
3cYgsAM7Ee8tdmhqkXdN20eP2kcgR/lnVlq7mnmuDK2JaTAidXjtSGvb6UH0Azk2
vZ4uklftPDrSza/YImcDDpuF0iRsCVllLjV4ACf2zz7qxp7DvzkhrxeHPz6GBYai
ae4GchwA6cWynAN2Q939Jc/6MfKe/02PNlOAJRYDDwAkpcWcNok+0j0c8VG3Ju2F
X8I2vG1fTk8Sh1dbuwwUgla5BZBnzqUdna7yp0FS4sl+bfEPr+Pj6bUU9fsgywcj
HN7jfCYWist6wsIsI5ffGrdQoQFSMa3nGLU4o+5vpzjulhfqoHkF9qI0fQLeAPiq
V4W7ZrPxoKKKxoKg7DT7p3ClZB54H+xVr/rqdKejBw6Oe9YqY+cFwQELOtECO9Zk
OxvMGxiG9QrizqoKz0Q+nAenkeO8KOgOYm4u0QYyUp2fn3FuupaiLKfJM4KZ3+qL
TK4cDRtY11u5tgEZuC5kUjslG5bu7L36ESK+tl8JZWzCj/MeyCoo7MFtDrpAv27s
XsuGXkHPQoI7CPdcV7gRnrw8ffUz5VtmDRpxoC7LHP04APzfNt89dfwJV0/4kwbv
V/6YGdvKfLWF5MmQQODB3rnpOBLF3/yi0Qxy5zj5NfOfLUtJxfEWNcqM0hqTh+p3
aSJKMFRXNQVmJbAUqAWEy9uJuWL/tk9aEtXhlkoGzfwJsDuVRQ57T/csm/6WZNjH
3FhqWfQeKIArlbNxk0ygnGyLag1UVbuf6IdM1plFQPAzAw01queGje3iFhlju7zv
CjpIRqATD1nwU8XiaYTfUJy8meemj8u3sxT16ix24O77cYTVFjMpfsDPbfgWTL6f
LifZ/mNFDBWBoENnjQN7/fPG/fIxisLh0pMMqJcIuUFxHMkBPFJzeqcLjqZpGS+Y
GmhpIZDz4vPA7kjHcW2Xo0nzriPyw53PCpGC/YFf9u0AEI6Xal9M3WYyNXSDidUS
jVserWxMP7Iy2ptPjFAIFobXbiQmL5u6nA+6q6b+tWInicgv5r8jQ8vst2NwvI6f
n948VVskHLHullf+XpfRWUPksCR3LbtMZYE7NKxZG9NXNStYJZPyfsPPo3LbhlAy
E98jn4br0B2IapytVs5ZXH0NWq0hUTpdwYk5xxJKdTcwcqJS3aE+KhGOaUx2Japh
43Isv5rrlzLnDhbJYRBV+Z4eI4N8zUTXUHNTBexwTLwbXKmwuCgRTfC1DRO/PIsl
UDcHEu0Hovzua/x36uvj1kawrbVIfSVnbZ84u7ioon64owHPpDkGaVc/Jn+6ihll
vmgYrM8l2XhAMCp7GZlnVQksWTWAveSr8tMcS5qh+diNhXT7NznxPEoJjn5WerTZ
1TRbBSdKZFjoJvagnjJ5imWvwCw6NECtWMcUkcpJ8VPyqETWyLyxEN8PTb4dV4GT
tpz5v4jvKuNHY36kZ+7SkZvP4n1E2DkelT/DS5y7403Uud5TOuASvHddcIX5pksa
0yAmPB/7lYBXRm0RfLyMW2jjJ1kei78Q3VoQka6JgQNoZI/fYMEY38E4JTsQLv1N
MEF5PY1pzfNJykQOicgRj+/7eiUPDihKASzGgMg3D0Ixv+aEH6OvW4JBLC8nc9yH
f215CUeTTLGB2oXeje4eLPLJQi4Ozz9O8LcrzHJLpuMFj4ZwW9DsiCD6f6pZSqC+
X6wMpf0/giqng4nL/P+oqVcTGTWSQT+CzkzelZHZd0EbtdhHafn7RPrmMwtpDbEj
OsVOOBY1jG+/6ttABfvONocT/5R59lD5icOVSELn468/yxp5RX64yrC0Wwdxiu9N
rgWzZCWTNbtIMnOs/Pw6+ylJs8Egxip0QBhothb7Ie7ddoNFJPRolzpru9AWYxtW
P4U5Vc9PWOaexefDWEg9joqBOVsni/vQRhzhEEqdBCwRVPCD0LdEiuFTLLzXp013
luESHT8tTcg2TXSr0EVnxMcHFC1oyyHpF5tjju1dRq9pevC1Cu2kfAO5BYnBRQhx
Kz7yjOHp34tgrNlEF8qxeRNzeyay4H1z/BsgwvHkqd9wJ89HkgkkhbgQIIrIpCxR
LhuGrpizLtoAY9thXJVmqLOSrwUUVQ3lSkhG2KgU8qZG9mwXhjP86QR3BFmcdI1Q
Cko2+ZC54ZFLq7TNIK8fYHoy/TckAeznUEQlP6SlFN/i55gThuUdVGiRZuEfpAEr
IfwHdkTetcgDFduKVzBJ3ZByRMYdBdAcnZkRVsAsmkQSWkc3nXJesHnLlCl6K1Lu
nsuYrSlFVhMuruU/dnt5e3K2ASvqQB/DsGWsZmED4/xfW0kh/CD1d51BSwKNMi08
DNchKRmV6xg8PdHnP4+Abc2VJ+7QbuiSsY/lTVaB+MXla/O8s2xaooWT7rGWM5Hd
gkeNwCe91Yxf5TR0yMVWyR+JleosCjBwzjTXPvkKkVfeo+aiVRD+FxJ1EmdtB8aP
BWHiyE7a1BsptEo0SazLajgToR1ppfv2ChyTNHDiCq2Yn6kQk+zCnUke852LRb9u
KXTyOgjqVBrPyuqx540nA0pRW+8JAuloqwv4JexJZ7Bs8UvH5sxan45NdfciLZ5r
Mxo7Tze/YLE7rbeMDvqNExdvLNjDwvUk4sYHc/Og159Vs5VWQrYNcCiNToFYo06Y
44vlwfgyXuDPp3f9smnZThnkXFkYW5Nn+HAnI3dlyuCtjRLLlSUbrwh/oj6FWeLT
PjyFyeB4isCHC+Oh5W2gVFyrTdyko6M4VTau4ulUnmEe8RyT8OLyi2E9jDGB0/cJ
/ugK+Uljt3hdNa6bCmACdkBXanrYVDAC+AsYOpiw5Et4y9Bu1lbGn54AnkuQSmGx
A/6uRaREw+KZi63YU5x7TvPgTOit/2GpVj3iu+t+yQX+N/TbkN0IdfCr4d2FsEjy
PsvkYoE2d4jxXe+nURkObUwouC1gqhCoInGKPyoelps8nIvClDC3VAoW+H9HW8YM
Rlgn4Ji02vS5fOGSIaxV8IDJWg5nQBC9MhRL+vItmQwTrsY+Fes1Og2Ny2XyGHT7
J256Zb6Uu4V4eQr0yk5NpDmHMC63Ou+nbZcsCve+spL8egwv/7iKtY1p5wxQjwxx
3VjL8aTokPNkZ6PBTRPY3Hj7HJok43JPvH00CYL8dPP/l3tWTm0lKMl2kmZhlfzL
S+cZNuozgrSL1g2rOXzpyjCUEplRqw2m2d6pvKj5+awKmlSbqHlfdXb4gIevFUZR
4tV0fhmQpkbyzC1808cbbaVVRgPvZrsLDc7FzGXwN0PCpFTuSegQ7L1u4yo9WfA9
Cyfny61t2cSI6uZ+r3T8ipj78C1aLhKkNgs+umlMAWqFk5pKWHUlxMB3VZqXCHfc
lOQl0HqZ2X2Jw0vsgKwa2xZUozu5l+EL5X/Tp4BEd4oLwxoNkEVFQZ5LkUUNtvlI
EYIu5wDvBQjdzK1ZdtTvghU+DwpBCZKViTtAJVoIIDEKsweiGNI2qwZODR+VwVfJ
NBUwgVMvEwwsWnvkonPbE4YluWp7edi38erH7Jm7b+530mSlztl+ayXGalaOZgjH
GVjT+o3rxGJqXShav3MdYFACH6iENGrxj0i2/mDTwuTamAatBp21atZovq4krdYp
Ff0E/OlBIfy86/FOwyaebGqbuU+GNHJvrNURq+38YcOR9BhssYAjvW+S384XMNSf
LL/v1eIrcYbM0/f7TUxCAaTDDc/HSM6WaD75sfLEuaI3y0eoK8rVAttT9Z1io/l1
nenZx1cm57tYK0JH1z7pEXtmKeTm5RA4Ut9yJXq3OEBUD/dWuOYQMoJ1TipjBkWT
ct7wgncuxl3j8KmlONomLmEPDjpJw5kZ11bhPGmJaOCdLe1DX+tzKLOCqZ9KdWPM
8r71JP3woWUDdeadYHxTvnXlsswLjsjX6J4whMlOxwpl+0gLaW3FbVp6CwgiiCPs
fFwz30RNf2dzC3TAlr0bwj0Bjq/j7Cw3st01LR12hDADDgFhMxBERxTzE0RNE0zD
BmZNENEt8os7iVNGQ8FyZjBNf3Zmddz+dtW1iQ4TbHFfPr0U7T3I8fZXDJgOG6Dc
bUVmncNJU+3QUD8QtYYbqrFR9fSHkfDA6arqLv9oeZRbpxpzCCHZRmZ/Dhwchyno
eF5xtUeL/Hxhok3kofR+NvuoboHW4GNp4eQDJXjRMw7usrUXQeYpHqw6HHeQKeQg
5u5WKXaytVb9/pQBjNix/6d7Fj+3LbQN0EfnQhElrl+fNBQu2G9H3rVrlVkkuC5O
Ar41WbBMdWuV2qJhjcz/b8vAff9N9n4NGBEUPZDkXGE/v+9gkYkoy4Et1EOrN6Q9
cD3zecAlsaAR5Kv6RpQGjIJED1kHqe0dY/2HgdY2nBlmIO/wVr+KnlGqdzeJCgm2
gU6LhN511wCvtQmv0lo8YAp6dmthiuqvdWkEt1awERBmyUXJpx9aRD0udF/4R9xH
qj5QEtC1NlMAHhvlxl3s+iqRje/9A2i736peuiHPGx/UwsJ0ItL/DuQiNRouehjy
8ZyC1VX5l0iSzZxgT6I/LTUIvU9zFuYtxw5sHZS8srxcjGWwmAPxFiBgbM3RBdd7
o6uPUCN7npI9PUN2m7XVYCX5J+J23hZirqkuclqWUFbIdK1XZaArW0eBxsX5zxIg
En5Ij6kwDE7jWZmwE2lmCeoSY8GwVHvVqHx7ZDzu8u3kE92DEz0QHLbUywA//+fw
UMZp9UtCVBHv3KYDM6K/ZXwynurEpJXCe8RUg0K0uBGVL/U2IeQD19SPrz818qGz
XEUBniolOy7PjskbxKssSEVgYHcGKYSeYYE9i2OixFiJBlbt8PzBPn3kkt57+hr9
KDGID3ZI3U4beJ3cFbPalzGfAbESvp7lcvgtVp2nSbDBnjWrlB9NuPc+QR8KjZl3
3GtP0j/JtY12oPcdPfyzluUbAWf/Irb7kYI52YmVmtBi6UAysgIvQEp8PMcCPtMh
jQp7tnz0rphYXHw0jjXG2ljSai09dmEyKglBFJzrtGtAOy/oFs6vQtqp3bPKS9Ic
v8zSLCbj8nMTL1ZQyN+5bhRcPu72A2sR0fVROAsG94QFcBNBcENaeCy/AZkmKbIX
b78SAdVa/svsrprL8oBGZb/oRGBR3ex1L3EhSz9vxpBwJHk7NS65ja34YxW4ENih
x+m7KiOHarYmR/JwnrF6iAd3qNyInEUfrQxBaHy3/ppjNFCKvaQfNDWo9NVSoI3I
U783yPJDjTZLC7b9h0EBmB0/JdcLGSYIBLRC5MQsdPTLc3eb0WnaVN7yuS0Bgaqc
FprF8ryI0dXHGUYQH9oMiPSQicPhxZRBhvxiG/S2uJCOWIo1baUAGRAkl0mOO+bs
mBI66yQp1x1pnCKymLDuOomOFt8q+kgetGV+R/y3Bd9+5CaHbwlGkzv4g8wjvtCT
tIYZiz3mvtXARsBaXBhM9XMC7rXRTN2B/z0Rral2oUiUCtuNlne3mtkMgfAdBSk/
pB23xs+C8zklGy3FMQauvaqnFdtCkClUbzQIW1oGTsugohs1aXh/MrmsjAotlSYW
TgRL7Vl/zvP3Zb93ErclgCg1xaSwzmN+19oT6HHS0xfuia0mJyFi7+xn88NRPfVH
EZEzV4CJSQ4ZgK8G0uLRWupV6WZw4N2ChP272pOLgnND3iJRV9HC7xIxmBOyWXe2
lhxi/F6ZNoNFQ9XP1H+S49djKgh9piRxyEJmy7ZzzE2MwwA7BzYB3EGVJHoK+Fc8
yZmnPSxlDTb3938Z5t1PCx4rCI6JRYR/CHB3Pc180m7Mxo5ZtcmvGo15TelR0i7B
D1CPTH3eNYGh3ro6LfKOi1t3MMTcOzGHBTKBYeNYhwB4UhsE2eTEjTbj97ISYmlb
n1sq8V8j05g2ysbTCQA7JD7zdoNlkj1qZSuJsfi3qDN90lcEc0gX2m447aMls9vi
6JozoLOQ6z83QTOo4LRI7f/5ZVDhmIJ1KHwjPCv8MPh0WjNEXZuJ1zsTfI3qFePh
T5CV6I4MDHsJq6qSPzLBznLSOgYmnpGGWe79lhl8XfIFkm23x47UukmjWAFgGUus
hEJFZYcFIqO3cvDJZuCq7uwVM6+2fzaqLfX+ZFhHwWh1Os8+8lEHUQ8j1wSPWq5h
oS/30go5M6OGb5Ueuy9baKGpVWBf3apY+uSldlZiP6MyQBxPrhEn4BhWQZ7Hin8m
IkQta0chAqA4LVkCLMXS2hSz4qDuNQHsfyZLXbxqPUiW9H2lI4l5EnBEHMndSD7I
FigUi/LjYnn776/akRryWe02cOUITJ2v4rcMtOJ6Gw1FMdMGqcWsnC3t2kUIh0av
Huyu9cboL2j+xsJ789xTb3Y1C1KRJsDFAxuig9rj+DqUmDyX5TS9s+RRSYo90IlD
rN4bbVJM6pKI+W7gL6ihnC1Gdm9PV5iwDt25SvSRYJv3x4MzyqukjWbgunH7K/UZ
wuhxnx6NXT1/eVdiNbzK5YOtsprIBAheowXfVTFZWgki/NsrZqBm2IfDHY6t72zQ
wnUBkNDNnbFoR1LnOot8zGAHkx2cKYfSYyVmRUZDG/4HMGUDRg0NSJODWxWtzW0p
Pb5fw/l4pqYX/XZZTkSzeLMxapX6SElnEEdChzQ5txiB/7mIg8gkRSD0Az0uixhs
A6L+e6RgnZ4G+cVP8HSRRIVqxbhUKYzrmX2I82rnQK4IDLEf0EZccQmlzeQc/2Go
CjVpA9wlKtqJirPHsZM+dSpO/JD6cVBe8Ijd68C+xICPJzXYp+2oRh1gVvfXujln
sLqrQ6fU+Iv9ojR2dWWzKO/QDqPOGvlEuK6d0ljTDS+rDbXEFgJsdwxLVblIcP8L
EcQKXmo/JAbE91YZtTvbWMCbc4rDCVBSHltqRYsTl0szjpLsJ2E3EdSV6J0M/sKl
H5YzQ53itQUGJ+RNuT59497YQRktRvvQaeu34AaVPLEdEwYs+LjbRmsQ4+Lmm6+e
ZxJfiLYtUtbW6moMDjvH8gEpVIRFKuOdHP3Gsx6eoQg1VyhhIuTUK5rtcx90TVsp
M6tH/4wM3yNX2UmmNbfaxuJLyYtcYR36z1uCfl7olZaLrhiUZdgI+8QvN0zTaFkw
41JPQ0ktG7frl6sOmYMPRudWOaCRMF6Hr1lu/mEPVa7vFgSXZx15COCijd/iKWsK
OY93qDhzDV7vFqmRNaJqYf0qvn9qU0vMZqGc+mEj4Etx4m9JcTXR/JUyK/VJ/UE1
3dcbOsxypIxqI80gmvdgcGCmzXokWvPZIgst9mJ7gM+DgdvnboyD+Lut+jpfY3eL
iqUoy/r6kvIICJMd3ov3WKSiY3Jv4Vdg6G36vZAPwbL5i+6AtuwdeTRFWsxj8vQH
5MdD4qe9z0WU5rQ5zq+38ulvaSjaoFftOTl6f3FW8vKX45aCnGcntTJ/n3cwI777
E06rU2AOYaHUsbn4pKTBB3xfVFVSD7egLzdc4dQnZ27YiuNS5+YxuYjEu8Dt6CkC
vNtlKD90uzMe2zwLjtsBDq0C+B/1ZCSBL7L3zB+ihIn9zfwJIucejO2+yDtaVyIe
Btj2c9BwxWj69M/MG4bx81ertafJ4WYU2gvQ/pJZJmllC7Y5RuvWlwBDXo/kmq+P
wAIrRR5GTPPOcprBZMGsN9lNoizV9mHV68xq0dtZXGAZ7oEAlZfiMjm0yFmgbWWm
Hfl3fPf86QSURl6Q8xCekoAbySZzvPpgjpr56jKzr7FKIWqAztv8p8X2kozabAUS
CRtRwz4W2sSv1jy+QMykoPY2BIGoNU8dvRCSjpNxye22Ne49ZNImsy9IV1VqzH1K
xmFFlm2i3CS2KXs8dXrWtbpyarnd7o8JTjkEwSMwq4XgtLzh8fb5P372UJ7+NPUh
pbtjVbj50ZJXVY37nXvgXziTWbPrgaXztqDGEPn3aP32fOOZgTofKq72WgBWnjq4
XrLdSuJWMxCiCtPDpCS9njX9QTHUJSFoeB1gkJps2FsEUyAsAjjPh9hK9h+dLwWr
/oVL+6wubXjkfO9X+A4uzlbKgGHZ33GhbKv5CrqK8OG9azwQZumgzYZy3kmdjXej
tgOGolmNtdiv6cweCQnI5WMsZBORte6zRRhmcQTawMx0+2DzZ/kEGHGv+J27U3o+
3/Z+Q7R9HOwS+hFqORjNJC+XMfTN30PlTfd+K/vlSd1ujYF1VbWMBoprMg1sETRX
L/MYMCNDnEuE0BlVyrs+wwSGRrMBck8iGSDkftYdp5Vubut7dzODuLz2O3gHvSr9
czJodC/8Eh2redXNImHvkFdmu7HTnCQ+CeKxSIrFQOvRpsKG9Y1MIMXPDgLCfORw
b+lqfljP6mUerR9QBIov2POd9lGOq9AKGd0fknangEDPbNXY8YX2wUATUcLuHZIK
p+DQeY/jKhOt3V+164mSOJAAxuO6SgBv1g76h4MAGCibamS75QqY3pXkYMlIOG4r
6AyzCUeFsmzqqr9sKnTC+d1NMR4FRhvBePfRWZSEEArAz3RB949nwxah9uHnjIgS
G0y7hq/ecgs8C+XkYX4QV8zdNTX6JN6xg7Q+opRvRqRKBc+MUA+1eSYNeLpD4qMO
uUluvZDGFGicQZjqIlKNzJCu4gjDtfAEB6r6r/R4In7rbxlWkU3hIq/oOavonO+4
zWUXT1nCK1XDG9wLnZmAyiedOljr9wIlQSOq/kEUQxM+WWotMLVQDtsoTe9o+cTV
nUm8TI8cvU7t/WmGEoxNbox0JmKByAtGDng6pfZXij1rcLy4GsREEE5e7e7qLRx7
n7FKuHdV3BYmFK+NpOnqoT4+JwY+pVGkSnF0JIwljqm9KAJVGoPCYJFrUV46NrzA
gOJ3scpJ0UXKIHSrU1VRJgghCpufgQ7QOwb2quGRX82XmwbaJ1Ky5WZ8WH8QCqsD
PODvZtFox7E0TwY9PPnwBECk1+qCjGcbtYiCp0va6720qN/mVdDwUhEQ4B6i2QEg
3Sk8Y3oYDbK7u3zuSGl1Q/eE4c/gsSNelhw29XlCsbEf2LYYs2P/zM4CJOuf9mD1
eN1lwPUpgnjL7Y1wuw/pxOv/GnF6frozyOpS3iwPK444fJYxUQdial32CA9b8Xab
4T0SlE4vX88C93pRr77yllvL7PogBsaa2etZt7kTw2xkiHVVMVgotX+179AT394d
8nw1nDFhvcwxx5vr6x3q8ACNPx8vZROnpnq9rb1jvu/nL2xTTNFe+9cvXwFOsDjR
3duFSeOjizQIjHQBgG9yKIFmhCyrNbR4BJOJoCc5by+wqTYKtkzrWryBFAx3LWAm
rAmJGVOvGFlgfg/Ss12izQWaoiGj4RDwTgbe4vw3KWgqKbG38Hk/How3v+GJEexV
29mlpZXXLytQG8+TdWwKEBrWuN7sWs/d1LwCotUpcnundIcfwKCLJ1LGPdANGxCV
BZRLXXXsXVaZBsoT7p8n7HiuMCbKWPBmLMXfTRbyFDg/SSdp0j9yryByv6sTQzAm
7BcH3tNF5o+xsFZuv+uB0/Tlajwd1WGrqNmFPFmn7ZRISabyc0KrRkfiH7l3pxje
k8AYWion+h/MLdRT9f5NP/L0yxROnWB7iDe032neyoW2kXeIQfJ0RMEdFHhk0P7/
hhhraiRTn316RhqKa/u4xVhrOeYz3/bA49OuoGkhIdZUHPIvogOmZpoMOwbavkOk
nvFfNwaJZtyFVNTSq9t3ngg58rBWxgdd8RXbJzG7ZrvTAvt7htMsgmVwiW0Ir/z8
o2JIi5N3/QqRO/T3O0/LXbEhQgfYPWDJkcEWExxWU2pe4aFB/IJ5qRG7lk/VlpWZ
m1dVNkmNfufHrnsTqicwlmmX/WAtESmSJ07KvdQX4vQuonyN+RPpfFjYh8CbGc2o
Hg/N5sH6D2prBqODmgl2f33s3ouTUKoIlQA2j2xVtcnolweypMN15OPjnF5TJK5q
thQx4tOPy2wF6Swk6W3pvChttp1Rkz3JJtd/0gF3dJ/Xry51oailUMEyVwu1cq/j
TNzT/4nLtA+qQluW76FncjuwpWf9XYdGGwzTnLG2H9xrjQDgU6+xXP+o6Wl7Tcfi
SbeLnVmbvdLFpyjJDv2uYAMu/qwShFCcGmwhs6frwwRhqozJmM6IhulSm8ZGAbIy
4LX7OCwjsaVJS7Bk1W+hAgV4ORIPnFgQ1gaWZwrrLzt4e64cXLHXIVKx7ra9Dch0
yM3P+21qI3H8MyhuZUAtHuTWvXiKKrK9om5jb8p2O7s8CUxdR17YDXOjN7ZwGXrL
2heeDOT4+hZOCXBWHkuQmRaJUDiEYCLEWzLk8n6M6HXU82OIfBwWewukSVmpISBF
2VcdBWZ2lNSw6azMfiotvPJQOMPKFWurhrkMl8MZWYk/qkxc6mcG87jk/o4g9V/l
OUVm3rPfTAo58xPwYukJDMQ7d/fn6uoR5kkkO2lhR61WbLhNbHnajMGfw+YH5J7i
+Cc+mDNyLbc6SwMauBEJDqEBSdYCNYyfI9Dput3iD5vWaAFEFyA2XllpAMhNpsq2
/sRzJnkglSQzgNIhHiXP7lLzlhxFYv+eAU6MkweTJMp58WczV0/NMZBC8Bby6zwZ
++7vlGPv0t3lRmhaaCnaP/HOlhidafKxrl7FxZlUazvdFwz1E2T0AcVE7c+2IMGS
Tl57elMk+WGC4ONUhHyV3U0H8phoP1WfRCqZm7qPM3PQDNOKOlWd9BsLMy2qDHZd
WilEwVzdmpz5++NmMJ3aBe4LfOeiJMoAnW2mr7YuDh4fzINtaR/M39XlsRMI6L2y
EIFEMAaFS8CbXwzyOoJjq0E3Ae19HmNDgvYGPYQ+9B+pVBm86TtxLZ3WieItUv7w
p+LKj2Bd1hP0y3XAgo2jaWyugvpFke2uEBnVTmlwR+f0PR19B30Fs/NAIvYPW7mv
TnJZ3knaE8bOJYnI7OR+bmFvgNeyLJyQmsAhKmbowauI2GEQrE9y+qwbkQVIQU3n
fSNF50Uqs3rFhT4im1I7NVkKH8FL/Z7I4X/rqpO2A3Y/gFUHUKLGQ1LPJVUUGJsV
L8BC01NTyGQsFZzoDqdfEyF1/INUWla+PL0kHApGHZFmuvkTVHgVgmnYI9WgUyrU
o8KSbUnBPFUx0lLZsUa2gdtYJmGcakEsefgPc3xI14h1JZNazU6qlr3BwzCoEccH
N0GLROX8i+T6pkYlfNiuq2xnJEOa/tzYrUm49ZkOEAczI2Tzq1KYBfErfz1CCUKW
TaKVtdUiYNfe94L1X/T39nCDF17LOTfSo6+O6UJbPSs6uGoTCEkWqpBkj5/BaBik
7OEz+u8ZxbSJvgaGe9e+gKPl/uoOei1eX054sh3kX9+VDWZcpYiPBMUtwiDJy0ab
DCffw9lvA9A5AES5+c1fkyvsJoAjxLscQH4qlPwf7sGVWv+sqc72L06DmJLqFK/D
erYKUM0a9RyS1VgDqDklAOBAEPr5cnOn7pSr3y2DzWgYieLvrPMmSqxRpcHDjrbu
W9LIf16b/Y/DLM9huFVl6EsePiFcu9VKK7kXiPQ/2t5YkXg96uk4WoEu2wZ11gwS
xRQNRA/oPWtWQHQ05EToHnYUVnAvboS8UG91KcY0qLEdOj51sMy7zPnZodl3BZMe
x/rSKkK5Bc4BC0NWcIzVsenkyQTwAbEQq895Idew5SR35TrXQkuxI+hQwdMASqQ/
vEUOIV2XlkLr3POd/35JmzoW+RG7zhaFbywF6IQrxuhtJmaxkApEmjrGQYYiZHvP
PB0/lklYql7eXbxkQXf1PpGzYdX/6eKIq9DZ/jF0HxAeC8bgawIRdU4znarHGQfq
Resq3wN47aqBnFXWR1wkpaY8IwH61M6PtwnsNn5fzxBS0S3Fpq46apTXnUUNRllT
AOF4A/BVWwjwIGgeBZl1KFxDirqgHjRaWR7VQzYuzVgk4MeJ9dhqExk7mUasvR97
yW18V2TBwpJRBiMI2bTjfAf4ou2U+lsG1p0m56KDT0mejKWJoL4OZZ1JbYVu+eGo
bcjrtbP4mN4eMkDPVPKXOLwnofz3UBksZ+aIZdcgaZNo7GVve0sPFD4ZOxfs19Be
UNyibD5IhPwvx/uO9wAqPdL3fhvdXyf8fAzK9RcWBvSPZPNF9OU+kh9Fj1kfjhY+
rIDSZtRe5CuGQArZ8jf35ImoyjizhdtU+bQFFXZRkj4sPKTtTW/bWrCronYj4dok
DsObD5MoDGdwLZzgL9vSx9IZpcOWGZ+w4FghyWzuO7H3KU82YG5wm71DxbjgLAM4
MJydDDcjan2X2/A72aNu9so4GCL3WumAJmESeEBXRm0LVCGbADAyTp0ZvAM5JMxb
Sf7wNTuDVfF+ia+9DqX94QeK5PutLaNoi86up0Zjlcljs+333hg3KxrlwcNOn7U5
L8xfieVL5yg3Gnl9RRkAiQ93mShKdTun4ArtWJlp54D16nB5zfdgk7TmlTLHWd4F
YniimiqvabiRJNk3d+QMZbOQx1uu5CWL/S+D2wyulWnoVAikxp6zh/rrOOu33/RT
Pg+4vPF07AM+J8n6itDW6HMyIP7BrjOfe7B/a/m3+F9lrNlUvljB+oHQfZW6CQuS
1Vc9QxI80pMYSSUD0TKFqcIPPeauEvr5TuLxunc8vWnLPlwA+qTt4bZ5vCJ2nwNi
uJ7tgYqLUWy7phNtDS/4mk+YIojYP06Upt8pFmgHUPvuWmzSMknhQXmG4JncbeJ/
qAjXufhMEbdwFyDKVODVDh42QQ4pxNPTds4qGl/SIIlTIUHKadsvr+sUKTOYAusp
kTCu/F9I+/oSRx0hfqaJMoAmUw4am2EODfRRtcomH8v38fiouVLJ6gfk12QqzzKb
kzCRFo0rVmv59lHMv0XFXec1OVWJafI24TuZ273rDWTAz2ZnlEkF01GQvtYP/Y4S
lqYvkyEYszVNfHoXQ2rymfqPObhBjRSFUrG6ODXUxRun7dfIKv6OyBygJugVT6VS
SGJDGhsTSanF3eZN1L/Tu1i3gt9AbJ98PJ/NcWHRI6ccekE6D9vcorP1OTPj67Jz
d7zgeGzcXhDVLWp1GqyW7blF7uXt3eZlYRAuiSa9anutpKuSTsJiPC1zIEUGBQYk
4dOBv2tKuybGpdx4pROvXe5SV8Q7hDqzHHMKbNkQr1kTuedrIrRd/fRJNJJRwG5U
tC3M2CvGK09iNyyrMBRYgwPJvbAvT9BhQ7IZi1U5TuopTeIRiOckYLSP6Qpb0mOw
qBgBY6wJIdG+BFPEDrp7321671HjvEKuRFDdl/w4bSkpx5RD0fnPuF9xViWCz+hr
h0PamYVCJApHWXXMa/Rmrvahc3J7mRiDyyCaJTV3GNiYTIrma8Ht9fOW3y1+8vJC
b0Yyv5j+tZgpgOwIQFQ/tiLjoAL2p8YD29c/VRe8AhFOgUSDdeY+hx56wkaDDV4a
hSqm6VL4QDD2AV58Wn8/Oiq/zVvth8QuDA73kxUENiI+vsHW+//UJoWjruq9PIzu
vv4w4aMBaepzdSoNbq3YsUfkEQQaGUyqGC+gyPO5PtP+En0Ds3K1NeJQCdMl1zmB
stQHcuHqUyQk6mFkw1QkJaocjY48D6+KhgJzWqD28V3hXO4X3tMqEShLEbolH8kr
zCw5FcYW1HHQQkYCHxrSnLLw34jRfxqZkmiTBBkeAEpdfrphq8Is4VNKRl+99Wzm
WymOn5Bicp1xV/oLVNnSadvGSR8eZdioocNJH7DzxxS5RgKnPypvSWnIJPyoKaC4
uML09+3NSust/LcJBSKyrc4ltXkFIq06LpaY6XIyTE42GaL2kQg5L1Al/bqYADhr
Pesngp/qNvaylFHaO6ptVLhAcQEms+6AZyJUY1eaxarTZIgXMU1MK9MPT4d/9GES
2Zxiu9S4a9uUJFt8R/+LJBmbIyGQ9dRS61TsRABOe2OxTlNAkdOo8ZPoSYBpIlEg
SGHEMQ7Bu14+o8aOmLlnmUGxlRkI5kCSs/GGq5r9A9bRr0uyGxcrB/FkQPHM2lLc
TIUf7W0DgKemnY0jkopreWjDYf84Dzo4tN1xxnsORoPRiSuL+JDUvT9FFxLFVWOu
zjyJt9tQ8M+sHVhLczWaY/n+ozNUcTz73CV/s5XOfki8yvRnkMkGNHKevHOuVapr
MPJd9mNZ7Szsllan5Wl/YeRLQCyUzp/9P9pQCeUo+Zjnzk43VKWt1hDXGh6zIkUn
Bjcvv2VlQbgo6G/AVaw5aM5Yuh/MZNyg/Y0s4Ov+RRl4xSDje0+Ee97rhZF/W4Up
pcmbLNzZFfWjxAk9cDpA1Iy71lkK6sOoBiCDDdGfidUgUTP/e82o8xp4N9AtGOuE
lxiJ9XVBI36QK9H0LBa8OlWALXH0KwCPdobhw6cKdEvPmEu025sXN5HK74bR0LGr
hwG33pJ+lLyq2puvuNOn7zdCuMmFuZcy8ZXcVbwbN5fZmwG6GkQne0/fo5mVsg/e
gxCfl9eF9uWfPGQuuKsXIMPpU4hwWGWlVYORPTC51qrPPNPZFspzRR6Ue2P8m4CB
VsmqsdHFJpvP6rVndTxSA0nQ6tOfMh1IlNJtlroDoDK9IGmv+A6gaL5X5XmKFhxz
EexhkdkRi0vs9RGhZOSp8ktNsHxB/9HIz4fWmR67t/1tIXuWa9J4OX/cHsuEUb4O
wnVWrRzGN3qUTjWQKKtSvqN+XIrLvclms07HFdnTIEzWcMvmY7BNJo+ukb+o5ODP
dpXB4exoTXu2dpzlFi5+ebg5GRm4Oc8eeXdv1JGqpDx11aPKM+4zLTegUuMeaijX
ivn+aH4Y3MwDM0uehVlD7V3GKWudRfYsBSIjj3SrpApVcwQdOX9hal2YsQSLpQGv
9lPDqt/pEEiH8wBXI2NQ0X4yvhO5p4t8gGzz45yMHYQV1sZwQWGBkB/8GPFl6pX8
4MrN2YoKgqV88YjuYDwC62QTRxia2PG0Db2wQaYV492BfS9cw3GvasL1P0IrR/9J
MRaRK8QCd1aR/ll4G+L2XrwGSil3IMzjOtKv9WpCF/xD6K2kkQlck5nsEcbZaBiM
1q6f9kVFbLNJ2sNOr3nJtQiHZ6ueXcKiPueVLQwkA39Qw8YzB6+Er229dyV6kGvU
L5lnTxTM0ty+PK5YZRyq4ZWFG7mUWNsTBlj5gGHOe3luvce0I8u5C9j+Ob5jX5y8
WwuL2WDbO5chjSXRR3aNcawB2q4rjeyuYmCzSnKEJqr+AQhpG9UjRR0qUwtk4Z9m
2vxJxNXRytIv177rsgO+1lGVAsPPcHREk1qAKmjsGp4KdnobePn6wr9sWNB9gcL8
lQLd6SrkiYMf7e029/BOeHy/vPve6CUYQGZtRxjBU3mB9+tgxDDqnLgW2F8KROlu
pjzTa2xpFZRzq3XluBP+oTS6J/8SAgCZM2UngAdaUUbTXCR0o8YnG95GQTcK+0ng
yrssJ5Ry0g48W9KDsp/hGdnnsmyjTCK9PfM051x7r59WaX+YnOF3WCO2CrAwmDdM
STPUdj/3x2XQWpkF9v6erncg0+tLA9KWCIokw5Uhy8VnpIFjZrolDThLxtUu9HBT
sxwjViq6zUVK7oQ98K1St/UYuMdAOCRgmQ/RLzhMp/1R/Zlnfe7fviWC0xW07CGX
IHCo7GGVx03oZBPEDsfxBuri2iJd9eulOU+YZGg6KiBod9hhqXp2rYeJmds7gGRW
GHr/xC0UiVHfceTomLtnkLdiTCjBJtdJMjVgl1QRiAG6SVW6SdaQjdY4Ph1xa5Uc
ym0RSpK/hnM5EBxwVEpnfSfDKoaie+zMQ/+Ud11vBE36TBymsasLgpJBcZ6uQLBW
VMe6N4TOrBXyenmpBgmL8SPVx+vNr++5g0yri3bujCjFaLRaNgS7Ep7xNrO50oOE
yYCoHejXK20AS5ARHwfruPpaqF0R/m7ST2nBvS8G53E+lAi5/hIn2XrK36WnJujB
fNqs0mI+4ZO/ilDx9lqWfy0EZaRgbNpUKPfMIEbeIJ4LIh98DPvUwcvJH6RlVtKL
tqIC9pDYXr8QP398Y/LcaNJQHI0K5br2F0LSot+ssj/3dqvaY+45/OPxGotw/mLD
FBm/vJKIvdty5eTbbmBaXiICvnVt2eznyBHZSwxhrbHL6x6k+abJUFaUTRBH17pQ
IeCnidSGbY19GbhadmNH5lpeU7FBTmMMlDgBE1Pwhz1J529S/V/h/SQ/BjiDAmst
mVMMN1IpOynPV60lphjipJiFU7lb20yRmQTBmB1fzJEHPIkxa0C9Xdvb/b09cGHq
mXZcVXPdC1t0BWSvpv6zD1leSjuG1KUTsyp2LAh4Z5gTWR9HGqpMfYMPah6Ll10Q
Oz6JTL2WxW+BF73hEL/CtEFNoqVDONSUeDgxletheMFgjNsHNx66BDKhv9zNonDi
gO5qo1E8ANAIgfFqSdm/hZaVmN6ZwPNIPf6lxowOaQHVww85bAQFjBVGQ+4Rwp1g
Zu8xzrTxgJPl4eAD6cd7w1Fo+oGtuO1C1K0TH+pMSTDXulf2GzvWuvvHmCC6yO80
zedVPjMwz2oJWYeFqfAn4ORIfS6IVfxkt5n+NgdqW7wEaB4EBSm5ahQnwdhh0xim
nDIDTn2TaBTJ+N5iHAf6Td1BNP5SfYz7vZ4PBVCfnX2+hg0AbZraqt7i4Z8h+v5j
01ShQzxyg7s2bLof9xh/zvqcNhamBDc3mzd1EKOPsWsY08iNKGMgnnQj++Mv3rNZ
NBYui9u6vSMsUk0cQBVc3i9fcdIhtO2UtpIWpcvi1l1CXVkeYuahm6FiU/Ky/IXF
zqx5mtauf+daMHGNQ0OflDBvo3+4cic1L79ImWaj15gFwBamgBTnbQvB6D9BZ01J
AvyglOAfzHA6PM4Z6tI1Xy0kZAr9J5uteHTH7vyqKSv4J5g9SKhikkaQouaypj2A
asuXhzTL3ujVao4DAfzgR5/+Je4oLh7CGdk629NM90cFSu84Qx7XiwKKhnBdq1Ht
9+qi05wHX8enf3uliMcKiMK2qALB7cL3peD5q3wqiwuyzg5pvIWj44Py161WmO9K
qip4TWThvpoTGYgjSCnUJRLvPk+S0al45/AunxJOg6VXB2roC0G7qz8skxr4jN6l
0IcuFrTXwUu4Wnvb/DiPDbEnsbw1m7gRt8VjlgjVjE6E2FjC6B1wbh3dIdGbJPRU
6aEgW/VXDzWp5ZyYvgxfEEurpPEocnj5nakw0S4KIExibJP+rY2Au2PI/Ng1Tz0M
1QY4d1g+QYXHV9VmxcbuQaDdH434CiaIDfRUqqi2r06FGgPSVDJuV3FTXH0y6bE6
sWmO1C1+hhADbipdKbQn0jsy0WhNWbLJhraPszGHpldfDjha+Cbt5SQ4CbwmtkfK
dTM2g7zeQvrPtGZ7S6NfdcPpTm9dPFNSvY04AFWAobG+gLVR3TujUMOCCLDPfXwU
sp1yODI5PTbwJNsJ/pzPSgPT8OpyhAsc1lLTc1cF1q73WIXj++zF2vXu23YcQ/OQ
EOIw0RhlZpcfazJf2suYud8pVBh1w9eX9+8C0ohizUb9RxOzsWBn/VOQWhBVRkEx
pLYDH/reuueraS9BfhVTXIb0VWoxtpOqOC90Wc3xXb9reeBuu22+2xEs3qMJ5SRe
zdvb/zvieqcWhbYXWAF9OGhGl5j6BqcYEDOCzwMczoSnkw7xSbX70WB8ohjqd1PC
u6ktbaRULinefzovwEX1vC1AvoqTSe78NBDjBp6mfdaFCv1AKUCw/n3Pj2ro9B5S
SbEnHrrQGTwrBKOWDIA7yq475ZP+shAMbAAfgjR/tM6QLZDB6LwlF20BpStnqldY
wfNJmGtgQvFb1FWakKK+MPORJrOdcvPjWXz0RewarTLiG8yzuPimGQ5biqwDpQTU
PBmoAzjNjVwuQ0ED/rQNIZxTWgbGdlpW93NCCZnpS6tthuRFebM+9Aajr+qJIIGA
rAUPqj4fxA280oC/nfE/UYztEXPFpAOXi5T/MR4037LEHykbMrk0viROi0T7q74y
+XT/tvXHO0EG0sgO4ac0JHKAjpwHNT07NHhNUiKLsZMTgsKSYY8GJL20LFyZl+jC
7ybJcxgbrQUcPMStniJd8bh5gcS68BDlAFpb7GUt+1SCqb9cD4OH2FHAsOWQ10w6
uhwGEZfD1tCEfnLIiCaUVt98PcAhJUtKy1CkBP5Qlf7F3Icm/EA9nM19iEEtgX2b
IHaPSr22mCE/URg5JXLdrKR8SaslJtkvedqne7IC5Pcco9pNN87F1Dqf4vmGKNRg
3BKAf/B+8ivX111GJVDqi/8bjT+fMYG8kRvgeBwxw1sL0/VYI4x2xI5pqpMKIHRo
ze93EP3sMJenFai+/KWZBf87/xL3NkNlAVQA4SrgfmhdLZw0eiiBmobNrL4W9i/D
6s6FjhEPUKmdKVfZEGuOJsssmGnRbczk2NUfO6B6H2t/7SdkW8d+tTrRPAe1O9uw
LhnKZePWp8u4aJY7Gw6MvvjmNN39TIYV/M7ZQIY1Yvb98I6rKtY5AMaqufsDstgO
sV/Cf+dFOCGQuDabbhcKl/qHuBJtREv4RaRQdFecz9QtNCYvf3LcpoE5paPcIVEl
eET1lcfXg+eUig0Eww245R/AutByJnDZy3M4osKbgUHYEVbil2xsolmr7KdCrZ64
XgpPWFXrU271f11QtG66/iu+0DejRdbAnSooqRM91tQrZIcPPR1FvMe4Bp0FM4sv
iQNXzCHbl/kGRMqr25949AYBbMW1N4Z2mOM66HWunTsVgQ8M9d1PZVkmP7ZhYCts
hiR32RjiUFUUcK6PCZGNBBHgiCj3n7ijxOnkSGuO8v8b/1gfsjSsTp0daF4CqqAm
JyYZKxuwtcc5ysFlrjnhLsXt79WPCbaco0dNOxj6WBQ+oQqWeVWgBty0+pg4L5KT
ODZIenSZegPVpPVOOv2BDgJ26dXR2lrXAsjPI8yBs3kZihRcJfeZQ4TPAAUKyg0u
D2htUzPmon9dt1bZxH86kQ/Z1bKJkcruLvwGrKKLUMNJQMGbJ04MNJO5/FOlTiAx
WzB4T7/nqAcZrWlYB4BlAYblsF0c0zVS87Ew0LnX2IMddGcvOdsXpFVS44R49h7Y
Jo57qEzVoBIOX+U2Eqn01Vfuxd/t2KDwDpdYcPE3bjZngUmNbB2ZHtyT2Y4J8ay5
w0k6op5icfCuJw95rhJAyP9ioW761ybabcQ590g1EXqGHURceE1E5P+do3RejF9E
i0tOFDmc5gIngo/cZlqbUIx4SZt6/T+ONr/fomW7I11SDwUZxJhUB2djyQ0ZVcm2
5IIZA7dyL/06ysV1ZVYTSzS++1C7HkV2pZ+VUG061qths7KKes4lPQPQY1nl0CDx
m0+d7wCKLkkV+ernmfsAByx2Wqz2kMd8LtRQGzC1RgHFglYO7w0XQYs3Bnx4mYMj
7jM6/sfcNX22ILPPkqZHV4AUT6czq4s8J+VusLqpgF91dM1U37+KfT7r7zbJkorc
+5VJUtbQNhJVZdI91ZEtRQoGkbTF0CS/ZOa5zpi6wwAZu1k4YzwI38J5344Vh+mn
oGSvJdCcB+9qvsX8AXdeWnCMKAE4aqJFrA9g0iF8FY80SY4aDTVDPxElxDp3dyo2
rz1B6trrR4ftpeQ2R1JLHFCbDhAZRU5oGVYEBoPq8e20TFTCYsdPI+sUO5HxTJxe
yMcq23ObGCkngwSeCMIS7cvpomsyTrbj8VvDS+mVqrGTq8bA2qb5++BG8D4Lx60c
RkSbp44rKr5mtqeX3s27yk8H4jiEABtHH/SnlcvGyGlXs+RYHAg4wHIeFRM9K3rR
WIpRrfzpwoQOeaBsiZv4OROOgLBNK3ijapwFCYWBGbp7rzOp/B1EQbLYcwoX3M68
8Y38IeG0mZyO30CyV+PiW03Xi0EhnvGtBlVZogYrv9YDY573N6Je3RbYIco359DV
uJj6Bn8EIOjJ5tNdBzBym3NhgwGverE5mUvsSgFSjqFdUEzQBFbWLoUY3JN6YLIb
ha7/c91IvPFZMMRmFNSKT8LEdIN3gy0YCuO+HrO9R+E2KJcQPl7nJw5Y1ggBrS8H
m7hkb8nayAHc+qubLLNcpeg4v1qUvEobj6UO1SZ9vCtaw8xvSIq28cDyaLYCya7/
tsPnbbkIny0O5JtIYt2vvR8CM1kCiBgd/NNhbBfQyZCxBx2xvi/N+OCyu7oBTgEV
XDOn9czxLrn+hoY1HdcMWFNgabYyssBBLWMxCyiFZ0Lty6WGGCrLFcU6JtZOWQvF
Qv8cww7ET8mPIj2vXHnE9ukA6gMHIHRtBG3wTF0aBprC/oUFVmW+BwHvIV7RSaPn
FNp9OjfKgoC0J1JoT0TqYeZVKjI5bKO5h7l6RxwCxAIHv5tPrAWboGitPmGPD5oF
mAoN/uWQbDu7htn7WZ7CzxlENGgnQVOJEQh2CuR90ujOzwrpdCH9Dts9MBXXoDbD
zdxFmdVL/0LTykFqOb8cygG3O02E8IV4cw3pcrDbQuiDzEm1Mq6WJ9EsBqLqXXjP
GfC7r/YlY4aDVuSRyW1Uy6qM5ck39uLyvWBYGJ8+UYy6LD3eKdz/sgbsRfkGzUNZ
RQ8a34gIwgHgCYApl11ekCBGQvGKNyFB6eUOW4HH0OMqOyjRSA+bHqS+oU1ael1U
3N0Cqa7jk1jw1KVoc8j08/urKUy5HY2EnPo2NnUJRlWnm5c2XPWvLPvnogxS58TG
1aIAe2b9A8HO5mKw38Rk/hvoTJszz4gsIxGcIOgU83OsQj6LabOcTydCvCAwCjRi
oxPFq/wGzv6aqg/f2Y3CdBOXv4qGwWZIjOqQVKgLi0yNKxbD+t5l8uBOe5ARsPp2
OadWzLb6JPweRqDTnjt8ayTQrIc0ABeN5k9iskWP6o5pQdK36+SVG1jQtrE9mXwA
VwB6O/mAXhCzNOURchobDZywgqeULS38x8JKNdEMIlksjMB1TXB6F/wHV00bPTgK
xXwxl76i3S+Nk7VZWCfqUb0UAfIALx9PykjSSMULdA0Ox8IuMzpCP8SWT6COnP1y
ZfjLUdKX9h01iFz6N6XjyBX5qQbO8s4LSxttloq8pjPoJZQEeThqWhhLiFSm8da6
7XEqmZ5i8vTRknuOWI2vdS2wqVwRr0Df7tikaTxN4MbKmIbO86BOX80ShRdWu0En
rORxbyTHwP/KoKPtVJJlrNJjmaU+lg0RmoCkZyRt7zjrhsbTokXjOTfE6owdWqpA
JGZxqRPnZ9Xlx5a6eQuGXOcXpb5Jt96gwxh6lgUrQ2x0RuR/M4QG3jsuQ5zLKp/f
ToBqdoj2cA0mTrdV3k9KHjaE37F5/xnfM4vRDiAZS3Y+hv6woQ6DNLQSTp9fBP9e
t80AhNKCOLVSV/4u+MDH4ETklzKkI1oygXttOLQNnaqKexLvUqn1Sn+oSwra1xOG
I8ASB0jbENiSHJ89YPMQ/tqUnUy9DjOvRQAbdam2njGojm3nboilGeuNhmovVT7M
sW0hf4UXzoydrTxv6ZXyJwQLS/YenYcH1dP31ySfCtCinkKt10DrYp0VhHKXcyrL
KwDrG+DuP9/Nn1yI1s25Rpjr1P0g3e0ZKDbbmd4dTJg/rZW1cR3CtRLluGHMsBtu
ox90KLpNQCA2r0Ejdtv8mJskdL5yeGZPBwBekCHEvhGKcL3tUy39sSRQG9alwpVu
F7NQ/FYIsgj8XyIxqZqHSIjnwSFqvjGdQOkz2qSWSCY9+yW+X7b7QZMldZCiJwvR
EV1NXXgIAc41fYVasYg4GgoOph7IvAt+d+j5iUtd8nePAOVGQ2kddqPs0JguuAu/
weEiIVC75cCMEHk+vYaDetx5YAZRfKFiRYomsdQ8CtDtUra5V58XxuLtElwiF3zm
WPJzGaAmxTsynbxKh079pEGpbd1/38U8W1R7KKrvJ4kqG12oyTsIfGo3nCIH9JUs
2g2DpMSJ2GVu1S+l2F+cYYl41XZp7ftgxEssvnSXvsfQnqKcbVx+M7KJqEj5/9I/
pbY396uXcdBjYLlvXjCWyTRWurnzejJBipnCik6/V8n1h70Fk2bWN1Ygp67BKgJ5
gDolFE8x3qHTjkABo2Ly+JNr0E/HgXIxQ9AOiTALUPglui6bDuxp6TAdzNnfYD9j
9uU8zC2M/ZSRmmjXfcpW0zUzBkrKHEkLcZAME1jFikkHSEr+rtDqbRWZGRdZpfoX
SqgmpLHgooLxKoM1e2t36x6dPgbwZXkDvoJ4wjzehNmzD9IcUR6kWI2Mbq2HbqUc
/oM6yo8qdljro7evaAUw92RDz+7iei5qadmGkeyMZoRb5JBWqKjiGsP/AjH8cevX
/PqYqO2VF07kVpYM3WQxXufm+UuVwNAPtK1QCUvYWghSrmRJ3WkuCQ+VtQMt8pt2
wflu3sj9Lbc8Iv4or2BAQqFaj9/M8asVNLl0tGw92uR2yUmj9X1oKR58ppH8eqrr
cFU/ew3IiXbH9NUSfS81ea2xsoBEr89CQJCPa/AnxfsmQR/LE6Ij/DcLdRNRnh8r
/c6030WIQ8dxyWU2Os+eu5ceABuohzWWMHj+vARWY8wBtrmjBNxA6Le73bUckSQL
f5ddDxQktSYSEGUauBDKEtdIzgMHZBDtgWGry4VkR8cxrRCJS0/qEJBTgeMfriz8
1m1eRMDLCQMngzIJe+TzU3MAu8/bJ1SKG9ADZaf0NmCIzrLgzK5F068/ppbJaCM7
a1oJaniuG5QgkTJb7M7JFBkwtEg2pVNf0nIdqZqyumMo+ZVW3RMlwKP1bLq84QV+
bNMkTqJKOUB9kVkE8i1XQQtDMbGj0WMspfgxmtPbl4Pcoa1Bj+vZsB3//BGjeS/l
E3/wRbaJeJp4qNtCeBPUqZYbasqdQOpwE/WHc8+hhuozmiIkvZtaIV+nIDgnm2N6
bC4eLwpJzRgo7/PyruOcNVS8RclTGTEyhmh+YC6FrQHUpxQ7wI7EChYFrr7Mv3qp
LxzknDNZ6PWotFny1RBo++20QT+CPNt0VF0eem8F+ZYvDNtB7MfAQgff5yvZCnzw
FPR02vCcW4+F/vwBs9UnHmEgJ9iGWiDbxMM+kfCRyHLU51jol6dvVo7O+2aJMlH0
vI8ZopPrub7Ac83h39H1+H9Ib8rTJ5lolUi0UvJUNlEfFNfsfZE1xwaKmxRpknoL
r27i+nCiAgy71lFgDX84+Xwjw18ukmsLETJRXScdw2nLX69DTUhcCcQkVGnTgWYF
eWUFp8RtpuubTn7sv17I1UsGRCUdgpizZib43elEuuXLdpLjOco3iwTAl+8sTDGP
jwWfE7uXFyYPSjach6Spr22vEUeJEDUBFXSXgACvSV9UrpEhHw4HwTIKO+/4WK6O
QO8iSfg310zpvCKJS8/SG10WeQPfcwBfwgoHE1OD0djqx8eE1EC5H+xNZjOXfRpP
dgH41wK2xnTXZjEVjEswGAXb2MznHI7r8XSrP/OPzzPgTsXEeXuEa1B3rJHp3b9d
F7id93hM5Z5qQUoAVN7oQvoaCG9sENSTzpJG9QHFV1MTrmRzSRL4MCRE12mWFEJj
95ILPA93L0tDO5svCZGj//gJbkUljGFqzKPFcgiNLYtP1Up4LpXAD/FE1Q1G1ovG
XQxjTbukWDYqFbDWRm9xrf7byIlVf6fjBehDemxgdC25YRbNhiHAOb8+O9CwTnbP
FunwBoypu7Ng+x2sE2mZBrLaK8WFApTKzusKeyAmgIOGuc5Nx7qWpwD1GEDRanKy
2cfqv2S3M3jaPDdGTkT2Qcbvwke5owTlUXIoZo8Pony3gm2+J6HZgwxAKq7Z+rvp
BlX+ELcNy1PGUWVJ4JzLRGurRya83BUAm0yr2i8+6p78/EtrvDLIv4uvuAI8DUY5
JTwCj31A23UJ1+ppwObTGEJX6kmCpz0ez9Np8SPHVIHChDHhjOxDW8g/JJ85QNEI
m6CA+eK6d4XCBJjjzxryHX9vh438qkv6IT0Cvr3A1n0F8t9GMsqHhxX/n3+a6dXI
hDfieuft0HuOKI4ehgZqxfQAFL0wU1GKnkshRTebkWarZSXIi1pS8NkG+dj9enGn
Z5vqSjoV2/n78rog32fRlW4aA7jg1lJ1u1BxGQYxCaEdoAexnZC+rKWQ4oirIsBH
KDD/MSTth/TPsOPhRx+7pRACymkd3Dm/8qBvvtz0tDNE9uU1xIRaJnB8bSiEKFMg
vsYK9ArB1o9v2vcgtRiR71YO77seqNs8pnq5kPxcv5vAV43Cfo3ekyNHLBKegJMr
Q7u0U4Vb9c2pAPmaYBFj2OgBz6/KGYWVDBzHH8MXMw8ImvoozkVOshCDQIshFc+s
GGYiTICPIteUAGhbNrrwISqTjZicFEnjN6s3yv3wJ4hwP7Lkhmnk64fM/J02435V
j0AvSt8IgYtm6IJdoi7MjHEmXv0aSQmfq6BpOqIfNQp69DTQBZB4JKt7+GqqPy/n
Ml4hc5GUNpyNeVCvHCaIq1bpQzcKXOd7lDH5go6+H7eq/tg6MftOCSsa6xLlywC+
F82p8iqtKILpNOwSBXxv8gxRSx+nhLRTwbuaW3VBpjA07GJ4OErVNcFCNrg3KHcu
5km6zD4/zowNenGSgfA7d/1y6ZnNbE0SERAiZcopcpFZu+iJnH+U3N9NBaD9cYZT
QdIG01WvtUmVYmMU7tEZvHppIIcfM7qWAk3/hKAjHdZ8xcALRKJSA2kIANSnv4xU
COz778hSaFQr4DQEP5K8OcOWjY3wIJO7PAm0z54pBE78qc+t+EZH/ru5f0Ti8IoX
tj5D3k5EJ+2QbL/KMMLcHLG+LBymHinttVOpEGUDrXyS0qppDDWAV0AXQPlqdbKm
1N/Fx9yPtvAJbXsbBw8BZ+iWBdHzpbG/aCoNBepAWKpT6GlpqZZZRrNSCpQF+F0V
HKoW6yelS8UcK++6wyiZHKV3wRH/VJqQ4QSUYOVf6qcW0kK9o3wYnjygtPfndlkL
KI0CgZ651niE1ViddHfOrfl1W91JOCbucGCDYOKuYGIp19fq8K6MxGhN+aiaaY8j
OTsSwlDYj7AUznBAQk+EAq5KenOYGhILtNXH2AXX+THsa2U+kdsBLaID++iMT3tg
cFUqDizrZ1Rd9ujFFHh+r7R/A55aOC9o/e6Lp9xHG8RSMtWmP4ztRyfX5SDcrhxQ
JiC6WXvOTKFyHPWI2F/FZ7/rVGaPdlgoJLMTDGtB/rc/JitN7W22nawUjHh7pvIW
Id+HormFeI+4154jl3yoXPyX/XYdezld/zO1aq3YKkjK35ujVFsLy5mZaZOnGYKU
bTBow1oW4ED9B2JpmE5gRO0+0sr12eP4uUVUbYbnecRnNBfDe2ucBWAJmD5BrrEq
J5e92Ls5ZeTGd/mH/w3KrQ7U4bT5ucpTgs3e2W8dFzixi/Mgot9vEvkHpTi+mLzj
aie1Yrv5wkE1UOROO6hRij78XYIZLpxLV4G+Z+1C0mTZGxfPD4Uy6aPVhVttrLnA
96laLY5VaLjzXho3CF89rbsVIM0dSIsWQ3q/+iYoJoSMWAqq2rdoKVWWPRPbYkmU
R7Jpo+RVfpoYBwvQ+6tHZJ334eoCygvqFkPSK4lqNlmuiqdGWbPrWLLPH0sLLPL4
y6K/t6zcSJKMqet9oK1+Sra0EwsIeZHrrg00xiNtF1lWHOl79FMVSLy0C1yYJmzi
NHVymKjva4Pscl77C2HMJxs5uwz3xY3xGevuFxpAWdpZq7+nDMNDomKYeGloHYZT
fY8ba1Wi9CNd5fWiO/8907wC6m8AN3xZXrZsFwojmmej2b3Y935enXG+gd1DpZnj
GMRL4u7Enf8Ou4mYunuXlyVxlck9idTalG4JPGIm+rTJsZ7tAAnsVlpGVVF6tCan
JuD/SMu8U/0gQ54M8mnItVijUKcxigeLGTzRw2kjJXFx4aX8j5dcMK9MJ+U4Qk8q
JnPrIjl6tbJjfPzHxPZ0H9I2sS66vJPd9Ys2gEM7erDnFN8aqCZwan8GgLaafdAO
/TeKUvi9FWPAsZZW6b6xzVGbHPVXMZFHz9YO2KJ/QwhZr+8f3f+l9c6RwH6dkwYc
gbG9EGbtYtzlP117C7YboUJ0oLVFkr61pxFkwtrHQfAceRh/0RrB86vQMYjY5WWi
0j7sZiJoXoq5nyKL64R8OvVWGdPF7K/sFZN/NH13ADB2T0j6IsD1kC+vkl0TaOP2
ti9uVSSBs1YiRpJMXUqnp1FP1BGsJ2qh60MbwewiLx7Ohqy47lNu9DLqetqNshR1
h63g7siSzX0w7y45lUizGXviugn5GnIdS9lrfrX7TWAmXWwFZyaexSIWxVI/ZWLa
5oLgOr65ZKWPTkF6Epx1W5hMwsbV2lL/oPf59LrEbO85eomxaGHx4y9R0X/HT7N6
9w/K1O2NUozHqAFc5/FM+h7lt4w73zMuo96jeSFNyvXiHKJVW0y8dqYvjhR8mPHM
pGY/jW9L2smPPf/gmIoSK3BEBkCflwO+f/8XXofuXSoZjSQDPLseIyXl9xfaZIVN
Hud09Y0paBVVO8EtOZT7b5nzGjBk120Rh3/LmMtMs9mWGExK5PMb3xFlccwgxI2x
0kPDMS113ayrf8trHMLlwpnZM+nkswcvoj5mUr3I3WOep4J+4YoUEZgb9AjrkBiq
+0naCNdA8AoZWJH1RH+UtmQtPZ96UNmt/pe9oYXERh3KZKHVd6SV1UicnpgI9MEE
0rsSAgou+l/9kfg+V3b7RQN80e6o+msv42/QVg1uqOKgxOZJAzEQCGOAN8WBXlWP
OwBGUxJ5Dn8Byl55sYCqfAW+NFWeImnZXtCy1x1/eG8kxvMQXYG2IUM7eGH7GpsG
Eg8IKabvwEzH2RFUkg0WWy47ijs9BRZTuvk4zXmPybQGmSTewMCH1A2G6YUyvaKg
etTocIa/gVE9TlWYQOXQu6jTsot6O2zQk3pZhOcHNDQrC5J3ZY3i83FujBRpVze6
3eBAupRTXDbFyT98fPTt9J6YWcfeIZ3Ti6jxZ6CchIju4cEEBmWrL70OI2+k+KRh
b2uouSokiHNfWxxd55LGGyH7rIrpEyoEeCw3TOjsgazrGFn/tJ97A1lJOrWGeY6P
sDTvmgdRT8FAq1yOE6g82+cgBzviFNvl9iB5Cvt4XGxphVEMpqLWWMp5Vw481gDy
ZQvE/a64P+iSgOBlPy6K1fgDKuAsyU0+j0my9iZRvMu1SdsinbG+IO0E5bT7MciZ
RnJgdI9YvarOmuXrOP2RUxQ1zrw13ROoKx75HAfrpIk6FU1mfvEL8LVSvBdeTLfT
bG2xnuzx8k37yE/erL4vCES1wyQL5YJVFpbMZHjZ4D8J8Vx2fPwZKCL43GyAiE0U
kBaEBzNRyhk5lWNas2+8JW/RN7Kn5hD1UphfDOcjPEg+om1cOQS5WmMzrDGYI01Z
bFT9JSNWTs4Ya+SdRippO6wq4ioqFyqPWyXITxdeRw49ZfNjK3b2grPh8S0Xd3GF
FWjXc37XY1IWx3la2oNKxAW62VytCoiEPXlHn2MGJbqd9g63Z6bP1+GKtcBy7hM0
5HIDc6e1VkfAQ4KXW9x+3EjKQMvr220SbuvnG/IKy0HVNex8XhUykUbODteNgvO5
ycAF0u2mgDke1+X+G7oaHzNrcjSLnfmWcWSDo4TqmV6V1IrHjkLJdZEOJ2RIPUl6
/Gbw765owXDwKTjlPVWI/qEdXm6TTYxuubc3TH7EYJmuU9S8ht5kUwiHVwxsYGXF
m6/H+moMCv3mz5oEVeHBVSGabdxOMNYIK/a1d4yrqvHP8pB5lEAFZjVJBafG9J9H
Jbjs5MOGdkkz1RrLQjYJlGPBkZp4AsBfcyNU/cUwXjpXAm9yTOzKablmNJXRvMbA
J6J5fKClRL3DGfct+a3l6ZYwKRpMClXbZMptpo5QW/5LOK5eUQ1mxarkS2uJghuD
NWXgbLFfqNvGMKjDvNa+z8nt3nqfBolrcYeEPOOwbwvI0zBTHFrw0pIAORzsC76s
GfW13lAlWYVOc4/Fb67r0I9V2tRNDaTKwAdUxUwASkYUSuCFPyZ8+vV8pl9KRG3c
2bM7zhfwsuOtdett+IX9o82Ju8/aY2S/MNMy4sYKR4J5qr9EVNUKM4H1GAie0naD
m8V1T6hE3WtaU3Rq+lCiZsBcm1ESjaFymND31lLjCtKAKqbQUh9btxXIGFxuSfmI
BF5DrzdjlTL4t1fzCjApscQ5x5fX1WvWbn8Qdel/WCvGzTdTl56Vg6NLEcXgV1kG
0LukptH/5tzw/CBMTwc6CXLQzHWeTDNe4FlFhuDpfknxgdBP0/wi9sxzfSt7y4Jh
fElXsSr4hUntZ0Va0eYcxGs3gTO77PDqv22s5oUguKsEj9UUwp/hkAcvBgK1V0KW
zhuKQQqa7ZLOXMObsP5mEtAD3FPM2i+Fe4m9SdLWjkXZxoGUs1bOevK//rv/Zehk
z8MnrMO/BoDZNYDcw0m/QTBcz+BoG5++6HWsOKEg+y5JCxe8x5MltoMAuB4XYcVM
tCTQea+LM7HHiO0GZ+HjPghtoJeqG+hQmUhNY6E8bFfZWAEmmYBJaacCh53pMIwE
BjmCzJgBpAupnDh/RWlrUECg975Bo7d7W6r30p5BU4k9LErX/G/a+3QuMhl4SX6h
JDhvDxQidXIjvyYAzyHIYgCrUKy0rLljbJLT95i09J5fMPs/rY0p/zbY0+Z2EDIM
zOJe6rvNjmPrIs/cNl9CqP2pE2M3ffUjkq6/yRF2zp0nR88AW0LPINH0WSyQzkjL
VGFaZ09ooL4nynwhOKEAGgmayEXANzRLc7SVEd51yDYFwnezRetvSpBWYx5TRI7d
kIGtzFWrGheiLsCB7ZDOeb6VM9o7Gh8Ngc0e1CdNMVHYgAWLtpqTwkNMzFlEvolM
NYSNok21SkKuHWj27W8klVBZCAURtrIh5AqYLhj3rCQGISRwx/tPchfgOJcjPwdg
dKeBHcdRzpEuWguBo3pcfsUq9/hFhZ8P7mYYqyiTcKbhbloXpZWinwhUNqcY9VtZ
0BMbr6NxiRtoQy0U4MK2MjKCISruh7/eOm1R5N6Mo6Da+0ZrbIj5KMy64hN5R94S
tCOL66ob7jepdQwJprvTc95pyV/X80MyUr9f1ox1A/DYjBeFbmaa6Zv5AprA7J4k
2lcN7pSB2QnZ9fnhLOBuiDmsGP/S+HLDull0jrg3+I+Zt2nEXeC55P7hY+TBp5j0
Ley0B0TJHHrMVQI8CYzGzBHGUDcv7d8rN5gAxsxbrQe+e36m5XiIwYKZFHcozH9Z
cCYpSleJ0w7t8SF8aZifgQs4ycYfAKQN5SCrQK8anZ9GIOuiU0IrbM2Quh/k/e96
CDRcx+nJl9WHtrkZnPMjRfYsudkbVtT1n1w9TB6OTjqYV7FKI+UWXSWeRbRzL7zu
f/jfJCeHDCklpR/pIIP5hZm2lO6ssk4L2pA9jMlQelcUGP6MDMo/IFmlcSKTMasw
roh+DYBBx2bnwdfHM0p27RTKq3gYMqdnBtgXuHmVajAyio/6dqZ50IF8uBG91VVF
9K4tJM1xRmZ4bEYPYqJmNBB6oBU4jM+9umN2eg2hNI0xZlIsxVoDiLnRB09V9/Pi
rYZCWv5LIqEqTKkM3Js/sq1IfpWYwoInDxsqDLkzRx/jlNOAXj9fPKGgwQaTY9gJ
RNm11WYLTVjyng0qAzfS8RvUIfrGtrCXzxoVyK4gwQduSKnnLuAO0IuyZANrYvpi
RHVRWQYsASli/gTnajazz4DZ/6wsy0fPH2wsXHeGhFZWuf98A6rU0n3jIy+gdoSu
AVmZzSoFFgSQ17BiTRlrOXJmAn4vZ9epeZ+m1zwlmzLLlbQiMSSOCqJcPv7w5t5l
3dYPt3reFhPO+sZRqPaZIPC8eP2KZzRJV3wCid5P2avs/1OvhtFcPHwPsOKiAzow
kjqaP6vZNxUEuCzfOeMDyvLAV4BHGJBtuJ5JCinWYD1vLStRMVDMtboGqpuRIBmo
fekg8zq3IILDKPiEOfdZ048rk4Y2PBfXasTcUXkTvQRQhMgeWalpEpXAnfuqyK+A
bUV52OZny6T1PZeEtyDJjc7lGuE64MASNKXn2mQTjiwU74QyEVZ+IQT9r/H4HuO2
xHNAnV8Hxx9i7g2W0F/7xEcKshWCRDhIviHqRvnp4fqe+K0gERdfP44INTiIJhKQ
/cQAsM4C39hHM2EyXR4dc97mOm7f0okUyMJXlPZqk7LIkcccNPDJmU3ihCN73QFR
EhUHShfZwtlEnwixkbsfiq5POEaclCufjP0+2rPU6e68DdvMWL5YupYqcLd5k3yz
ENc6Grme1/smG2Q43q4wm/s49/S+XAPKtE4Bhu6OO8N0AaD12n9oHr5UY630sATX
hzc7jkWXyswMiWa90o0Iu7m1cexEEn5feYqEb0WMVQrRLuYpBxW1OLK99P5uwSFS
E3CT/C+0ySh31pgSMDqEu03dUD8jI9ZEeIXlFhiplZKnkfV59hxrFQ9PSxU4PvH+
R2EgxdTjBpntsX9dgEINpGJACLjf7vmKzyUWxvj4wP6baddWPJmaZ0PugaBhU5UI
yZFpcvchOsonWhxNEPz/HMfeF4LJ9ih5gF4xXdb8nmDwo8C/mHgIaO77BSzjN0pZ
H783cCLkY41Gvs4A8dPAJb+auTzE3HYdRmJdKcfsZiv6D7Zd6nIEibXzYWfCA3Tl
fR3M2nvquCLP/+2l0Dij9j2QfERii5wAV8meO4fNjc3g4gLqQg8WS2b+1u3e/Z04
/2PSMfWyjaqyW5mZQZZgYnwWCwjFCJKuMmVme2HDBneJmdAgiEgE4XdO53/bszyb
4ttuakB/IfyzaFjavFQpjtDiuNRVszvBaLWgHtRe6hcYxGXJfzel7dZh3n6y78a4
ZDxmqf+ltgGQ7iXUQlg7P3qFiQT0LuvST32k55BwEZvwjTg5/ebEKge6HlgPKvsb
Xjl7AneA0XuLuYuIAXBL8rMsVk6ohrAhxcEOZnDdY5jAODNwTsIMsIFu7bGHargy
LNR/2GK57dg/lUZ2JAG/P4ALTsIqxs5pBr52vGUzJlCt0tltVRQugLwZ6xvFFABb
hfjEAzNQ1LTHgaXtc/IqudFlJDWYn2lDIX09l6BkoAsPrKluH1t8ul0BJ2IVXdnM
lkOaLEKBUDWqYMGYbfLIo0R4lm1VZ6iRtObT0jn3k1Llo9ubAk5zN+QCIaNKuo8n
9XIm1IB5o7biB0VJZOvsX4wF/hYh0ehR0pDyZYTKTMKsPsLuEWWlIdVBwyZiB6M8
pZ1bR1/id2j1uDHX0sR8rpTOc8crB0Ppj17jDtp0rKNmp3L+/9A1SYtyHvRJAyl4
orr27IV0n70h1wYJ++m014ciazrZBJNt15s8Q8cYC2/6O/YRi1J2eqde+lq01Rvl
t39E+itiaJTavFFzMbgQMKb94THAavCAuUHqHtw5vNF9VwXOKYgfiYs96L43q8PV
RLLhw7jrTlU14lxcA7SYi6UNC8q2XKHK50/zyvM7pVYPxzbAvphrY8P0upADO+Vz
h20ZMXquctwMdg8glx5ANHsj3eXj2DwzEaA9ELtCvQhhCR5XAV2UxeC/Qte+Lhvr
4KnoujTWVwLbqdtGZvju+EzJmEYoDGQ2+EbmShHepE7n8SJIjKVtFCqjwNs7nQss
UjiLG7mgfcaIFK+LFxFm8Q/p+Crv+3mIWmbNxSEnlNa+uh8OpR9pqVWPskGw/3dj
XF907cTZ3l5xj/mO3sdqhrHtfHW3/WGkmpL3JM/HTEmAAIlBfQWSAm1HKF9u6Hbn
PbT29Cc8cJJuaXLktKEzUJ+9ADj1oxDlDAmkmrZTzSw3S8klH5VaVzxD4Mv33Gce
Sb3Z9WyH8TJgEAR5oc/UOgjudfCZLSSxmbJx/v+dKcnM5Lx88kGqpDjz3ONMnRZz
IyGWkur13dtGjXHAx5SkvuRhz4rqQna07g+CZzA9dhjrcBoXEIPdGmQPEUAwbw6u
NChrN+LXdh8OJjuFCAnFKX3g0Y1ZIkSmY/SiKHbfQZ6cSSoYf8Q98qpG/zirrywB
3vU3F86pLcjg08K3XiOyvJ/5MAD3eGq0/tQ2dB+kO/YosiUX7CKmU07oeoBt1lgD
SC/X8vqo6Uiw4Qdte0keWdzSKobi+JBdkYqugY9ApXc1FlwJQvo9OtVhcSKJ6NmR
sb4nqump95AoR5da6qUzmVdjjpa1vKo4bpUH0fQgKrhWzsom+Qb9At4w5XdvJ7Au
WKyz+VjxNysow/UBFdHmdxcdqSD8ltZnycVQOOA3NRvcBnaBnIpa4T6bZ+hN/R2+
oTkK7+zy1ULQD3OBTt+DuSv3u8IZUeO1PyNcciEiBj/09UmAUrDUEYK7iV8N9yga
xCANcFkMHzpMeo7afYRA0It7e7joJb0uJJV0suxyos+lCw8cV5hAGXf9zkLem5lq
anvmdr5TXOmWjbItwcjLEkWRsDCycGuVlVvUtdBTkXN7KEIKToWgH1d+nT1/SGCS
SS7brnEhani3JaoWY4LxAPLounmZQDFNbqEKnFIAeNjJTRY/O84knLagU+qVd4WF
F3dPMGegSvavr3CsVZjLW5t5f5yLopI2FsWuqCodRMV6oSkf7MypJhd+3xVN/5LX
vBpH7pwmFs9N6SQmg+DL2TmW0KDOg+DWljeKFDaQ9bntJUehGaIi9qkmDD/V1jI8
+kETrBvmFL7pSLE99206S2RpXQcemkcVj9+e3uH4GQE/DtguJAfpLoU/wMfhPMA4
XNPCNnjBQoQ+LkE1u3lC9kd2aL8pPgav6QUB57SrA0xtZnj6PBcJIOBZcV0+v3Jm
X1zgSgOg5WocWE3Hk3c0Uf5pk14FuTlI86gDY6Bd5zQDXvoW0SOL6u9OrAJwYQ0G
0wzZfGj+AIcUKPalTYW4drB8r1wFMBWpcLysARcyJvrSnd3liz3SbVAYzE6n/+IN
4RKyAVSmRkC232YPwnrO4FCFD9nhAfr2aKk0hSOHzwzkz6MRfl7VTgzAKChDW4QY
DZ9jrPjFFCABjNj06TEJAphHUrYN8dyNzS6WM1bvVk+6ns/fpyp58Xj2rcbX5Bhg
HdDHYoIjWw9cv9V1aT/joO8Mfx3N2yxtro8BX4OoWUo/cduZFEScyLwLBarL0eZm
iJaoOMdWWle2+gdV++D8KZvqzBlWBzRlEKES8pVJlUw35pNrG/nQ3Y0bs5NeZxQ8
QyEb5pu4x3DyLXuI7Qz6AIuGUxFEMhgFjKEoB64Egen1T/tFZDXGX4sO9gn8fJ8q
Pee1VvUEN2OUtM2ELj0IuDJ9YhvY53Uqs4C+S1mKC8T1Q/pEhVpPQxUqEDMF7wEu
XuEgi8z2K4ZzhjpolQUlr1wplX9i20GO6Gyad/430BOxDwimxt3I3veGyRqGW15U
WnmWaCLlVs4f4zsvrGU+6EcauU/7y2A+MWhlekrGCq8LKLQ3bsfIUsCowGlOx2Y7
YznywXqkShIBrZBqs6SXJP20PfCBogcTu7KCrnK0U+/T/ErEj3imQOSmbiI01CVz
NebFc2YNgNJ8paIbsD++gfcG9oBa1YCiGgbyTfLYEF7E8Rn9xUZ9gZ1OpiYgbtjj
293TL3gp72bnS4fTaKO87FXG0tmiBurNHvyQf3PFeauyJr/viPoz88spJFL3ScMV
h5V+/+Shh0bfYapSVCzPdDf7F1RrLnVdfr9pC/8ByaKqDJeUyPDEBWw4a5wCkMSp
zwvyRDCIIMUxc1D+7RVbvxFXuOIaT1Bgddh8yVD0a5HHxAVfrLE1TEZefBef3seu
eBsYcQY4ZAuh/syX50hdHMQx/l5JFEAnW8DE4/qI8ln9rIkVaeoDT6iz4oAMZupx
J4HbxeCg/L9FbyNRWPPkE03IHjUeLKJVOB+ywCk5vm0o9j+O3uyXrhb2RKUmdbF8
ATBX1Wl9EDLpzswqEfam0zyOBz8bhKfAIc8vjRu0Imt40jUa5oSbNpKUIYuIKdBp
6hJQ7wYlcxQdgguBdhe4RuifVgeh2Lm4L7ImboVbSb4zBlYtOsyTQ+sCNE6Oj+T4
Mkw1M6Lejis5Kd7MdncPZox9wDx1V6H3bqU8Wxs1kv3jQjAZr1UB0a2x8yvpmGv3
ROr0FKEAY5vj81BwCliov0ASr5sMgsHBvJ0tp2qqM+qup3tuJQrVoG37syWpt0gE
a11D6v9PeYM9zp/Hw2NRJPKVOy0AYFJcKzTR9CCbS2Mrb36UcBg2/ceXodj+YYnk
2DqbrQB2RV10/JdQFvgRaOuS6is8I0L00db5ebMVLSaBpAx4dqnad9m+zlaC1pKx
ssXb+YIUkRlA3TB/mGv7gsj3++7G2/50GM972457vcEv0K6WSPSA4W9GdaJLSK96
3NjgkLZCV8IJC0zm/RY8f7J8MVVR0+HzpRUd/sQYeZwoDtyfmE8X07jE7foull6n
SoXbwbtHFsZAU5G+HieLb94JqvvPBTbJDtR1re2GlmVI8SUNlXlzxMSPv4bvBh8C
LzK1sZYhPFCJM+HxNvfJKV5gPpsJfqBrM2OfUMX78iC/3LPlJ8M0U2NXl0uzxc1R
0bJCLH+y5J8XJSSnldYfnXJ2kjhd4I5CCJQUFFixsxLjj/meMjyepQuvPWMkcslx
8WOzLl3BZ35Z6MKPF4z8ovAKGagEcpePKkGgOkj6R0VxLw6AcKktEBWfIJYgiRjt
3Lw/cvI+NM9wtNu9ttJ9g0kgO7dt2f+Zqllcu7xSkertVeKG2GhZapqFvIvAqAlS
3KNIWnykYmqN+NrrM/YDVpqIMFj6c0DSvN+utOKGLJcwRfmvmAuNOYn5c6/jXNG+
5/RKmsWaG0OUhuECo3TyRA39ANutX7h4PFrAJcIz6trlz0Nat06TUD8izoxDT0ES
Ha+2coCy+ui17N4xaN9TadH84Hwfd3YA6V35qJvFBGLwTGjGq1OkA8DqlguzJTLt
hnQlgVd/CiUARCunn6vK8S8kDUbZffAYKmEufLfJpjyWOsydj3wqkH1CqkduU2bM
QAkIvpws60ONTJ9cnxakJU1ECmD6YXF1FclyxN29AWCH10wTdzJLbW4h6Q9S0BwP
veTI1QRvBMGGrtQoezXOVjQyyFMLSZ4fLteMuqcxHaWQdctFJjCzVcvuYE9CGbwb
GjFInkt9PPKSZDfZG83hwhvyIBQFaQmceFEoq9oAQGUPW9lHzb6x+2n0zpjBLuWG
Hw4CiE5C2zNx9n2kwQlet8gvGu5X9ylP7eYkbqCxee7nnZROAgk6c/hqvxKk0etD
JdG9M/Ephl56zXe3vmUHCa1XdrcKkeN06Jr4SN1YlsX3IKIn8w5fUumNwByEd9tS
TARmJUlW4J5xELPrdUFhHc/9OgbZjObzlrFjp0vFJP8EshA2Q6ED9hFuUNkPQPyw
vOjuBz9g87SyOh3uUfsYuo4+KWSMItgPajn21QBQ/Progdc1gL0FYjirLNOe/pdr
IJKb0+pDRNym8LMseK4VJ6vNkX/iltBaQn63e0uTDo9uXJ1c+VADl3hUuCc7CCzv
qEo0TtutRnHylzVZp8zIdgn/WbutnIzsCBAmPI0OesBNPItG+DEFoSsePre3f5tK
NKlXZoGijKp4KXmjxihstHyt/V16HwmIOXBBimEb2DIZu5r6NqFNljSBjIqYEksv
1r1ckB02nekK0k52QxwH/eT40RZ9r1+euVonHzJQI5cU6CX8mrB43LPKynU4Vl4o
qLfJzEXmk9l2xmaryrW4b+yJoR7hnKrLPx1VSKLjx/GDkMnz97XmlQBQd4uW4uCU
murTfuJaQsOtPKILFQNJTdprPzeR5RZ16yBnZwSWJS20iwhsqzCLvqY45kDuKR68
rdCUgyha0Q4bITQfUBbOZPw9ZYH6eREpv8r++fQSLl6xx1wd3eNsf/t7PB0LGgBW
QFZKEjldFFyg5/8zcAUlrwl6VX+U8kmsS2LoP8hC+fJ2kqbuJeG/7V897cK/waL4
8gqS11FxKOocOzBavvbgVHy8afFcV+bgSItZxDeY9nSaCE2NdYH6m3cogjHFAxEH
Ktd5mwcfpg0HbuS7SA9pqnV1rDm9RnnOjDVhTX1XRM+Y1J5Que3yQjzVq0PMNjGh
WWpMkxK2KWT34Di5otDQC/MkSxY5z7VK7/K2xefhHnLeg5RA/ftpm7KJVbwyag8/
Rpr2rx4S765o3eWlfM+Fc9zI/LM5NVNI0NbAS6Y+YltWYTHR7CGMhN/hFzAtEiKf
AYCamXBmLj2UAIW8inMnAF+2XSzGWdNAlObbJP8DNdj9tXIEmW3F0UuQaDPyXrEy
PxSkaiKygGH4l/HEY4vcQYeZPYOZnnqawG8/Nyyh7+BqxeuS30DEdJZz8pOyXdjD
Z8ersKUW1wbX8yZPJGw93Fig+R56JNO9qfH6EXe77CT89945sV3JHU+bbxRVsaak
KS53Ivm+GuG3spteWi77vq7K/YrMO+hmq6JYzglA89QPYj+ZuTBDz5FLfPtg569L
z26Bzw0FqVc+ezFCOaJHqODgSzAwZG8e6ZIS7bNtsjAt6ssPHJigl3kKDGh0EKIn
tZD18WrjqiU6hn9Fg+O7Vfw/3cnKWgEczX3U2DvqRsrPikkMfGzvSpWKe3Bmv2l3
FlZ3Omia5hx0TxZLinAp98KrzONX5TLbdL9pQpL00GVn9tNqWCVZviGpm/i3qNpC
7YsZg93+c7h4HSCWu8mPcZv/g8z7nlpqfsj8JRynJdlXAI0WaxJvgdtJd0X14IqQ
bzseTmkd0snxADkmoh9zJ4B7UJ3K30AK939NZDTwHvvMcyeDIIZB4XPYipSUOh3d
zscVpTTCjtc/CC9SL41Jrv0zcqJQYWe78R2d/dD/OMNT64wRk/CGBcw5+h/k7B0e
26mALNikq5BZ6nS9Molr+v37kIUpsftKSJ/eIVl5hqWUsfyFa6l6DtdO30k8DOeB
9aNixIUIbrMrEUN2eeFBn+611mZR278CxIMeiPycJITLbRvKuJMMTkeDDo6KWW6x
DPriek4oFK1C0W9WXBhbipa974lb5pQAzcICiD+MeY4ho+UgPBaFwASLJS2fxCgZ
lfVum4WJjIqFxUjPhjGGev54jy1J5uj3BNWfslVmM30JByJoNoVZtO4LfeEPHc2k
+Tp5gYCop6ShrhecxNUwAtqFcK9ntsCp0xMG1M7kqEiPf+GcBGsh8CX/64P29eIt
LMUVeq4I+8gHjqpXOD9dO2u2zSjGKNJGdLmDWacvirGXvpbpTjk2eJ9aXizwYjQb
8XJwi0+gwKy2ST2r1+pPAuxmZ71FMYdr3wuGhOpI0VAKZWw2G+exo6ugR/7BrYXo
pa2fjL6EobPcfTXfos/PNaqGvQJ3I2yRHuSk8FjTlbK/+8sag9+tPOwhGEhfhiRJ
tIiCh3eTg93yFCp3eojIi6oJwjrVbKA/hKeZIpvUEEmBPG+6rTyCdGlgdRmMaUt6
9crlKWMIsnkILplygOdSV2lCGxvncY41gEmrSWZPuJS57iN+mNCqWcRrXcvbiOD8
EkNyd0TsgTNyIofB/cIxIch+wRCTxAdMuWM/FpFGWjXokMWKoTCSclHktXaHO6rO
3AT763a+Lc7ZCq1ORRRA04WkwbPpoWW6iVgkgRm+npvabZGBzmYuJp014YsTAZkL
X7ik1VW2iNXwvy3HoGLaDvV7MhHi7qbKgAp1oExZk1o8iu/buRWC1KZsQls94z6b
Xnsb3ppHD0bwKUHiQSOIOVFKB3Y/wzvo3JxuWY1mLIZQmM0ZIA0YqsxCld8LTRDg
X5J6S4oj7RgLvaP0cDI2+5g8gS3vBZOQky0hO1VMmUwYdANvUgJG4QBHMkR9dsKf
FzvbnxHO2AliPaPyygGxdkHtMF7TswQ9d+3ymkOQPiVOPcdOSi06xCZoVg3in7X/
5Zflei3Cn+eFxmo4YgoKPhVlBzQTfkGs41/xc0RC8Lp1vuf77OUi8ei/cTIGd+MS
zI/OlwkuBMwj+RYrlzjS559s1u/K0kFmqVSJPzrSRyr4Yq5oJ8gWs5BPGilZosTo
lWkjJD1W2BBoXxPL+eOWIJ6dM//FA0RS+KNuDHibvYHsRqVrw7lhnsQFXqFpUhHn
57MGMfMVCTnE8xEX4G3u3Hjb9U79dPmMvmYpdOeqK2+W2VfoALORRikL/X5AtuZZ
HDcGF5v8M+Aq04IMsY+EpXUQ5z0cgKgorr4KMNPUuqt4PvQLsf0IkqRc86CJO6zY
tYM31MgpwlHEip4cvHff7FjNA/Oi3+/eQdkO03RLdFuiJefgCpyLQyO4gvpOGYpH
3uwaEXto+wI9JL6o+olXMUsqgO+dBdvC2gOuVmYHKjORLST3/M9LMldGBTldMo5A
Whq7pG7102ZvWY7LjD/BJwKntOI3feQtHrU6glZD5hSoElBCE69+shAfDbF3atzs
iJ1hBlxmpB2qXEZg5OXVUxzfqfyn77DnXHGpHSMoO3qJ+nmSmekGGGVRzlBOhP4d
5atbgh5o5HdjX2WV0Dga/Yo4QJgXxlOmswdVVW0WmXqSqfV45OG1CwweTG3K43ji
rQOw2Z8fiTwewWMccasEzeQnBywGk2kLJ05yoxZDvjqvwwMzzNHdPb6JOaduDHTr
Lv5gxaGQ8OV6UVpaiqfijFYx0O/sZlE8fAD6SPwjKYqZg19T+WNMFZHtrMo5mThu
w61oOrlyA4YJI0wsB6vJpMoenTyobgNJ+HUAY8YJrwkFhm6UI242S2EzL35A4//J
lmcEWHUhYu/fINCjmZDm4Hunz0epaaeHc71InPLEEGHpRZo/gFQCbC6tOjVRhLTV
fskkRTIIIWUZhxD0+WHaGNxvIn7bs6D6Wb/su8PfVVTaCYbKHstZyADUz+dM0EU9
A89U3k53GLVlZ91hOSDQEmO6ricikhneAXvpvYd5bfhM2uTmhNFvs402ucdINUa0
KeZwOs/K5hcxrpm0J3IeqZxuD8Fn/Ds+pDxNlMpaQMLWgywI/n7SaCbLwim2+S53
w5ATX2QgyFLIfT8EqwPAuXuk++no3kMf3prCL1oEytUTI3GaZuH+b629g9KIDEGO
EzybB1h+UEUzG0YA/8wVpsElnk9/vF/lk9IJl6vOhyoRB7QY0c/6NEK7fBW239dk
0gKX99YiyLbNVs064fZdCikqMlv+0jv4ORBLDWqIYPhSfMu9y//yoBUPOy5FP5HC
86sIp2JyJ+00rpYXgvpW3HpKa+/fafoM3ZTikDCrECRRE7W9XueTXZFaq23gVsiS
E0gvIAyFg7JHIfIjAI5sEgDHEe8SujMnQaA2Whc5O7o/fFX/9u8sapKv5FvLop+f
kkY75OmVdCDI9ixE3QJbQi0Smg+ZiciP2KjHK0TPIYssYVnhY9q1ZzGiyFOUja/g
wyiLsD75eQuZkExq5YPuWNvCvth/vIOKrH3o6w27d6esbOcJpmYTkEvI0D7T8rB8
XNRWIkYVnknSWMxHjfzFVh4CasKNCIKR1KiwgHtCbFM9wRAgK+NxpdNbbPt/rgAW
hdA59vHxbY8vS+qxMay3plrcekXablCb6DlUSH+QNxRmNEZTfWKyTjTaOeyT/IPf
MqlEYbhegHKjiIBTjc2ToOSt+M8s2BDUtz5ZIPS7O/utZtDF0HzKqYlUyS9QceoM
NMp6ewiDMnde8EbPIKjc2gVzDUXxXXUdwit8QoxWT/apZylv5V02/AXW/aXhvdo+
B177j0uWrknHX1QfYZ+3RThC0WlW8ZndOxEleGaIq7yx8TVJM9WW/D3wUU0FgFaE
H/wFsgMniIj7XlFbYpG71YLbQSVMmJMTV+loBGEz1QN8l3/0XmkbiOb35MnenmG2
6GfbZnhWvvgJjlZ+6oY+tluCP5twEh7PA7alb7OtDVjjOWoFH17VFQxZ9nb7Um+n
gCQfc6hRF/frUgAPgIpfEpiuR/35sDQByoDbM28PnDEot10mKEaQGeYuscYU6UbC
aoQB66gaUPHh1yIvgFxFk4DUdKd96qEqlnHbRd5aC1iJz9liJgVgZBbtxsJQjIhx
R52C/wZzQxE2kyr//vAw3Hu/UgrTie+OjNMZJZIaqvPNjtqfNF6+Zt/BKq6DPh6e
CVIyIUx2+fcJieOc67AszJ+f3CM5fAxJ1dmWd+0VBoRKldjchK0948n9jdo6ftJA
QGYI/Ct7BJwobJ2bSI+Bw8wrhVkJQbmQfmMEeB4XQmJVRwogVre9O6ExIVLGzlsF
ugSt1f8GraF9R9TQ6DiOFge5bdnC+iugsLXIT2++ArR8XUrdpsp9Fv1C0g63G60+
P4I0Elf2fkM/f4Cze53WZ5daMyWJKlQJkoHqXUEbESZXgYXtLlmiKabODFuRQ8jC
WU2czaeljRXWGcwsn+KOnMsBoUSFocDqEUDMwG/+jH+Tv6ZdeRapgC8D4+D+3KLG
QWEl/RVLM/u0qdaIolOiCh9lB9iM6FEEuvBX/Bp5QCH/xHxe5dqFP3eFt75j9w/s
BPC659lmDzIkc7nVN85wj0ue4l8ZgJE9ZIUtOhLg+9Bwm7XnJ7r7TOeHEQyoLjET
okIWrkHcnHwb1eAbBcILCen7OHZWKHycHxUv2V9Z3uS726wmTELvEooimoV56W1v
nFiqQbyvy8CESY2Eiy2NI4EEqQKzCGNAdrlKlo1NqG7EXGdIt+ALiqRMLAuL8UQB
Obk70vOHpF+Zfo+MYPnfJRNdFOT4dK3pICx7o9a44uV2OgDJvBj3oUkP5rYJ2I3a
j9I0x0R+N3GjdWCYXdps3eMclJ2ir5IPUXJI9o0cXcy4p0/RTQbQbue7D5WZMrIq
kvNVAsiMWsfe5S6XQcpAAipd/UgnJAdRapR3D6x0YKH9Kx2YyEEHPngWJwxoRP0y
O1sYYW9eUIVVlnGs9QSLvsNWHRatcaZ7qCEVH7E/5EVCUxonw+83JOIqK/3ZNT1d
RO3Qu9gfmRO6gCj6QCG8cW+2tGLps7z7uZW2Nh3/4V9TKtMd1rsaVilFEGr8Uilp
HxVdJhx6ECR9VrTDsAVQb1wAH81SZqbJwK2PqUSX4xyr3heLHQ95Jf550Je0qA+g
VztP0lihbsU8j6NpC8rEHD+snG/z1E0Ido/jmV7tdTSrH9HzLigAcE1x17XC01oB
t34s3swGcbuuctsv5ER7hyKRKmbl+CGsAW7BAHWQAuDyEVSME8EdR5z5EoQARRtA
YSF+S8S8LuL/TcHOsdbp72XwLatkDJ6FkW60FsmzkWQmDssuRrbY3KHa/pYENIGW
IWgA64VHGFq/ZNeg+FQMkYT+TMszPYNtKZ/26dbSb3I2tX+HZkUUa9ym7ApcJt8c
iPmxCxrv/CuWMlJN7Eqkc3CuUqpQnjFaZCKdrp5jOJCtMuif56kP12Vj0tqbwimZ
qw38Z2weO9bqqsYhCtsUCDCME35K26g4pqb2epSNg3f8o0Ji4Fw/Az6cmKN/GrmU
k9nJnrthiGsTlQ3yHl0t45lFrLfOuctmT/3NAjpfK0QwUhxCzWmT1nN1qT9kG58w
6BgDXjP6Q5llRnrxHK+CKocS9zC/AYSpSNJGdpdtJWucvxh8qvVITVPU2yVs1fQ+
pfJEV/mKrEfqYyHBeZwjs6JsGqb+91koRH3g/hqolFpWGdovpmALYeFxn5ooW//j
jz+8M3gYKGLfM0404dC9cuB0q02e46RVfJ8G4Wtn3WAZoObfhLrOpEGT4azAg7hA
PJoh9jeCPeR6ce0x4yVceToI0iqP42JCnBHaqWNseoHg+23a20LC18eSH2OYSLoE
KeJKy9eLrt3SLvcE7z4GISjnBv4V6zpWmrEehTIZ8kIPLjjP9JuBHjtao1ymqTk0
KPEyueNjvYEANxBI9JeD8JudM4kmYEME3r/UEQZwiha6bHK+CyXVQvahJeIGnIeZ
juYhTeErY6YtnIykimRVpgsDRvQ5DMswEInpapk9ChnGsQgodgFs0zLXPFI0HnYX
pQiPQD2REMwgG25vk+hP8Qv6FoaE4zX44nFjfbW4ZYEXEAXabg/Em5CfpfCzAdlb
OcFvqvfH76kuTywp3X/BTfB0N4A5yjSNxcUIW6v57LMCOB7ZJCVhe6qT8SR28jkk
T+S2NUZQbSkjI+UzSC1MTW7nBCcuHp56eD+E+KjkLmWIyMyx4r1X3rPHl4IrJRtw
tccgAPHY/dKlLnDKHVRWJ7essV9YX2epyicDO9dIZjRNbtHf3x5SSsRttTC1ACeD
VMlNdF+6jlniiZbVm2zTq6KYdmkAB+5F8TOa8JLKN8/yWGxYHRJdyUU2rBlnaIDD
N2O4fwlh4gKf/bn1R1YMbaLXitEJYxmYACyxmZdr9WpWwBXEQQ+wE32kDUc4kXSG
oMCzwxrUgLp6UF8KQulmXlYi7JSZT5W1JSh2ON8snWORJ5LRdjv9SYXivlPqPXvg
fgfpeMhsz6yqz22OZBM90dGx27nPeS7WyhdeMWBGqZJhbC6ijccyZixX45H0+/pI
w39oEc7DNkTkEZp/AW/g4Xy84hrlL2HWk6guqdF8iZf+YHGCe7Y9AlSk2h9DH9UU
IwyZkJQQABTodXfCbIeRL96pAHePFoJO18Z+TfvdnIBILA8FpZEot5KYUEAsPnOU
PkRpU9pDOIEi9suBK5yxtLfG4Q5h/wx77mFcweOx7P2EIbJpt9JmD/Wg8IRMu7pa
nSSh4BnD/xJr/xGkKwqIL/AYYtD0z28w53RttaUuFVr0eDwhLCx4Ks5T7n7hhIM9
QrNxPuN56+gkANDWjjwT6CIzDCnvBd1Wj7Q4pwJexx1tyuFR95Bo6RH7gIcWBEnu
AetGZ8CvMANPpkW7hgB/XIe/4Yr6ZCQ/AkfFo+nitER3T7acjXp583NzI8AgbHdP
6hpPQm8y53IuW0DgZuTt2fXVZVwhGYW2wj2FPQ4+Ncq/PoNCc+fIAEki0tSmG5Tr
PZFTV1GTMnmM/i7RfWFENwzTrbsmJvF62LeODdANrRo2Bo/5WvIs58xNxTGYnE9H
gWJFXJOHikNdmcCxEKkc9OwnmX52DkNw6zv3dv61ppK7Ak4pJtU0AKUQmuI7Ad8U
RPpn1GngHvReh6JerVB1w96xlbLB8plZQ2m4MvcoUtsQ9ybPsiyW+sj9Q0PjbEXd
afL3GAEOl5h+5Jdw0u8SMZ/qsOsgSn9svImEW72Kcyr5FldihdzP4bxRp0QSSxcI
B8qYEjTyEKUreeIbfHp8TGzpY0V7ovvbPBC91geitDVMpcVYp/JD9Hp4GTYzvtUQ
EgSJF8DXTRBDB8KMzR9LU3ZG0syz2kZwtKVcgkpg5N6Fhlue1j2epCOd4kNZ3HFm
V5LjgJ2EOxcJurGRDwobOQnQ+atDTxMBIlKMu7Uuf/CYEG9QEeToU7o/vTfSH8YG
VqrGpM5PZxLmxGsQOg6GcapHDzvwW4muJpDQwQoDWWTRVPSS45ckigtKTHYiIClj
iPmlr6L7zUNZ5S6dppKXqJtPfa8WWcGMuZiA/5sOeGj1sgOgyKBo2X2xR6x6sbm7
x1DbTUXA6Xdv19oTz/yqadvJ+F3+bf4JyYxWE/1YcLVDcrr8Q1Pi58CPu0iAq3hT
KdDhiBLHjB4ZdtDhyHbXVY36wxygU8ZzMUPzLvzrbKDFhFq2qn68KJnZhqC9FJ6n
pQCyxa7GXuFcozkPQufMskOxofUazYNSK1NubZim11Mhl69Lc6om1EYvatSwu+Jv
hFGTOCl/xjkzuTC+RSmfIL3DLQS6kSCndQUA44CysD1HSBSevUYNgIHa6odWa3w9
KI0iWUZUsEwQ+QZLuVJt+jlPEwVdOJPIHjXRqCkY1tODdJ4EKjWHElZANIwHON+W
OnKY4sjJZlVE7CbnxviXqmZlVgDJrLYEtEIJiC46E+bjW7v6e6KFnHVuzxcZWCkZ
UitYX/91YlGqfaN9MLrCpkHXHK88hR+e5cjqa3bBYwjfsJ4fDxP5GFlfE7I19TB+
r1j2WPWpow1r5rqYF3mwyDu8mERG7si9UWaWL0tfIJyWiekcbbTXjMAN61GWnFI9
2SevKbcGIa/Nj/7EVzEp9ifG6dLMxlId5PnK5Jx+UR8E1T3rOuC1S1XYBqstyhFZ
h4yiZ+Ai87xydtuVtmh1MwGE0vLIwN8cKn9WCuAp8VJtJMzqEZ2+opvmEcC8go1N
w3+DK4yujrmJoF0/qVUHRT0G87v9GT5lApCFrGxBjE7S4l5yqq3POHBdl1d4X0SS
O+vm517UM3aRm4a6bsuKId5oM/CG5zYhXR36vrRBEcpmYarJK45bx21oH4ERsf6j
YPOwHbZqPVp7nRJRiztlxQJRdc/HB0YonU4r1j+q+Vg141EdN+wibs6G16rJm2OT
6JxEj4tJQirfUox2q/x35CcKaHtq0S5U/4sGaeCbbC+WlzMhDo7PP0oCCCTt4I3e
ZRBiOhYdGbin04YT6SqSy7Z1iNKCJL5ZoM7/P9WrCYwsbiuu0IO0MEHUsRzkQdq2
WksYlh8FiHTSBncKcPy1BujC9sIfd6IQl+Lq3c5jc7/i3OggLSV5/1DUAKcteTG1
8DyB0QGGhrfoTOKoyrzYtufXbkSdWmrHgM1NEnPDb+bjxEIQS9GNehFpv6CQl0xF
hLdUQgcH9oPK4/B9O7BwVzitMd4BkaeB0brTW+v04dNtAXw+HDb+6bHzc4L+oki6
g6b53FAHg58ZidpKfVYGT+/mQZ5i1d0vtBHvZLvYxWuyim1+a8Gt2awyBSMU4GkU
YonoaGgLoNhZ/4ZUOMX10TKnG1gQgQJ67a8bPkl82FttsEvLRmYE1jkUO+OENpLo
voLvnbRX3cD2RYyI2Xkp5dnf08cs25i31L/5ItGpZncSR+YN1fJxVNFDduLGjMnj
2BgOhLvQCZA09sBM13+ZzKT3ny0zirnWk9AiQ8yzyq6zR1zzcXcsYXJCg9ONlJHf
Bux5HOlExDcCsyXzHUileL0Od8GHF8MD3Uppjsohwpu3BDm5c/dOUg4MaZ+pzoef
xTEMW++4G+4nybR4ehkjT/eM5TJVmWsfs0hLQyp5qwAbKVuAzwDZqCo0b1xtyf+H
yPVeTYRxZf2qIx/o7xhioAhEXnhl8FnTV3evs1GBn+bJsofpVxWynkuIDdKwHRFg
S3bRTdQVlt1nfpDx3mAAombZS7UT6ittFHKPHmEKpqy72eAY1mJVw1ZwDN4aOB6m
Lo+x9RxgXkw/Xb8Q7v1xGmU6DlJdJFF/7y4dPVagRp4/uhOjeEKPGEUSIf6hBpWv
7cLR4Te8D7smPG34oyYnpNdUt9Ii8MS010l+2bxuTnm5/wEODrj3av5Z3bRUslsY
vkSzsSi+gqoBkFkAGV4hD5WQ0cW9zfh/lwW2rQ77SidTo0L5VyZWroZvdoxtQxVp
Koxo5UNKxUWJ3exadyIQ0oKBDVw1mUWhlViJwszw+eMAov41IYVAIPeRiOl7SrCm
T1n6Me3b51BMGraEJ+ymumkMIbs04W2y8+Hura/4tJkcqHgMnCbli28SmbnAwJtE
jBUYv/TodiCxhR3qF2F9gtgBrTpkZWuknMYuOCuupd7LC5T7yLMRcw7yrQy7bisK
tJzHP3aueo+fgMINI5FDSX51YTQn/hYpawo/+aYkKKz5s01e4dkQlDdBOWHr5xTb
lYENC46XAvTL5BaRDYd6JORJQR+tRBbBLldB42UAYmY8q5WxkwPuLwQTXp+qNNTI
yyw54svfMDczXZuFLm6hqy/tVoJ+poAJg+wbEHFGrcFqPSnyqH4XPKDvJzMjZsY4
rsHJD+kHdc59S0mNl97wQgeSMSSkCNnpWBagSR4zUJ41g3uSZPTWMHaU6qZ8PK7q
zMS8PKRpvZScT0DFgasOncaolcmgMrgcx7f1Sr+fPT+aHQ3zDSvrGPjYfKto/m7E
837sWmoU0KLvoHZI4LnPmemHi0I74xXlhNjSSp5JPnZgQjh/SdeP2kTK7smZ5K2l
GNd4C0u0Ptt8AuQfUxK5pLY3clOo7F/rdTB88ZjaQd8AH/SnL4oDVVO+voWIg8j3
1wwLBZs9BqXBTsKp6/InHl4cawRtKJpZC30ocylSEWdQKH0JKQyGuKve/B8tucu9
U4sSC29TMWrWbnHsXWMQjqaxXA1nfFDwtrti9BDAmdL2+5zIOYmV8VcAUs1IOEQU
0seGuobhQIsFTZt1JQ2Lm8FGvGRwBWL9vGMyDXZObxGaglx9Vg4Lynw3U5o5WQl1
rA7YevzQrf/gFtUJcHzZ7V35Aar8UYSk8VcneSgvnOsnbpcCJqIxEhDDXNDCoZvE
0DatoCWMnC8M2KrSuuvr+rS2yFEkhK9HwKb7yOhZzg69TgnQO3c+7v/11kLRRuDF
rF4D8Zv0TZIEz8Gc0BfJz/TkeZ815byqpVTvO+/aHThenPbnsRXMbAEw/7mPswo6
1Kpa4BmxsUTIJcGuOh4EOaMBPlb88b+G7InLyOEr0YxlF7+jAgkdiWQBC72ZyL8f
uoQJzBKF0xs/PFm+WPC8gN5znmUW3kU6L3RejNqHbrdkbfNATBOCdJq53hi/gaT9
VDDTqTe66rSH9OXZaUrbJqgxEGIIB0OB5k44sixFMiSmFpcPXUmP30HSAmpSMEP/
1E/rI5/Cam7sSutnfy/7G8Fg6oSYpMUwEp3RhHC1LEKzz1QDrj8FcJl6QWvaMLen
qdqsE5eSQtxVOmUOUOP8r81OBXZo/W1JVz782qjXBu0rkxiI4adVtjzVL64jdBXo
yH5QrDPA5cHwGdiNGBrOFF6egmGazYcg9J6JgaQ3J9vCcfNi9kVgRQjJuNOSoZDT
iuV3qn8JW0NAv1GxEL8BcOr+NmTjnPmCnLI1lWF/7CDtr0fvO4HVDMXa4B6RL4eW
78MIF0uSoLoJcgQoQHsZVYKdNnVuBqBVEEYRbr6I9knLtMYUoyOAZoFHoIjMTgJ4
FnbuWtjZpxdDSQ8LYHGTWry2BRTN1L1drM9ZYaf9SScfB89P6JTsh7PuYJKhei0j
ChtNimsPNYmNsyRHNk+jCATvllrlvZunS+rTA5xHlHA1/JTAwL5ncBpwNGnEfsH+
yr5fe7RhzvH0kifiX1LbNESmuilLQjQ+h5Ropt1H814T7bdLDAJFVVVc7gyvPs8t
j2haq2siJP07SfLyhLH5bxBQTRAc0aMWPCuQk5FkMHeZcMzLZYyiIpePzNMI4Ari
wZt8Ds03t/xBdu5Aqn52T1Qg0UxiQ+gPv2xB4Z2qWb/t6u/6xe9tsDCyXrroePsS
B4xNC8/p961Fk95VTEwUl2zoCTTsQlYrDM3wX1at0hlFcDO6plt//+OGQnbtU90A
InZq+QCL46w9juG3WnhfdmePHPL1CdzXEsQxVlcRHfDy9QyO0nyvUtxhqwzOpGag
XVTgLIKvSuyfvMdkE/nSCOM+Jns1CGDrH7w2hYoMRjoRMvsnMWmobQIbj1TZ/TIC
6NnuUcMyln5er/Eghcc/a+yUC7jwtgD2MPZGli3vgvyEoPGataeyxnrNbQ0KH+CW
+lAWHZ0GCBCb1nsrZlR0zwJINffwR6Hb/jgXOa5uMcNBh8m9kBa2KQaWeYmz/Glf
ux28OlXLD576RFNikXVcInXLIA7DG8doegLoY5Pl99+0jwgjB1R5LpkkHAWvQVUQ
uAqTnx3zVwSZ+rDMnvtISDuwsT4DLpVKfHXaLkjLwV4kZQZKNruJf0aF6dQ5c3+g
nra4nWLeMg+49lCGb/gmhzTAt0yqBhXHhOWBmXNFZwlzFF6PeG+MkHabRtW6OrLi
+8lHTjEUtQ06q+MRpHy/B64wAvZ/ADGgerjrIJJkJ58Cx41MvVASUfgRlO4lgyHS
QMo/kHrMXygtzOdpH4pycMkbjLXrQGqKX8bb2nXxIajRX4iTVifu7Drwu/gE6rcs
8AlLCSleCQ8MCN6spB7V8qFnUcuDxQDG4QWeivFI76MTzPuw5BTaIkhxeYy70o/5
Qv85yW6GIxfNhvNnLW4ZNC7z12MKtFE6z6IvRfycK2m8oFkukGfc8KbsFtTWPOi9
JzLUddvJ9JlQQS2+x8/2sJFUT9QY1h2gnP5D3rDxZa86vv6L1KbnKrYVNcVDm+Vz
fkkxYeOCOIqDKnqyPcCqawkg8fr1pkBqvUofwgth44sPBZjjWFHAtB9BDpaGpYWa
mjdEWibkgCOG6hzl0CJQwfwGrlvlCQA0KzHIMEcx8mgciAU6XgIregcN5m47p6i5
Nj/HVGk4UF4MBqHD2bCfhkcsaykFE8EV3KTwccMAPVf0AoXWtNYV97zQec7+TtV+
5AuMSauVAoNTq05T7BN8IKHSVvtilTyY0FonBjUby8kWAci9MiYM/HUdTH4UaKYG
qKDFQCqW8Cw4myxXiPQDBNgbXv+AfdiUJMTLrNgg/H+1qGA0S/ZYVEhZCENS0Jh6
FlIiM5TuSIYQ7iY2Cda1p6rCtCgmgxUopuSNKDUlBaCtuN1rUoK9X4hw7w2GCFbY
QujOueh4vXlP59LNICV7Q5F1scapDGxfsTKn0p08rXKQ9ENaeKsHJuW51/19fEKm
BnYYE+5oWdGNmG/Y/xvOjsqKSv2AgXNmuEHrxpu00sG0ZXPV5FhXEr6e5z+5txbU
miYTctuGTEPsImRo2tF6B+sh3lqXGC7sRHhMUSIxlUmaN33Mbgn+64DtaCV3l47L
VVZopFeaIx8XpUMwMxk1ZppKJE7yzKW5sbXMRvwmLh2chbLfgybgW70pvUOfqLkI
9Dc/tpA/g7L1EBAzlYUoWhMCgiUTyqMkonwQrleUcWySAwu/uFJ5K413KiK+l7ik
ZOLP5P2sVWQJ8medZt9/pX5q3lA6sq0EQAxpN2ExXfPZVew6WYSc1PbLXL8oz6J7
7MWAJq2bHLFA2o8jPBraijmAa2BrIKiwxHJJOayDaQNBvf7diq/YPPqOffLcqllv
mUJnbptkIz6T8QWfPJ21usPBBHXh0Aywt4JWyo9iWe+KX5+yru1MEJIyt8IIOLsS
GQcLXwUGgbBF2gg1g1yFnJgOB1pyvWFTbN0dHn5elhBH6aN5MBjIfcl1mJZlbLLt
nlDRCeLkhFnvMD5uKnxGKXbcplLD1bwMNC9//7zfCeq5c1g+m789YVEp0+gcHVcU
7uToGiAZnpCgbcQvx1NzdBU9Jw0J0IHZ4HOh77qfhzjrDELBZq/T9URH0gQ1H78o
iaRfA08ucAmo0Y9/97yy45Mc/YqYyjxBp1GgxayWsHOGr9neqc9b0F01iolzPBxo
foZZJqbnw1rjEq7mKHVvaBsSE+I/iSmcfj+ZaBsXNQ/DwX+Er+FaKnnGS8BV7+eU
FEYWCAdqA52SrYNDqcU4M8NxFNWXCS/30uwunikDNYjjhFCOIoN3Sn/WcFo0ohAz
aUGRk22vunPf79gnRhsPkJvKUlb0ggFYD0GaSedLd5Ha8WTYRUHMre7iglnsN3qJ
177CDzVDK+qoIJ1XK1dCvyvHsEDdGdfCGF4jpoiPfJ+ADGTmrXiekQzG63aKK/wN
SLn6u96QugL707AGp0CPMrfMOzZFm7VuNm3NdDu3kOStRUMFCxnUePgrb/VD5D5C
c/Tdq7q/b+vc4C8tajs66CuRZLGXz3RIZVMWa0INeUFjl7UM97IKHU87hF4zGWkp
pJe4eISvG+lh45nIYO5UGC+ZzhvkTlb5UOH+vioAiDKEdvWtIhNa1lI3twPBD7y8
fxrmXqW2SS4oBEwHkKmjdOegZFAGZAuokADWXBV0hFT2VljR0bvHEof/oGUlY1JZ
u8oKgKX+7+5zbjezPXrKlchXXKCFYoNc7rNDIQBI9PHfjKP38O2DVLvJ/kAZsG+d
7HhbwEPcAk48F0C3xvor7quqmlgpd8gGSw9X5/AyXACgu7d2ejHRRtWw2R7+SxOA
RQ15AvN4NP0p2cY5Dd1rqK/nO57dURSN5ohPxoB+XFEXi8e0tNueWxQrkY7sAIYW
mafp8jxCWsrteuwyQ+FOr+1VloYJpvaDh2LUTBCTFjO2NseV8QmUqRu2wKkXV4pN
PaHnBZyXIe5Cpvv+BKbHaJvuQh7sXEq7dE+PUGhb6WUoDPmbfvCWbVx+TUWbFQ24
yq5ujoVFWfNWJ3TJxLSm9B5etcpDrzCAf7CAD2c+UsyBA2pLVBiIAXqLps/3Z+8j
iE8EQgm9vKHGbZUrSn4FwXXVEikRlUWM1TMHmRT/5SvxIUpsqYVbqEM5HfukhYWJ
clSAy9n0VIUaRRu2GRZnZIpHhfSpuvBRJ4bxIl8071xt1uz+C55W5S0SdqzVUcK/
VpnFhY1xGr3peRZjceUAKtFuttQrGquCFIv272Jy9TtXt703OA6ZDObORyyqJ4WU
L0VGpcBfDmOFuxT40AS/KWNlxV2v4I7TJ4h4eIouiQ4brBkDbwVTzXeTvawsBu4G
iHixq/wjTon7W5aBIdhziCL9Y2+VC960h29zyo+9pVFDObfaNkan9KQrYiOqn0qg
sUjkWLNmJfOI0mDiLHRPAF37fCLlBk3FeNlY7LeUtHH/Fu6dnSAxMyJ+LoXpR1WQ
MUs32FWzLD+tno3lCFqTKTjNG0pOhrEXb6CwSV/8sj2V38I93xVN1LAkKV8ixG/8
0/U1vJFzV9Am6q4xU5xyFqICfXk95X7nqa7uI0oW08YQacEzxtCQDSw/YPkz6rZd
KH8i92iiP3VuquZ3aks7+7sf/WB+8oa4MH6VvvMd8LZwQTl2mhCIDZcLdJJK43fX
ww0DTGBQ6ZD8SkkQB9k0vjZzG9ZWZOpL1gosaIgQFMD6XNQJ09iMUetKKBmBaKc1
saoKd9lmSmRez8byryqIQ8JawWVY4ajow7SUMVUM0VBlEugjD5aHOqXsul/HzmbK
1eXvmNGc3cBvs7A2LH5ugzRa3FEC+DT0G2Ne2k16uryYoLdJ5bxHqKhw/UPLcLoi
PX4fdvubesaaT74ou9VVXxMez1Isk9wm5rrP/N9yW0llugGNAZvfcHR8xUA6Nk8q
ZVqI02BZ/ttxaFnmjchSp7EN48kx7S/Wohxhpb6NxQ/bXTzQoYvTulx+ASZphpwv
Kwn+UBuukKcQkLxLG0EVPGzB2ydf6zdGRf5+KyGwIXYiBCND9soAkNTPNUyA3JHW
Mbx3821PWZd0z+ooTgdYNYrRycfBfgRFSb75EwjXIxIuXVslb2i3TDXFnzItVtXK
2ePGWJT4SBxs8aMuZN93/HFY8vp7E5Rwel3ChhnI6BWwmnZV/i7LBUcQvA5OqVJ3
AZfUYPBF6RUwUrj/6EfpIDFzNp+ENKWoZZ4nxFzN/hr+JYRZyjzrZ0HOEkdOIBG+
KCuRljwCnEmecYvQqPw/6bR7YHNqafCz5VXR+6foHAypRTR2vfClKaf/hk8gtwJx
iEUClwatk+/T9sFd839iYdoYBwAM02oiTh8v2FrxLISrhQgAX1EK+AqGXDPTokeg
t2sJSvZiBJZLoO4AhRkS4n7dja4nmQGTVUTK2NOly1qBL2iNPYrs36qrqkGBV+YI
DxcLABPmHkUbXl3S2bOTWTH5RjFhqji2lu/MGPmxUQU12sIha4yVB1PVYqQah6N4
GdDlLwe2CV/erKhnN5KI1NZfu38oeUXwPI/QZka7oHY0NOD+OJB/qE/wmEE2/JWQ
K/BVQ3ZaLILV8gjkTVj1jVK0Xh7FsdgKwTtII7bimCkYpyi0WUaw5gmzZlli9EEn
c6+BUGAGF+BbMqIQ+lQn2hiuG2ffVYGRhhtvYdJ87GNTD3ssWnvaL6JTNjcVn1FW
NvE58NTIivixo+IBlMUaqmpi6FuLV6G1kZKPK94a5qEtnblWh82oCypz6purToRK
EMeHvk9wjfbQc2cEmQZqklRA8GArjMBVRdMJ0aCiHVhw3k0XxC/RS4lVTMyQ0dgb
Rq/4QRXDIupQOgvY2Buv3jd3FamIPue8qfQEZafuyMDkIN7ozzVT+paJ89VFtF5Y
ngcrnBNlw65x7D7ERarIXmy13vM2/HI5Gr0KPjNhEu+kcgzul48yHQM6lODaPWYn
0xcvMAtf2U/WZzQbdeYcC+Af9QHHz1BlIi2vnxiRtWKXNV5OZP19e8wu5vufL9Tq
/jgzypylCF2Dg7zPHSBJIk2obd0iII7VavnseGAvjoLhn+nCPeEHvHK4O7UiWBLk
qoz3g17AMJYiQpLRZAQNKyY4WiGPjmQ1fbzPyu0pQRtYk04uWkgBReNQvWuFR1hH
2rhBkYUt34XOuGlS0yAo+3pP27x9s62PrMgxdpgrZp361LMSasT2GD6Pwq7bHmuy
wjyHH3EF3BNo/SGolruU90QkkICFC2qGGmykW1k7zmNYLprhqHmd7e+7eX5ac5M3
AQPPhz3L5W+YrnxMRGl5IRQbAz39y7tfmsTmZcKA9314tc41uGTFqdR4ZmBcV2eJ
7/nZ486k1VABBZa5J1nCNI0/KutC8RFVXYDF0T736h/p9aRlQVZ+h9AMcLSpDwMO
E5HaICysz7ypIODOa8cQUvpHYDd2ad+0yb+YJtkMVh9b4GxS4TmvKG1g80Q3d90U
eOnyAjlmoU4/Rj0kK9QuvQ3/Ed3PzxEGByFkFfiKj+tCx178WKIWM57cf1PYpQ46
egPe1WML3RXjMQo1Si0+TDkrT/YvZYose/Ny5zwCBhC1IJrUp0kLgXocFFXMCQvC
aAEUlURemTGq1JIrbv7xJqDRE5ZCmHGHRB5/yX0ehx7S2mOnDRN8JLi1XKCtkLaZ
fftk8pl2FDeVyIA02pOVkYETLll8BKoCQSFfb/4JPZpyQOGNAtF+YazfnQRJ445v
k0xQM6udo9L0W5Pj6ovr3+1NUUL3GCYFxN8pvKkRO9C6aaH0JNqYK5jdme0FS9sC
pAx4zKk442Xdt2/loLEEyZLMzSA11DJv0Uhcce7h6em7RaaUR5NqKOZ2ZYDH2BZL
0nKvUYzz46JAUkU1K2xUT9f0potoaz1QGP5zhNItLpsXRXijUwImklY8N1BrpdGL
6A5gsSSRc/LNt/aCU7iSnStQYDxr44OvPWNi1Q63HaBmsGb36dse8lRO3Tv7YSDS
YzPW/aStCuwT7BxZR6jDQFVveA0ET5QcHaIuw84YEoiz9gsCCGRQcneKrIIDqhXl
HfXfLYKP+LfpccpWWdBfqG5ltPwvooDLE71ecmB8hfR5VElu3ayMdOKqNR/kHb6O
UP9QBgcFL4PuRrHEz9lcEzNRzCOW4MF2KaOs87DBWnncuDAFNUVWxbseio9oP1/T
DsBdqEjCbu/YrpYj6JkRnYgME+8WnIcOLm4nexQ0069OaZuNMehCtatg8kA+ByWc
oB19FlGTNPf56oLFySHwYiDUFLebhwZhIpQpYloKVW/73vEHPXPXF17OSZ6pYpHj
cRRQnUkwXU7Xo8Z8ynbu6Aej8QyEZdwhDG8+oU5YAK5ZfGMJdavtxy6qxF4UF90M
LFEgt5AH6XZ48FtIvlyUB5ILEsKgTkS9hf+ArT1na+XbqQKkQa1D6koef8+43zp4
L04c5zlsdWIzqyZLE7AZT9qYHZJ+mQ6mI4CyyK6f2YFUQrh2Q7rD3UePP1UVkc/q
SrL0dU/nHydQ9NfZVGncrR2Jo8RVAiAJTyEj+ngtC3kP2bNbQa35KOkTFgSpoj0C
ob1fjqnHcfhIynBANhhS8wR41VSoYtFHq+mfel1iiomlAbwcO7PUoP89+Uas3Dun
mGgeqNptSOKMHpbOwqT06irol6TNKZEURyKbz8MYOCTEEMKb2P/o2PNyOVP7Bd0c
ayiKi4iiy8JL8dBlx+WcO+0++ig5J/9AU+Au9vmjl76pbcRuNMF1nSQUYAcZ4CMO
fU9THXDluBjGMrDLmQKy6xewEbR/TCPgjzPZ63tt9bI0UDDa5hFhZEvtUv3lpyj3
tpqTJG4MeTuwPhVFbUkTJadN1D3OFe8ciJ/JNLVLoyxMDtuAtY4X7aP3QPuu7CRe
f4cW8oaouJtipXkeWQipEoddW3X6BldE+2zaW2+DE4jjuXne3zVJ52bwK0hSmVa4
1wwFQekORnZOY2UNtNkQJJ8cjWNHxNnqEG1UwvH+bY3nLSUKYbewkDxfYjxazKdL
Stbxwxmbj3Lp46KG6TGoIauPLclqdP8tweSqq6b47xGnQopHHdzH6ullzLxt7rGb
5nJ2P8ZvlNRl5dtAyWWNTbCR+cuYvmfh5aHg+6rssWrxq39so+PyZ/vRBcH10lXK
gTq/F8ujEQu7uGuys/w7Btrs4JwlZW0QanqzOolC3w5tXVAGJU4W7KjHBSJjjGxP
smdFu4ZQ0FGuOjy1XwhkfBWotgzIbBeV82JTFeaghnZzr7IVEJdL/8Mn1P0b2aQ+
TEBiarUiLUqx1Hc8q5DH4LFR3BlNGz2d++E2EnF7gKRxZgLQj0T0gvMbNU5jHR+6
PCkAhYgUcO+JS9REmlr5lmu3RxALpfTE/8hh5hBsZEYMtKF+CYPhRu1LOI3IT8HQ
+HXwFyZ3icbf1bgPFftrVluv7rv867DZjMOxilPAlOwRhss/5/pDRcxdBqSyceNV
PIyaFz6RB2pYQFTYqLiHw81JCuza1uT0pD9U1JcE0e5CH/VJYNl+8z74p/EL8sqF
/y1hloMxwCpEHZC7o5yEtcZ+2e9e8Lu9Q2YPXS5ix4O+1uQa4bjYD5r17nCFPd+2
+nn+3PbCI2fLGE1YLPiYtqCMiPsxHUMVoBZbv+RhNl3WaW10BPe8pK4niXT1ZmeV
mYMa5XUJHwtxNsbtSMOXaKxo0GgM9y7ura7qB6ls/v8B3gRjzbazMYjkYUF1p84t
SuffAnDovduBgRNgZEZYFXftZpRAtPOmX7DdIZhXqWX7uSlJJb5zhp9VTzurK+XS
wZZjpXKHkxkdsGEDwSuspgE+2tkHFHuXV4mnfX/EM/HD/8brpZUbPBDEjvgU0ZMu
DeUYHxbMrepNv++ppycif9fkgUr7rr/nEhlXxF9y1k/cvMoFrLsQhgOLnXsKjZFt
P+4/eJIvk5sBAQ8/So0wVsL7CVsM7Il3gPT4qTcn34UWhkcVSdTGtT/eP5ve4Xex
LsqcnKumMXpBfWIam5gMrr+f4i6WLLkQlLnZ1EAEu242jhotWQnQ0egBaGgiZf2h
F/eKYf+MazsZMx725fWJJzD1MF25/5fAw1H7tg163T2y3kklDSfwzDvGgR0eFccA
H6KQkTqRC4xlOZcI/WKkS28eh4hzY95dHdlNclynPX9LFN/ntJwCoaThNvr/gM68
oYwuhtFQwxHIryGS0ai0oS/ZiwW3k6HYTyVvKi/auHZYLo8ajaBHOwZbxnY8shAh
wBHVILeZY7MTu8AGC7aOlViByNtpli7oX2VYinER+8Cv5OIaZfkP7x9haumm6jKp
nMp2tAD0oLksy7slYMDo+6mIyWxNJrqHSBdOjMEGEVrBxL6Sg8XmByYUxploZXoF
6NeyHzK//IlMyJQxPdrP6N4zOXQVNv+93zOC5OD4Eus7Pl2SFqe1BXpbsqza58sK
UGH5qP9mBIzGd+GOV4NRXzvxKZJaQ3XixCa7VZDdNgmVutYe8fEi8SBfWBoqB7t5
fw8TfK8CVTkDWuMH+Ykkd0NECiGeOvtoDxNZqtqzeuuKoEeqNEVo3uv2hGBotfch
c1P3UgBkFXYZeOnTtx6j6TftVAH4Tc56g3l2vNtlvXD1HurRPeXJooxuLbmOrYob
at7LwyH4QMIpiaoFreAkoenQ+m0oQMw0SunvXdMh0EtAlk4S1djCVCeJgtLGDA7d
qSqAVXAY/ZjEwZhH/p5a+v2g6jWpTGtNXT30zDQyjWTuTvXa8/e3gegvERrfbUjy
S2XydidkhC0VCByM8eUzOl1Txai+zgGq36WOmF9QHufrWeK0HuyP9jHZ3yzYwiyg
RoOPcGCCYiAlRPtEDytDTFTPA51cnjQmML/XRw+KLmNksd4DFSyT/um1r6iPHCGH
c486Dbl41uAF3gXW7yugOUAobdt/Gq9EbCzq1RM2YXkzV2eG5GGgDeGorgBny2kU
TjpdI+f8YR9gZM5od+M91DhRGmeFNGeFzgIxPMdLq8zaLf5K4g0lk+FMuxLJYJLz
57etwfoPMFdwr/df3Txokjx5zSAOpvdiMQV7j0enerZ96iaKN5Anycc5ydchLY6d
k1mTHlTv5pA97EG1q7uL/4Kd+V/z6WjuKNAU9c0B1jmdRBMAbukafnc/qKe8+gTA
hlNpvrHaYFZi5hgkr0VJAIea12JIOk+xxRH+TDo9iF6g1Q7p/z9zzBWlKqG2PyqZ
xhsKYn9f6EvHFqcSCX3BX541wvJXYsOi+mPjSjo4CchoxZxFstD0dnoOAAI6hr75
YNGBs7EYnsfMZlosWVeA2m5+wK8q9Akn+TLewjyNOGns8z8ok9QnsNSyZJClcLJM
L7HWkHELJSC5lGSKanOOFBCvpYvcTSOjYtRkteW2sEV2JFn3O3+l4Ij49GrexJmM
x44gl6aKOsl5BRM92NUbwOEn0YTq6DuKILEt5/QYRozbyVgeLGd6t1/iAhbrLgdR
aBzjUoVgHTbKOF0D1Vkjzz2VMDl8PE2glPLera4mw+9+ExdBaxls9E45sBF63buZ
rbL/z62Xo/E32Belj2befaZSyESMmgn7q+EQRYJq/olV0fAfjIFjd+AQDxbOMXXu
nA4QcIp33kMbkAyN4UZuGOrx7qLlOoPif6qv/tCoMkQ7iseqTkTdt02bwyxQMNd3
iXwCM6R7bjwwgBqDzSCJrN7ieMqw9LPPsyGBq4UFzBt4EkIDWj4BbBxUHfiiz28i
xMZGGapT35jgTPk/GuvBoewEEYxiGSbWxUV9xLHwdB03Q+tKEe4qzzMVqXoTUfwH
q18qiHsrqW4ZcXOciixP+iTYR9gtJ/6HeCzw5gHjhpNDMc5Qr5TNWHxWfM6h2EJ4
xy6Xm1u0LEWCiQ2iCJD0K4qo56jfph7W7ka3JvY8CfLhcuZzhePXsRr4mwMDWCUM
oONYu1HuIrhDns6YBZ4FxF6cumcT2TFOvZE7Grm7h3FTISOWyr/dFWM4FzPdJGvl
rvP+W8LeVzLXXRNDF3zOSex5Ym3waM4ukPYPlrgdFSfFU2wtHiWMZG5FRdAbAfLb
4CbDVgPQR914/PInOeyNBWn5V9EMrMx0voHblUpeRgMStvxXCQz+269z/DvkFDeW
indJIbNPggtHzLUyxZbepORVPt2WBIEo9bWBiRMNk37SOfME/uYVJRp932mMZQNe
dVzTJcUjZs3tYeSP+ajyE7fV3aI2P5d+fPVwx+rA1UVOQB8owmfJPNYtqk9XKyq1
kmWU6jC5rV2KxKrtLXGWc0hiVilyAM+czkcwHyBurQDskDhCZb5s1JjQqAXcnLW+
9laQLR0FedQLOIWslar4q3f9l34d82SDm+qCFua83Jrb71HvUxFvmEDQSL6RJpQL
anHMkn/VerNHvUb9MXGpTV43Ukf6ECfnSIPGJItv1QIRNKtdcMadOffZ+FcPPyXz
qfYx5832+K3z5nvBxIW+Nt4EZQh5/CzpZuGHa/JOEiYFDKZO4hwRUxATOAmQNw8K
xxw9Bu5MJtM7yiPajAI/XSjV+hcbZ6oV/b36y0P31fB5FTs86Bj6pTJHRIpT3IHv
PskNZwYZM/uN76XFDaA6HI52udaecgK3RZKgzK5HSjOvUcnEwVgobATIDKmTqdYU
YrwGT5OS0LmGo1vZS8U5tk1CMiuoqtuW29ypc+TjvkuDSSLMgFcnZ/KsunnTzJAg
jzHZXVJ8XNsx6r6SS8MwzzAii8IDl5iR3xMowMaPbnw6xe8vR+pvTbYFLtIUAhG/
HpL/X8SeJwic3RA78Zdcnbor7T+i9JxDYz4ruS2Kpw2wHgz11eQodi6V3YQMdWIz
MaXh/rVntqRyZ7X4OHRRV0t8xd7AsrbSgaluHYBdRQL3oIwJPFvPLgLIMBPgwA5j
Joy0uDa9DU0HqzxT6RWrtldl5MUwVlhnFNApgu9qUsED1n9JOxaBSYtgpFgYWT7J
J1yLx/unICkxwpaElkTPw60ITixP4aBs8FTo1eWRC0b+zUc7DiqX9Q2WyWf2RIUx
4L3u4I4C9tF3kI9xWNFh6XjCCHmKoKf2Fi9kNKOKAJZIxuyzj6sQH5blhl2JyD1f
12skDFof6vYJRujv+ecWtHVr4TNHRU3o97iFAdIsQ2orQKRfOmlCtP0Fk07DC8pB
KbeBnO7zOMTT5GT6a1W7aMBJSTRaA4KrTeAhlBMxQPz5Atdv7l5CGACMgs09X9gV
ezkAegofxyhYxWEAD2pvVBknfsmHtfdw6+W82MZBkrXuGiv4PqnsWZmAKq4QuloO
V7O97+OdsZGr+zYvPj2Usd/0fz3mG6CThrYPPwvGLOU6168dHpuS6WZZXb1m3Vj4
YxDJwl4HnBbGKc+1iphakM0EbTORxeEvUbnyPPglTwFwe5pcEi+pv5uJcbvhu15O
TJuRtySJHFBjf4EFi2EjJsHsd5HNhaJk2lOHfm0HI1cIdgwbDgujQ4foW/fM22cr
jcyWClDji8SKleqGDZyWOy/pJjWnwRXL+Mkx3mgfA1DX2CGfN6ODS0da1/Ng4pyr
bvCimhFTRSWdxvWV6b1VK6Ghw4ktASupZ10hiawwvTlQuOhge6SJdESYiTq3bTZ5
pZUJtOK0FyjeQCRHsvvVxNEOGYSGaf2egOMIawCySf7h77jBBgZRdSl4BCOA9u8l
gNlQkoaIKq1qkrnG74qxmK81NIpjFvJ2nyq/1zRmWMpTrfYrzIBSs7QMCGWg4NB9
8RRG17K27Jjbr1+Zg5ta4A9aKoPinLWpWOdcauZtyX552o8z3y5cS0OcbPx2m+hY
0rjAf33bgdCwqwT8mtv+qt4PbShn5utCPToKYNrcysDAX1XPphvK28dlbs1y9sXm
cXM79xGHqk9/hJ4gIQzzbrc6LlHZ4WW/vPICeQTdLl2IobaEovLMwKbkCjxJY9u5
clPPgWWhWPJ6zM39rlOFfn3wbU8VDTjVymQKsD16Afv8N3lgpRaZGtw0kJofoTcu
PIotuP9WU/IxNbh7iUwDbNswOiV7/GEdjEFQJiIhX3EjgPO/wmMM9rhg8fMAYZFT
qoB/d245dOstr/PcYpIqkFLZBn7CcMPR7CM+I/DiCSQDmAFSxukZI8trmU32Vjpk
VrvJKd0b6cx/Nfvinvhx95ojyK9wBpZwzCy4MBx33bKyaRotF6JHicRCGtgmP/YG
Xu8Ipa/52tPze1uLF3ZXddHgG1+vZfVtbjEZ66ck8/m3gLJxaE7jHnp4tgjFNGMJ
maH4ogN6cMHbsKbRDWHFY+EIOCMhS1EMdWqEp7N42EtzKjbWTpe5gOccIwor+58q
mZuoL3C/JlGFQ9y0t4hH4uMmmzm+4iFls1wf8CA48/bJzWTpdYZTw46ELR1ZNHOi
rmaTr/kEGLGHJld9wibFfIdVz8Oaqmr58hV3gKekjQcAv9r6Dl52FYFVitMJVVWe
hWL3bBl2naBT4SGXl7mw03pJDTzny22XgZ/QgOn5jgHNHUySzy39tJt7QT8XsuT2
eNF+ghfkxElGT8ZSFHzzFXRLmAPHS6z+dWIpTkmaT0xSVhTJN2yyU4N2TWaYXst+
knnAB+CU9Hdp+rwJbXraZLCxgA9EoGcQBmIP5hCxfN/UcVP9l96Q7hNyQnXx721G
v97uSonwWxLdOsFybS0Y+kHk1LgdBKha9uKPz40bSPXMdwwa4fOhxIG/cL1ivldG
NxB4oEr2T77OxrqO4aVSbRB7f/y1gbxqvr/o/8SpjOeiEpqxtmSoeBI2tN+kEuO5
B4LHaR6qAjE6nv/6D7QPcj6U4Tobri+kMqJElTc//fc3GzBm1aoGcos1wR/ZkNNC
3DaET8VkiAzJP2UlazxYQE75kJ+2uv8hOsM0Sp3erYc8wCGloz9HfhFLR1F6A5B+
dr+fKtvUeNxC6eeELvOC6yjksV7s9zdvGJGOUHceAfbnd5ViaosuihxU+5Q7mTI8
ktUo1a1C2IM6zBne90HFT9hVMpBcWkIRiLygPBty1GCEE6t/4qZFnapTwNwqZ5lQ
6FzZO2dlRbI8+DvliFE671rwfguha7EFrmDIffqZjTzI28iiKfkkiG0bWJk7e5cV
Cqzu9vciUaCo6vICi8v+uSuLETzR3+CeOggbCyJTAgSJ/FfHWNogoKe6NjmKni6u
2hRM9/gMm60OyquYNmd1iSgmtD01OjU69h0nniAcLE/DN2r1oP9yVQMNm/h7I8Iy
IZOFwaguMVuq2CLvbuB8aGmODpC60nJTPdXb1ahvFY2VrrQqZAGxB7WLIcBqtXSN
+1PxkIrLsRPFM8dV83UffhKAq31zjrpmhzjqHmGNHgtu7Rr8ZocL5Rt4SRiCCqVV
dp7N3ErcjmllVOSkqiF05HUq6a+C1qUmlAKBg04lbGxPdLDrfzwmlgJXL1+fQ6q5
DfjpJb2NAQB8UhwmRUz3XIFdOhni7v02Zov4USjf7yXGLY3bjiDUETWMbhS35nt5
Nu7yhpzx0Rj/PI9sYbiwe13VaFBUcz9pKr25Ra0hbZ6njqS/7Xph7bccBqPmGHwN
leawGAT0mQIzSxnU0ZYWJ/xmVbgWOEg5BkZ20gONx8EehDVT26Q6TodMBLLW6SOb
P28PEquL2Oc2AhrfjKUKAnfYxeSexfSpEyIeOAKVUXr3wAx7/mIH6DO/kOxu4i3t
kU5IW6uz0kKdOrmhD5C+69yu9EHU3WgGHQZdyZBowmiPxJ291aWx4ZUrzCGFsucR
JdRuRiOsyut5HQ9XaC0xKmDSCP5VDgTwj5G/s2MfAvUXch28f8L7E9O06535ohi+
K56LCkRWKfBcEX2nMy+jxFLUfHY7VjXn+ofpSXGOZmU2suTfMNpt4PAtzdRsgDHq
3DA3s5R0KTdJIZlzsDMuU3/PSLeJcfMWyovC2RObnC+rPc9bTF0j64r8uUaNpfQR
Ki6KIYRpipSJm+Ef1DBU1Tmc1t9W6AacJexwcrzH4zfmvYbvM8mS+SKCE9jdSkoh
m8jL/xZVzSmHKxSVJiPDT4T8oawYQYUdCZoHt8ecNarI0dOPmFuklDfjBfIRP1HW
CgESKxnE15f7bsHdqE00uD2I9JGyj6F63BozuxlgOR70KxEPD/XZmQaADdx/pZz0
QJVEO4Q8kFfBbe/Mn+KYw1p3C4xMM7TnRD6DuELpoNgaRfYP+RuAjoIqW2VFBNg9
oAo0OxipMX+XQvMnUlcZUvNwus1ub7hyOZkCgmocDhDzkCz8qAcT8I+Blrs1j/PA
ypNWwJwxbqY4+rKtEk7aYT9Y+0apBV4qdNwrA44XdqbKkwDMSV78t4IsKAG020DJ
jnrJlMcOuUaIpMg+9Mig6XAPHAmYq2rbIfOI5W4DNdBXwvJR7u4CKa2uVP/mSB9O
HdPgUlqbNltCo5FycMjf5Ccf33ORnI+x5yxMs2IjkNHV+mIY1ETELWz1f4vdXRWi
qAEpOFM/FXKFGWvGQvhi2sqIqKiIn3fet73/XutTak0oAg7C49U67wjFRwRSkpc1
AK2Oi2mgnRIQPh3SBVSMVou+DzdCmJZhNL6OtbWhvTeSuTgyzH7xvU9al5It5KUU
bEFwpbgrTPD8t77YczYNU/np3vdWmCBphqM6d6TAhKd3YXPT3tgi/O5fn6lfRnlh
xwT13LkEuV6/ieDzlZCDJOoLtW7qyjyJE9X5E0UcWz8t4cUQlcZsqAg2/Kp4yjhW
TZxAQGwUoh0x5qP+DaSmzqboalKZRLmOrvLMxKeKO3mZ7V6FziV62P4cIt65QYHw
oukWTOQSCHRpqC5XI8bj6WyfJFb87EP5TNnWFJ1FdyzqnrWBAOQPcmNzn0UahM3+
7vU4irB5KyFSR9dcrne0CT0Rbvd3WWXDsbcZkBlVutTNh4epVldgC4UkHe15sbun
wN+L7mmhXxk7zFj0tRmwVlK5d2HfVd6Akh/1ZmZ/+fKQpCyLtthqhl7Cfpx4Fsg3
c9wCnmycKLOwOXSolrdKWMGfTVXuZDM7CU33X6YgFNoV3NO4HBzX7mCNG5nfKuH9
fBbcKSAluzeOJUX6lMx7NS+MULmQrzAq6pffOAcEQRNMWHRHKN59wqL96vJFR1Ww
SLtQZDsBqLzJ5iuVWjM9Ird0K5rkHGFhBHDQtmiGivrbT9qMIsTaWaBh7u0KXQsP
AXGLsJGivlB+cs8eNbP6b48cyMc16IhWK39p1OLPdNgrBDlDMcOlsQTV+uQm7wDD
/mxjFQ5L0B8Hi0LVhFZggOCzpUDDV+aPCQI2tUMySa/TxalwjRK4VCIlnn1O9ajg
lHMPLnpEENU47w7Y5G5J1fzbXSxJorUqq+Lh0y+fn1LEfbjmbX0qRRGWW/cV7En+
5JItxSlW8ckGj0HYkSpsxUQOZrIdsktI1aJ199N/2Nvvq5xieh+MFl+7ODPuPqFb
zAWleSJBUIMJryosb+L+mZ/mXYPBnElpJ8OxiJPyD9RQkAYWWUD5hgRxhsfIHCj4
us1t3P+wuDWAOIJjJ3F/Dt4M+k/tSwX00awf9DcnW2Rqn19P5/IlUCxrC+e9ueAT
YdgZM3jQB35WG+aMhcBndZaoeA1d4B/nOOgYKa1Dow4auSUmjGbgHHr+N5JHLiNc
a2GDU4jgQJXIClW1G/j0Nc+vx3qdtk45sizLlh09F/w2IW9l6/MRv3a8c1Uz9L5E
utA1zkQ5c72DkSjZmjDYd9HZ00hrQYQ33Ok17jiOTRlbDbJ2hsDQbyNPJDnZue9t
awkkI3Hq1gn+lOHLABntv6wq5B4FN+9YRKDaT0g99Q4HWwcJz8GUW/h6YwVp8pdl
+F5NXAP52QXrfSGjjLxzuJQ9uNTvsBFup9PFTavHzbL7ez1aR53E/buG3SFxgCca
zzzSc4OUdwVsS3qDjrXvh18OFLKmkrQWj4tmwlMUXDt7r7EeWWrKWs0uh5Ke4nIw
dv00xvsk1xyUj9eDgqPq9hiN/XKyIF8kk9DnP4kwBvemOHyfhUhPFLNoI8PiPJ38
zYw1sl5ecpAuEXCvC0UItc7eqj6b1wnNpRP5UecdY/X/9bFDoFcneN5rDRttllzG
rhTq/FZ75LWSo0KlyyZYXkJqCcQfu4NvmF2R3q6shBUfdDw+MWKUs8+9TZJ39v1U
0CHZOQgV39bL+qpc1m+VHvUD5eFumAiXpvOEHtXMYvykSFYUjeNwmBtd3pN8wkVZ
5/cY9jucVvWIxqRxYRWNevtZy47u7Nnp6jej2f0BDNSNLNfgUCgptcKIIFqaSRzM
qll8DZpjryb95D5y0Oc0zclluysiNRyjaIDBc00bthsmDA98hjm1CBK1BznIpXy+
Qhb7wOMqXR3S1SicOOMNopPEt7AT7JPZDq21PBiw327L1v9BrrQYG4G7XO+NeZL9
qzQle/QZ6zZLOAjnnMYWWceNomJH9CM6mBnWcPyAGCHZF6eGVC+y7DwdEMNdQjVV
oHqDUz8/9knHk2I7Gtn99423yDetn1V+RHx7zdeo1TyfC8yaN4+1yucfv15kWx4G
6mDw9rPpGKQjMVyMrgQ79qZbkLdkrv89J04yBDFxTYFW6DMo1rlsgExHSGKnAO8+
/4UN9McXsDofkTDaro/SDiyvFH5vAb+RIpX9fJWKIFWn89Yv9nwvuDOrHfAWN2y3
OkrKC5bZRkpoUYbHKqCCu2CxCVowIETuJH+WVrHzDtSsWLQEd8noxTjjazQnBc4i
8KbxFpwEfEVWCBATukDRknFaa3dex5SmKJbRvh0x9cc/e4SGp6esV+6CmFgvXMr8
K7sVXuby1bpY7JeCWNOT7NqBK/FibfeKwQ71UyTTNuCTHgyztQsEaK6GLIgrB2na
ip5m1HIQxyctJTwkbWv/rRgRPtwtjyE7XWc0UXN+IadRZaxAvNtEFmTHIJK3zc/E
9UasNDR8nZHbcyXfR+Q+hoAjU4yQzR9OUvlY14elRwZYYTcQhpTRijjWFaY2eHzS
qQB7wnJJO+BLA+zar7gN7rbILXS1z+dgwzUvOVG8CBhmhpqvCcIgSmqt/ZsWgGPR
U1RARZFYdY32rU2UCoCi70iohFYHHuaam5VZ6SguaKkqUKmQuXAR7vAf9slAl7+6
RG1E9pHNg0NebvEqsq8GlkmS4FUMMZrTM1V1kLol0sg2kA+w8pIvN1LjaFAkeuPt
5EqtP5pnRUUnZQjjJFpVVglxKUyd4smXzfaDXKRRvSgnYiqM6zgLDWIBJUno1jrj
RnQcL5raPpqozQe9foQm4i8T9aX1NsQzxTpRxXSz3iKocDOqi2w9Qd//d8iuidyr
vlEcu2WuvvITd0O/S1bQmCILpg7l/4VyJOfv7dCOHKlaaiSzlVRa0yWkuj/W8PfG
dZj9bjEkbuGHdKYV6Bf1bai3jwFwJB2kiYosOlrh9N/ZJiS64TzBXPM1z7G8q1mZ
O/yBEfg0tVKT4ATZ/a7OEOGqEkchJhdROxauzbySUaDyO7+zXFTpXVniX2drvKMu
B/sSM36e4FoUYMQktCuv5GeBlrj+Su+M3xj6Nph1YH+o3jolCXJrTknO4hjt1CTk
FqsK506trFQ+nEREryoyHfKF/p0dprrKA6vKdve80ZIh1etwP1RFv+bJAFJa0Rkp
BXnt8LHK8tSm7r3y0L1mA9TTtkLQhIefgZOut78ikxBrT15Iy3r7o0KY49YH9UF4
WRHS7Y2Z70CyFOsNmkORp/HsxxAjh/lpGwQi4+I8LpeN7K1VP0zg1DoJh4JMbTho
VUlXgDSLJtnjtaer7jHjPG6/ejXA5k7PEnwHq2oD3vSlGO8WBrgJ6MfPIgBGt9YW
g2E/PlqU3DDuAw8q6SCNZYsDeTHuRspwIQu8tnB5SdT8ZK+zNDPmeGIYiHd+sf81
4R9YC9HBSpWKO5M7VDQ68mxW8X8DNsMvIsjLZKeGMYxk2pJhU8S09/WXKIU5zdv3
h8XPLWU98ha54iFwOS6MShvWx1t+edrRkaUTVWdJqwaIUJmpT9JIU1RnESDiGl1T
wzaYOZZe8wZs42wiYp/dXvQfjOUlNc14ZPkZAhlLqS3w1VunbHxWHhW2EBIa47nh
IeyHX+Mrf6IKQLZAf1/mLYdNzx/N1aRfwQ2aPyNLxfju+n10dh+ML6oKQVNjeRX7
c7Ajo/f5fv4jg9fyYFGTXEqT7AfWBDt8BH108YxnJ2kudO2Jmf3faZyhIRnZiqfv
ob0/3yRMSLGIUE6wxRqs4cV9faSIiv5zebHiMOStdE31F+j0Ki71NMIBuh48P8qp
42Z+bCn1Bpzd38ETfeWPJ3eh4duZzf/zsOkDFan4MPAGR58hh1WMgXz6xmZLIEeU
3JxVhWualwFVauvLF7uV66YiVsuLTgGQoIuYIpEpHLviZhZL8XmJSw0+R655X3CM
jEWXz62AC0zZ0pK903ONAnYv9tZ/8NW0YULfS1G2qNlyPJc3IsHFjz//kNQrKvsQ
WoqdhXmLFDX19vaWzUGC2JZAZG+ppm6GcYnz0pEM+z7t0q6qX09eYj/lw3sdvtAx
LllqUo4jJ794bAaIMcufzsc4fC6oZrdQAS3gK6BXhxEYOWstqcnCNl5BGZ4TmDj/
CueQlj1NDGVDJdKP+ODX5FfqbEzVTLJvxeMFBpVSGWxQJC0L1vV4iMhg0hS5PVbA
lwjRwEPgfytxYLX6aI10BWpoTZNEc6SKthGUVmeDqthkSkrGfspHgtNI2cn2Ywig
sJiS4LGNl6s4It6nSOXorpLAb/dk8S3GXrnt7wCIi7xVbEhXP6jzL2ARNp8c3lL7
WRfQw2HLsqZDWtwADThV0qQLPohhz6Ay5CAjAncwfPh9WSnlAR9vOTqBPqXOmXKf
YBDSgEPjqQaDKVhkxiQGs1zyIDKbnCzsDKbtNoSRlBTEOQ9R/Ys/nwXuQVoA8bdq
mLNh7Hqho+oSXi3CQKZSmlzmBStf2DcJOzo9y05sS75t/ZhzcFI/b+O9v66aiB74
Yx8wlJ/Nbz5iP3EKHfwJgdDCBBrpO1SWbz/ouHRpZqpf/XYuQ8AmSeiP7kjo8RI3
RaOY31V2gb7jc4qW3Cuu0ZxjouDPykBaNBqfO98V4t1tsGrsXxI5p5KxTluigEg8
UikiGq5Sq9nzjaQyzAH78WIL4Txg1s/BMkj/NL5ZlPvnUWauqRbJdpq1lAtVDGiU
HkIX09+Z9v6PAblzCuPWtjcVv6SmzqzCjhTW7BmuVr3BZMw5w9fkXNnz93A1Mmvb
Vd3O8TVyo5z5zNP86c7lAR4+JqSn6aBdJIsWWrd7X/bzRKMM8sFDIa4Lnnq1HQLE
8pWDS2Hp9yhezzUx7zW2leoRiUjviaZkAy6SEo1g8C4k5uKIVZdnLSZfCH0h3Nfj
a9WJCVCtsOA2ZuisMOzaHWcReDCB9bf6no9jaIq0Rr1WdysoHZHZ7Z1MDEKNxGDv
3CTjZr7I9u3cDMC0Zx1VqBxqEHeXHXjOEcJdAemlUA/XSn30fL/HI05cxKOk53wL
WtC/TkSHyPeYGoITpu9+HwB1JIb3P0Jutr1+OW2ovjA9ihCgT0gq/MIQNqhAe1qM
HATCbcAUd2cwmgyWDA/XnaECIgOsgsMAvlH+C0B9UW2DarzTIDMlC465xoshfHgD
Hs0rBNDkl2petBchshN74HfbfR0bspvKCNLB3Z1YmD7lxfNNFt8Au+OGMBV8UZ5O
cnl3aW/vx6jyg7MGTZyTMWJEO8LK5VZi2hUjnHBaVUwxle91F92pjL0h8y3Gcuvl
klFd28QqcF2UmdW4dGIWKFTbPDeR8Pz2lYZIoOB2rcVj8wTmXcIHmx+O+qzOQmY+
PVH7PZjia8i2Sf46MWxncJXrLlenDMdhz+bb/pWW2n5J1NMykQoU+PWgd8ox2UQl
Pwx9opZyBifP8M8xA9Z57GMsSNU69wI3Sf1E3nUCh7GLwcCfmj65Fd/FbG5u+WcP
VxpbyNM0dF6dbtfBLuJl/59ST9O2PIPoKMNtFlQFJB6wazU6sN1v8iS2dJJ+EEKp
ycTe+FW65CJ+hEZ8GWE6HS904OkxgD3Z6SgNntaDrIN+B7y+ZiMfR1T3xG8tTUgB
iXff3YmCT7hOKjmhhFmkDT1+KcpeCP3U+EeWfg2jiJRUbLXmqgLIID1qjPo+3sDS
tx+FTeLdnsSgL71cKbmidJphz+KB19Lx8D0xcI5+xSt+M9pqw9irl13/cM3URwU5
I1+2apZiWB9S1Mw3nMf1WXclcpnBVNm1Ur1voMm5pdPwwkL5Zre0cMh9KKJBCOwO
nQaugPRESFMSMv5N/qRGrYzvFv8rISId0Ze9hYZ1nDZ8cPLxRcB1OVKKXvTFbrA8
idv1GHWjespe2A/6Xb05/NDRbouEaNG0tGh2oB3i0gO65nVYXP8nepiZUoJS55wd
RpPIzu8+M8lWj2z5arfzu72E+n+/U3qdfddXfMVhsU8vNB17wq8gkIY6Nh1vXmG2
nLk5kZSZAFoNWlyYUAz0MY9rLUUYxyKOxt3eB7aB04o7PxTrT1Bm4GiJ+DgB3Z2+
2XqChbTuMu6uivAYj3uHh/ztKwqvCtTPwKGiwOWKYYovLbIiGfxyhbT5d1yrbZIT
Z7EmF7cwz2v23DJZnp95DmmrG/R0NcUDjF06w/kjPivU+wY4GLAJCvhjJdKbJkuS
sB27z9QvzhQ6wffHxq391SKzl0RJqlCGALLnjBhPR1qMYF2xe9DrGhYBAbkfuXe9
/vSPr3HQWhWnlc5bSGV6lzP9OlJn2RUixcW95ZMMLnOpnH5Y88QU7R4I3oVt7FYd
5wBlklESi5Bwa3O4i2fxnZWD3GFmzQOrSs92bLOMApWQx3VN+d3vf8pkRfhI1xlq
UMdS1SH5sLxUiQ/p0ldFcvlvWjIE+l944KH+6kw30DOGB6m5od/2V7tzU+BjWX+7
ANVI1ojz6HEDdQJqoT4dtK8QXI+Uj31w7dN1rdMOWorbH5oFxY/g7pnPdU+e/NcJ
0nFASJVD63jOAbrwShnN4L2bJZrgGs37er7XwryT2qXC3kFu6Li6oIRh1pc0o7ls
Bmvay6i1ItLkBjrnP/Gkw6LZtBDyGgzAGhL4BmQ1lfGfH+E77HkilfgPEmyFLR1g
RqNuL6jwuUp49UGfMyTBr9SQ9ywPjbtPtsj4OwHbSf7Cy2zig/ckKy4x6PA16lKI
twcEtHIU1rIHoX9zZOzPyEtLzmIbKUNivrLxuGNsswENl5lO2iFLh4a1xlGxpUUh
EhC2PyO4rfUo0c8PPYIWbaU8by6fqlZeC2yn8AhOxQN+k5QUf44tHXQvIJOE8TaV
LJIvChh3NAatCFZEEBakfjTgXPAlDaaxQjhjy6Y5iaxAjuTpIo3gSgnqcqr1PipX
RHJmj+ecUgsgWqo1obeiBT2I75wAISama3m0RGUHN/fEq8wqk+fo/lTJQPIXQi/b
muVS3HDLwXb1VPw3sCJSa0v5ChasKqHB9sj+htmw55sk47FA15Uum435KIdOGYLm
x40v/u9es14CpjIfhGRelCoUZvl3RdpQlTdQ1AyKiILPNtnLpo1N4nj4ecNfIokO
ZgZs9d0WJPHUhTJbDXHywX4R6AHXeHZLtjt4qcqGHE4/JuSYuDLyl0JJmc7TbpV1
ri3fIffJsRZSLScyw0Gn0qDkOvBSUFReD9MyHJpvy6myH6KKnSc1/ZP+B5Wm4CB6
H+XslELglhA6JwXAjG9m7+By+HYoavU9z5r5axtplenPKuynJG0IPvNGCb45pRKW
ceglkq1zlFOpu/YHM1RgehGQZQHPjVLc0lidTyCSa32OSSoliS97WavRZKFaRmEH
6rzDSgUufqGcFk4r4IqVY8anlUARGwkAiqD8rg1n4DP/IEmgdBGxDF+nIbo4O862
CkHNOrf72aFcWpiO921OFmwdSNt1o3SCkgquUTGLEtb3bDdlF93mZJCUVnXJ4BdW
xF/zSku14cTI4kf5v0W2p8mb3J91skYzXeAKig4h3M8IakEkkRJ/DvoiT2wuXXts
EDMoPhuhlSSndnun1YUt9Z71oDNwfhTooIDySgC/IMb19uyIfxQ5JbOsHi5JcgO5
gU7wkcB9f0dzfxQuNc5bnaM1cJMgmgrpcsTgLIY3TJ6pvII5chWWTt4AmYxQUy25
OPLuJlwCnXKVzHX7dT6Pk3O8X1cnQyR6eFE9LRf+r9XawSuJC/hmKDj3rJjY29b4
bijr7OodXeCNh6VltQAuUrnow2ebMMgeUtWy5yLWZ9JYwY/cQqnN7BKZz2vfWpbn
neAQVZ+7oRWHWjBjk5aVdVozKiJsPqgEbjzMJI88jGxcCW2k3QEzS6/zOMTc07k/
5QNs1GCVt/rvT1Hbjx0dNyrg9Ot/WCUE9xVbuyngjAn/E9tsn166bS+whgAFnLnS
Ttu8MGdvmAvnaogUJRy1nHEyL01aiMtioGZKQptLQJidjcQvrRKdMxpP5H4X6NhR
TaRvSmUE71Gftzpd1M/T7yAbC3qLUFKsBY9ByAnKle/fktjIRRw89/HihR7trA66
n7/siK7ACw6lFa8xtw6jOZwX1GEMXvQU/+GqzXuXJ3OGN/CacbQ5ZmNvP6aJv/q/
fvDaWijvm7rLmVOKoSJf2TB2zB1qL93/5GPmOxvFqBZEohPSPRifH7AtqN90UNlz
b1i2trccw/9+abMK6Hd4TR7nP0eHp4XTr6Oaf9EXzxzosGES2K50jo0v2uKu94U0
xzlJB0Rkm7DOCxTtj9UxQ9cOaE3+8l8NbEtXg1X2WRv7BFjNSZFe5WOzysyBqswt
SDGWB+/pYYhxc/G95htw5/ows6rXbwFIYew2y94jul3XFKAf0PavhjIsuT1tSWS9
lw6CjP0XpE81bakEfJLC6aCVBR+LHOuYNyJmF69yBZCieiOvMkFBkQMXERTGFwR8
9nVgT9yGjWhTuS0+JG7bSnOAaCCqq0miPzGUf2kY2k+n7mQ+/j6GGijwfaUXDHYu
XdwD+lPF+gfDJYDgqWXJFtxWbhQshSInRZBVuK+aWJJlYmEK97GMkUdBZKR2FEas
1/3+knztu67m86DX94FLyrYzwycd7kWz36X4IPBQWH3uySOLsK5ML8f1aUUt5H3S
mbmwJqPbRGaDz8Dc9m3uZlKFRw7Ay/A8IhxLrCxs55sSxCXBpWH/IrwVvfKWl2yo
9GZMXAJgJck8YTgff88top3unjHy2m5Ob1S71F5gWee3EhUU5hITcHo9KFGW48AO
wRDUw4eW+tDfz6jDLOTPCGNoYwB4IKuGS/GEBKUz0IZxMmsSaYeGQu2FRmEhlCg0
+rY63hDbhNcaQD/Tpjqone2WuH2yxOlNNUYk+BqCEqHs9J+Zz1aP8WmGHpAA/7Ci
HVeXdxhjZqZbwtvOaxvcq+QWlkqg6IhDI3ucaZRoc8cNf8g6EO5UP8VCPRvOKgi3
JBddsF7A9NYb7fe/CqAAIeVTFnPv3sBr+W14KgUTavTmPHT2ZNYijUr4SFqW50d6
38crgjdE5Yxt11U+poWVCn6umSOHoRPzBZ1GJFFXRbL76W1GplRQYAUVKkvPSvUl
y/+CuUKkU4QG1teVQguV/Xa+EFcIKJTBA923fmygP+AOL0VbZebDCTaqm6qb67yP
jZ2fm/Um3iinsOAY0a67Lvvn3PNIppi7y8DqD6VAESb48ptoHaVpldtz16h36WYD
eOxD68hkNK7CC+7MB03p+Zo1jK0g01B98L9fmYb26YY91hS0JljqeNpbPzrmQKP/
4Fp9MRoRYBnQ/llm95Ri7uuunEOk1A5TsC5JJVxemlhdTWEYTq8CzB/cMzl7bztc
dFYxoOJcSNdzYT+Lzs+MJiBgraxHW0NmV7Tgh860hiZxkRM8/KoH+Q16VzNqzcja
Z14QICeaEXc2+hmL/w95Lv8Fck/4nudf/zQ9m238MkEuEvHlLwrZI4RYyZxeMnQK
WtsEVQHRgxHIAZjxda/PlKYFeOOrsokQ8698JOCHP6WRIG2XnFxdxRpR2qpDXBlt
TNF55mffIIZgwLkjx9jz0ozJYmwmuQVQSaLHEwDGRiy68xP5BIK1fNcz612AZQpo
AY7uVw4ZqpIdxnD2MqDPPFiKojkNmLbJNjde8x1PbSMbq+7HzmZKNKasfcfZa7wk
fl0HLb5XbNidBqkWi+EWza9vwmaaeW7LZhUzqm4hKoWD1jB86gxz0Kz4ikGZZm4Q
JfQYApIInmbNOpBnw9/3Ld1M+VLTmATpeTnHyDJT4UaF5+/YrPBSQ+j/29jB3Bvd
GXwZzXF0aFYOHjDMCm40vc2lIjoOQyVEFGtzs2mNxmCg/5cTWqIuevmkq8copSes
GlpwMm9Mm0NRpldR0vVsVtmuA3tG5iU2Kfk5wpVqAJW36W84150PPvZIfk+U+ie4
0+oWUmxFM6M6RMr99iNqVSq0hTRBbxv1hUq/eDwEWcK095a1XOa1BK1mPJeG0Ija
m3Qaux65JcmVigAHtLOsUwzBpMBfqR1WmEpwUdcuwexgAib3NtL/1rhvD+w7Mm3f
un+B5rq+FjAkxwPLjTthTKTsESzU1/1e4GccQzIoPFdUxli9knC0MZYTwjto3uZA
1nfMwY234cVZw4LTRkRoBu2TS+Ci/ukxKE+BYCKB2Xk/EvWi699fS1IyQR5EhnGm
hRJuAm1IZx5N7zhUmEQKFkqRUv+NLQVqz72hgnh3WL/G51r3s+9udgDLUkfXcAcZ
5q0WukrBaKJGKUcOWjV3p3Wb4ZWuvKIu08AsFeEE5cf1QbRe4kjlzgk8xyy8jlNq
L9YnRFyWjcAtzXoxcgqYoA9epVemQ1QCPlgb0uVLOUTHEjagxF12iKoceDOlf0Tt
dLzmluiztVbght6WpddCtnYT0zOXHxgl4grN9keR/70hsso+HiRCTGwE7Tr+LvaD
2RhL3f1vZ4qEa1PpbXVxZ5KC8LUIuj+2hzJeZ+s6xDbPX2gl3v3LwuowqLm64bUG
xxS4lKDXswZ0n3I9rRYBJUjCjq0dqMEtKs7yXm/Cs810f1WFz9jBx6U+z4zXbQns
8DkbIkktTCPE6lXYFJyu+KYIAoY/4cms95JXfcOSSNpA3r1v/WZ8KP93rQTRwFdx
4GhiXOJbmP8RHGnUoLOAfZ3ixiiHeTqqC5ZUzd7oP1CgDQjMPAh9A/4qyfs6lai9
M35sAuVQJfNOpuxtdDJJfbK12tcq/Cjgf7/X/wvH74ZNwRPS39knzEi0aIDNlele
OyZEve/35+jY4tZqE1ZaWDgzvwxQdlLtT0qJ5zKFEqMwu+t69HPw8F/mX0oJbi/X
tFuqoJtIWZ7rDE/EmjUy2MxnKy251cIVRJTYZfqmWZ6QjhQCdW/P95MTC+LpfwG0
R2afOKImF3HDhih7RFJZzIo7hs3WD3dJpmBNz3mN/ePDfhESySv17GcdOQrLsfYQ
NvwyN9BVumZ7ARaWFT+OLez3oBhlT3zakv4sMcrOhNJrylqCsRyHXdO/bZT27ubt
p077Oi4t1d106zSLMXglbdRTLzKxRF3DxdPLHY6f/x1Oy46zTh3GWY4Ao6oRHjFs
orz1I6UNryLgHVy7CXZ4axomk2CWewFuZ/PnEli4Mxhhr0wIZJzNL793wT7XQjdv
wZYv0rGngDVO1lyJqpAuGiJ2VRRVuYCaJtsclquFmn+nMBgZiMBT84X8+kuMBZCu
dg7R+jfNC+uFV1CmC2906xzaD+r0uRHe2fQZisoSiGKLNpvVtcdB1ybC/HiY5f9Q
yQDXUtKVYK5ly8JiJGv84rm7k9dsFUWMahMNwqbavLBj8vKnpuNvz6uDCX81viys
9yKtxfUZRJIqBEC0CgayYdVS9Q8jR5rTpzo5yjQuVJwxAx3V7DMLtEipbWq1cmXy
2lBwltM1MXm+I7EN0GEVVhDqgLHBJ+otwj8QtfR2pugLkDWtTlKB/eOjaY7voLgN
P871F1+OcJNT1fO3tpsWgZKe53aWMdu7oO+UI7ASfedsYB+o3xgPEjSgB2xYz6Vg
n9IVNetK/Ji2j7NTgazaqzMlvRb6/bR/LycA+WD8QUEuZPAyYPJEKIcTE/0h0+V6
78FuWpC1oDQ2ud/lOIDSQg3uQ/0jQw1NE0YpeDuaPIkPUrGHQqkliQkml/iBG/Ir
VNsJOLm0gJrN9kKWJq4PLvL5nUGJhCZ++6f/WL9XFNBC/wazLeaXamXz1tf5XAO9
RTEc9tocg97yptMnxkkQRzuvsRtSGHAm6BPrplP75iuH8H7E/QVl+LN/3e+995Pp
HEW0cZPZP1sskxflu4JGNW4ODFjUqfvR0VsfOcGom2EgqSe9uqWQUNWXmpw4gjEO
RnSHCXJMW7MnwO/0Q6xjGAJzKTQCTZd1Z2TzHKXPaG2i1AgwrZ+UF8lCkIMDrGZH
R/ynVxzTGYj29JBFbGRCtHAkRHyssvCCTgpdnqqkQR5LZ079K5XCh3Yws/U1rxSk
LREQmCthQwGsLL7qEQMsAqOzzhzOnEmiB3YVa/r2zqCwFVct4PSH0JCDf0bJnh+g
KryaBtKdO10lVk1b7I5uDwHZzE1RsvTNHtaSsCWWHXTtqV1I2rsiQToDhpaBFi+B
s574ZO2NK3ABqFKPsOtCcZkw1WTEvYrLboD+6B2lf/IbSzC9mtdo4bMoKT7lR6zt
VTy6wnL8zbxOLiRHhY6QEAwCd9v2aLFgV6nrS383ptsWxprUeBGZhabU0eP5MKZa
lf1doiVIvxCXhtKu8tHULk9Va/DQayPtOzA+SVz2uurr/zJXnCSO4Zc6n06hMSpA
fExXqGUPp40MYFL9FxoqgsSx4fx7cG9fIefQsXnHsVylyfvg/5VFrPlzDLCBLWWF
nMF2YoBucHKP/BMeduuHxMI3jvjhspYnZElES5BXNRiWYX0BxVjMs7hAe4kvM13w
H7RRxMuUt9ZSUTTOtiFTiQYsf/tev0bFydHD7PWCzZ47lmxkgOhQLb+HKB3RWAV2
toHQbOvzgGNCttXePGhzaRt/bqJgmcIJoBrM99xB8VxutqP97hKes87E3B+BMBET
5eo6YbjUDkM3i8MehfnEKMpfpWtUKIhxqs2Q64+Ho412X+EUKxjkJsy/rZuorpml
CIoxnupm8ysmeeaZHDSYRFIH5Cjm36i/x01iABfGJWMJ0LZyZk2Kx1XqMG/V5vg7
egeVoSe94qfNIeqj3rQppfl2dgbRPFD5wWdi5XMv7ozF5qvcV6CDKIHaHwHeShOu
Nc6MTNRH3gSZDpoT+vZwnHZyXVSjSv6r29Ltz4lgWlt8zgPkm7KliJiYp1A3y8BA
e5NKmqPDrrbpPtMOiuXsdiPZvfmq2Q4PMPPrW2BH9NaaGxhcVc3Jf8xyRXLiD/bl
ncERXiOT3M8mhI2gb2nKTemEdEwbiX+fIXKd8yo/Euw2ba6csF8DRaYY91jMTfrS
d9GUbw+Pk10Vs/P4a5FZ1OGVr1sjDNXpx/znTegHH9czqKmEiwA5Xq6YDVwhhJJn
ZSTyU2TPoSvx1C0Un9/vBDx01Zojv+tCYLrjPf0RvLhYJ0AlIkYOAle+JrqsDako
Uhgd5NRY6zf8HOjD2L9//gWQqlA3vpbQr7dYpQDFj/c+1EYReGnxkj50IaUR+DJp
z0CVjeTHOBpqpppM4BMtnFoBI1On/jjrwbGOGR9/vnDlhVS9vFZ1k8O7vt620VsB
a7BunxvSZuipfXxwiZAVqkt+VR5uxDU0/DXnnJRlAFnu0K15NL2cB1PqukimVeqx
hApL2HhZeMOYFepUJXl8RN5IOzp0YOqFLmkBEz8nFCZ3AXK8MlE6W2b42nLRvuSu
KO5GzBxi181kDWLpt1wf/DNGA/4e1sK9NLIiiQKZYUAv8ezL+UeMe9NRUk4N2i7X
BhbOtwICgnQ8600y9bcd4r1FoEQhCWwvqQYqc8e3pIp6riYMgDgWiM8+0SjTJ934
+2fyLp6yMtcgpErMw+U0CWtluPPtfI8znzXZ1PzHN3pIga+M2SkvGu5IvBSj6EJV
qaFQIC2IlQ5J0bCzn+G9pIsM2jqsjUvS+2SmU/e7ShpT3kkG2UIpIhyObGDsaRoz
ZZR+3zp9h62ai0d63RFRNpwnOzW81jgGxZ/Rn97bOqtL1TEGiSDftQD9MCmjQ4jq
LI+QduJmUJB0XhF6QgCmOHKiKxcDno3aA6X/qEAC4FZ16gVPQruNmlpAE+v4WLDv
iozzT1FG9CORextr7CYNI4xcRZgIutwIcKFPZiH0DJEHyP7MIM1kHEaRfdwePClL
TXyvjSRCyGLNWaAzFCUhJWNFqrKwMgzz8r1iCflCmx3d8j+HGoxxHXTljxyLTbTD
EbTMJ3lBA9oChTdMQw3vv+885GA7ebrx+jbMXOH5zJXRDQ1k4OrpcP9GntyUTaS8
Krs5/5DXkTjmpGdTk+LpxhiVuG17qWRJQGssf6cY3jJ+YWH9GRpeLMBvaeRw3ECy
NLWT2/6zs7Q6x4c8LqRbXJmrP/KH9LD5OOBI0RYxkuvF8k1tvgDixIxCHlUZOwBt
vtz8Us4v3P54fY//yAPv1vjAug5IkxAN+41J3KoHIltcNTNzCqk82YUW7vQWKY6N
hoyhCHO7zD3LWTE1u9pkVjGQ6Uo+Qg/MRV6Wp5CQHzT34osG4FU6RvVnLRI3hvxT
cm/rb3k4QpRzBGndg0KaAtC7U3ifibiFf8uUlf2gVJl1ZWJZAOWInIIAHgQdQoua
QvCt1aaOXrQwq7Tq8+QIr+b8vNzCM326PasEHmG/KAdFupCc06PI4ZiyZpGEt2dK
HNmerVygfUWVglHMDtOKgsApr4QCsRCP73e3gctXuWRldrAblDU6MIWeXZtwCmaX
GXQNXKPVuGMex8QXunFrmS7bhDIMpZ5sURePMtMDykWyoU8KTpgK3B6U9FOlEFnN
SY2AB07h/Dy46KkDtrII1y+tULyL/lscxGdrlYocR2PdIsUmXKsuYvFTLaLAUhpA
lKO0YRa5k/3Buhsevu2dyhYaJ+LqUxMuuFohBkDgSlfsaqx+Y+0XXW3eW5YuvSo1
hTOy8eOS2eogPn2LeQT8ivkcXaZVNzUDudbczECqm7pzPr/UPdjgOalksNs3hVMu
Q0yjxbh/L1QEUNTCB0SNT5jtat+M73r0HPr9CpYkHKanddrDgIP6As5cxAqiwUsY
5ncJf6WFviC3Yx7j4QFxLmaStZXOjGBFx9j1948WRHbWWWa91MrtQYhBYwk4eOas
UoOyUxTKnnNfn9GItm8e9hlBdik80ULMJ10G0uiAjpbEY3u1DNeKVmIfu5b4vS5O
ZWEReyHOiaNJoweid1HOV/DuP2Ekaus2VPFdB61HEe+NLMXjRQfv6tL8VewAGNF/
KXTms55eNTtDmLZXbNL++tfHEtCvGBY61bKWFi82NIA0hwCDxE4NZOZoyKGRJhds
c1VXXD8KDWDDV7C5NxczZSENAMTlkFVcKhZTH4m3DgRTRuHTUaQu8nxIJkPS+bHU
yxZsYyxWyZfcQhgha5PkOsqZEAji4Q7f+vr3Ud9Nbq1VPvA/eBldhWCLMNq8AKQh
NZz1VPdSJKckKjjjnTSm+PRl0n/VdGWTUcNBt5hFFScLJT/S+VJYTJAZ7b0Y8Z4y
sWnqw5cTw+uS+DGLHQZiFjb9hTc2dmeqFYF63ndgRpwucmlvpULGe02941DHcf3u
UkEp14zJrmCL5kkbIHZLjm2g3m1U8er7GVxI5u8EGP4v2AxpyLnU4gyrSVoBpQyC
zJr5YiZNHgJTFuWwfLaA88UTPRd6tX1yx7kV7T3i/9lIke+tThkL0qM7wAt9xBPG
Mjb1sYGPo7zduN/7eKp2B5yWfnv84rYsiT4TJXRn1Z2Iy+5TGVexmJs3Cpa9s22E
11PVhgDW4XJgFv5+2m2CtyYM4rqIRh4hSCFqoyZJ6pycdYdPB9sCS1W5lPgwkagl
YyqNAO8q54ekLTHlAlF7XvPTOJbR7kuoxFh/1EJzGncj5pMnKjpG9uK+driHSaIK
0upZs0QzS6dPijQItpi8Xv1Ra06RHy0WW23ETOgupV1+SjwItcAvxBq06LmK1u88
dSbmwSPmH491lzowo0YxqtOOqZ//YKIWD+1wefW1k/IhaBWOp9ect3voBl6lmF17
nsaq0RyOWlDJFcPTG5B65AeQN7w/H4C9Wv9IUUrkURstmDbv2jYLVqJI2pIh7oTi
8muSKCrx8yIYlSn5X4WedTx1o/U+Ftv2rDGUP8Ll3LFBXiPKCc+su4OLsXG5JEtl
oMVpuK+JGTvRobWacHjAerD/Qz37Hk7at7dchw8FcrbCkQKSWPT8Asp6AeFY+V2p
K4Tiv70kpdRcHrr+snx6aJubFFeurshdVKY3jtmEwjJKnNAaf14ouwkmLse5CBZ9
s99MFVRVs1xaa6KsSX0AQ4WbavX+6/0l1L3WgHV/qg+U3s0PlcWcGkEzrZkkFoAY
+kr1Mzc7uV47ZbbcgmUU2dC78gUdfRAfdv5OZ3Tcjs03GQN5GEpMxV/4pL+ncU0s
X1tkWDwLJTtZoSqwpNC9DRrb9XG1L3q4mQOzSb8unS2vJ1CldVhKOWLKRcONOsYt
O3EsVrvvgF4dTGx6IxtvoJbG0Z0OPMwrbkZ6KfdXMvR+XWjL/YEdi6Z+NAy+hm+H
F9RZy6V5Zxi+IiTBSfnyDepJDmibYFYQ4tlkuV0pFwWVJuWC2R9eJlPwn4i+o4Yc
X4DHzcsKfm6BIw3h8cxDuX1Y7uNA1QtlZJ6gxJgfyat67Ck+enH/TB6Aq2kWcDsl
bMlM7vO/5tbeAJIwvrVWWrB0BNNcYkyDevMEul17E3hVBGk59H1UP/tIYDUrtvjv
DJQCfpwM21jx7FA40H9oU7GO1ZGs2Z3Z0Y4JDKkrUyjjJrg3DP4cnn9f6Ub4Yu+E
0JFZVyiDezLNhOWXqR9y9WbOeRuk2eHnFjKDPJzTfLefGphm8YMdFC9mYeY50caM
Ae9v+xRZJQTiYMT+NQGAX7V9x1OGz0bEkTWrMLHDsbd4cTS2b8Xz2RJdJQhzg97M
3ahsPGGKDxgrIvhCmavzIswqwKR0rIUrDvjyYBq/4DGUVfjWRHzIgDNQfTduyLu6
+rjHfSd0FOnawwZmK9yh9jzatOepRRQPmqwHyoTMOfjOZAqB6esyVKo4n6pck11Z
Ulv2pJu3Gn8m5fJdH04kCGpW2SPp0y+Qc3owptWqsHtc5Y/9kbQ0mYbUEoIKVQeK
m/rOAQFKjysVPodIb9tTKYq50OeQXjb8IY3h5cydcdCXZvZ9QIxdm2/kxvf1evZg
a5/Zn/nJGYWSsL9bUOdggu8ZD3Rw/FvKsmTLG25ia7bn66FWw7Av9nGSLbZU5kL2
H/MDdLJ/TMMZOIzFrr+lt/06enaJxZRWMivPmRhvfOWXvx8mUO5AlpX3gV0vWJ9F
Tx6yZBt+BIfv0Qa8o3ecE62zso9+RxEjkejRoRqP9g+HlRBhTejVprHZRBdfvXy6
fyPFGph3FGinD8qEFvPBSjPeC0thKQLays3DG2v8Nw5P9wRP27LXas4ii/XgsPo+
5iNJfevuQb9rFk/sUH6invc8dKd+Uxe3Xt1sGaFV4RVrPJ+0Ipedqmp14Ux+O4dL
9MF8wen21+D7KRjhV7ijXjPCEKeRn7IQcPNlYhghLP3ObkGBWr7Oo+wInRk/U+hv
UOyGetNvukQ61nJQwWQyt/rJHC+ja/kCoJZs+Yqb9fL8InC8X9mz+ENpE8CLfYSB
2APQIIacRZKJQm8sGpuecv/gNgt16JeVRwzb5A2PV6kVXRe9mwSY/skcH83ll+W7
yt8KAExLEam4Eyi8cZ8YSxEHnfJKQqXq7DUu0dyZ6U8XC32yOKRkseqBhrLVliE5
/caEp17SWEm7j5lcWxZQFtGDWxvp9K6Vq7al6p3kOSNjp0d3gFHfzoCSL5cASunM
TT7yCM7UFtzVELmnb2199t90t3yPWPXeZSJzoRK8kX/0G1v6GGffGXg8BoV/GLkK
msZAutl3v+46RsbZDd7HlriiJiig0/KWMjSJPP8CJuiMfn/YaCPAfZQku+uX+tVZ
/2gjV0m7eH8vnaSyiznracce8bz5W+YZ0lyckwMrY7AsoiWn4WIjRQdNAPnPwy+6
VQ9GSGqQooMNk8kZjDcEheCUlFH9aoqIRNWlFrKV1AaO2Hh3UAoUEZr6JekckVon
r8skhuS4xkOtdTDm59kg45jV+ArHDov4IB6ZRmIvBauUpOXytsSjlItbTdEf9i0Q
fPhb8VMVa/JJE/2rtk1d+lKt9IEcOvQNqEoOuSdNdzdIlfHSqH4uH/lxr2IgjmUf
TBm6kkQqf1H/N29IUHlZ4+ET7wV8ZAoFuw7Trn380A2ceU31t6N9/QiHFLf1UtXC
cp/e20QlC3h4jgWTyqMc0wlsQ1MhWxBDUeXrpMtQiosPcfLPbw48oUiyX1zLX8tM
2643OBr1312hBCNmkNygCbTXKD8/VPU3S7K+nF5hLZ68/XbxSGVjaSANm04oY3Rf
mOP8K7hWqOtOBimyw6k38d9r8k6xAXdAbdkYVAg8H3bcShuWWCOWlY2Vkw6ITf3b
L6Cxha1PccqgUAKQhT6rskZdk+lsIvCrunLxRm387zJhI74BrpA39ff77WuQepwa
ycrLMeb8JX5WkegMMCYSUctMKtCmWjLIzOn96vPYi4ayMiYjq+DvK2u9y1WOPNbH
sY4+UlJIs1xwrmoba2YS+vxvdWhtXTM0kWXOSRODIA7IsqfhVXfHZqZHT1vyYHDW
aT9XRUdn+KYyD5PFt3CntoeGCQMhdkuuQ5y/PGBkXsZks25+NUDjQn26o+NMYQDS
bQs79xOTTi00tli+vOhssJmOb6HDpNsiu5ewm2diyQemzhImakS1bpiN5kbDMfGk
WbxwHT7+UV2HFz5VWtvmtJHD6qNkcs4gLcDbpdiWPIVMLmKnuaI3QPpIojb4dSHJ
0QovR/7gl9ZJe9d91xtJq4euN8wZKZzd1KkcNreLYeOojSXZO2TRun2RL6OZMEnG
3YefsQPcEaXBFuCfLm8go/wwai2ki4Vk/johzYMKhQbyfBtcWmh5aDdC2Zkwi4mC
VjhykHneMQ5SWgRu/k80J4Ga3No/+8qVIZqIO/pGS7q0jw9ZenK5ImAP3t5n3qJb
DxXroAA1cI5x63HbesbrjvCz+JLWv44XGw1Ktd1tbbr7DjjprzBmILYB56peHGJY
ZflnvoRVPGL93OKtBgvYnRLxfJwDSOV7npbcb97RGiSRUbobgzqxvHPujELcARNJ
iZ0wc5Ib/w/uvK0TSPkFWD18OrPa1fW8lmVkqNHloU/5gB7fMyndw95DVu21voYj
BkM6qTL73jMH3LoeGbuuz9v9Gg2ibBn3N7bjwt43fJqsN1W7RPofhmuESju/o9bm
SIYVJDSvxszY3PxtzLYvQB1jkCznCi5HEsYnc2Btv4ucmhxPvmWP8CzAPdWSAGeF
lpcsfoTSLSPv8sW3IE09WMYFPExZzRWW+I+Ivfe+ygL/L+X+V3WeE9UaU+JF9Res
YqFWTznR9QQIt+vUi4qMONIfRtqRPhmCj197v3dgBJ+X5S1ZTAYlCSU1byJJ+1WN
Kv/y1bx4+gzindmoXLl6GgJNpqgcyWKZD6DiSiChTVBM+Ui1hBiqFe53OAYT0MD0
JyT7P/hwiXMogOsvw2/ONoZREFDJEvgRevEDwS8ssDwcBZtdao0JZCJZohB4ULqe
sGUy2gXamXAuqaAvE7UpUxrQ6JKYOdelNu69pqbCvuGORgSRPdlCl/rb4YF1z2JR
lf0l+0fyA7zEfyPqgZsJzBSPeqVC2/AH/8aNfGnP3r6xIvvNC3T1xsV4e3D4moh6
LRGSPKcQVSZVoQBBz/iYr7hfebHEwRjFxGagJrfhJ2whPsjb000Zo6HurMiE2Xd4
pTvRYamI0sgWnYvwDcGvtgElnoJRLloue1cpV5fx/3gFjhXOEYtdDuQcRMKMBMu2
fqiEPw4rYx2R+CIR8StkjmhkcNywxtp9TcmKHkNaP7ot3TL4XpMlDzFr31aK9nR8
RldI79g9/lOkJWfoiE1675KP+FkBz7B4dKziXrm7owhHMJdFtDFsJwrmP+P46cqh
bMA4CxiyboqKblTlJRhh44XXqIZzhDtFFkHHpKjgryi3hbOldssMLT5im7Z6dbym
AjOQo3bkaZ/7OImdxO4jljRF6lwzj1LC+vzdQYdfbPfL0+n/1MCjI+yeuOea+0Oa
BEf7A5q1Mjf52lMjl6g7L90vq0lgjDNJ/ae50l/Ly3xJm1Kyf+XjKlvpH58qoAie
QAiaY+EqQOc5IOWqHvpGINTpF2l7rfg41RFPn0rYpWcExPlWEORix47jBRITrJc8
dbvtoSpV9wkyWVILlUJHYLCJ+O0fHYTzLA2J3j7mdQ/nrbSeTLSEeA1sY906H/mk
L+nRig63ErQsOHSXYJ3vK/rqpFn0CWJBZRT6Nmi13OukUmnsIkmwVDNcogXYRRF7
LiMVt5AQVpx+NWw7zjQ/maRGyQB/4nwPC3dWaqtoPz5um7vjwAhzJcGheKwIprBF
Kuuuoiyv77oSwaJQvCNa0rsw6yiAToD9oFQKP4axto/59ukPr5uh+DlS6ne2G1/I
QY+5zw5UHCYhaWqrXC5l7c0KAA7idKXblsHUPhvJE9iBQvXc/2WZnB8tnwCP3YJV
lMlksYOwYJo6nVrWHVRY5gN2qPdjiMmUOtUJjvwJqONIkI9tg/x3a3DGwMuFKyNT
OW64avIzz3VJDE2EiwN9o2kd7sjAMc0ZC/SjlWTAJ/Hzl9//oyy+KywEpBfvkpAk
/tSNlU4hgB7BbXqqC5JIeQf3Q1hIMKpvQ9tsgdbjduDT+cZmGauiqLkvzc0JYZju
cWKDMBMmqwtXYriWqB4rrrfQQGIOS17jtmgJIQ9KecMWzxQvizt53bR5SGWY5tc3
/nPX2tXcn7GGYmTpY4QwmKaXo0VgCPLi/t2B3CPm5RFgNSmI4HjStg1dyd42GroD
T8gaV6BwQ2TZGRUr9xjs5xqTWSvlgZdsQ66Ouj/5cltmRV333JnikuI7JmkC5lnm
zVlj3zqWV+JtQK3o4HqwKXSHZdB65sj4RC5+cNJufoMUBDouLq4bmiwqcAmP08Rx
HbRIQkcPDySBCOUYIYzI/dJhXI1npmKIDmv4HjEbRoEt6uC1StNWDKUNuODhnB55
D5zjsKIG46TbQl2CuzdoBMiHT8F4aMlmQwpgUSZlQCsHXn+3tOFbFD2weCpU8ycy
2NEjSENgp2VAizdJEPGnz4iLOTaFewqgfMI2WifQ2WQSZLvEZeUA4aeeMjKUtz9r
dcXv75AUSJL1vEB74045oSKX+BnSVupndxqij5uMSzZdo9y2AaigocGm1MwbgYqm
QKpUKUb/ph7tVOxSw41soIP8y9biO69LEkqOdnWRwPF3XrH44EL7dBjvFPc85BVv
1DNo2LGhKYnybbZuMDL/i2ZroacJXKC+pld+Y+RKrhvj1iHNTi8iuL/civ74zelb
Gk2DNxMBjjou20sg0YqKHP/HhSHDjwGko1oTty3EuNojAyxr5lSJTAwm4sCleS1V
jJcBQK3etsyxfT5BHVJQrrTBFJuJU3tYuYxpKYa2RJunMpJLVJgRU6gOctWkH4s3
NgoscIMHqGsyyB5fvo+IV6ei0k8/HiOK0/3lhyQBqY+ZQxV/3WQzb9vpyXHzS54X
ar+zmnCSzgXb/TEZe5s/Ucn9rWoZF9cNY0yyMyO+cj79GNqUrMO42ypDFePwNCs2
iYj0xZ6Q0910+yHLcuIChA22BDSD1RyJ4l2U54yMTPkbqzL9A4sFByhS3q/KXVf5
vccRfWyFuhyUw0dfCli8e/EM6AdKVZFqOraE6+IbgejTgVwnnxRjwPbGvUoH3stX
sDmeg109QcC8Hp7FKQUwZKapdgfxM3xL+8uKuA12bc+mZDiP+j3yDn7OK1D8ShAd
MtJtG0mq6MiBtre7ycf0dkRtLdOydMYmGXv0c8IdtJ/zGvT2uN6cxYPiulCKqmSH
kxN34a2KbRhgqOjIz7qwtSjjeVROi4zqQZVRpRjqNMWLJXSOK5XhqBWTEnI7Nbzw
O4ynFuuwxvesWgp/2n7718p8nE3WKmx+M/+Hve6qdhnhTH05eQilKnhqabYzOJ/K
mmwYh50bM0UOlffGtjUBF8HJ0iuRoQ0i/JvgWlUKJBpo9Sigc6oU+WBsfY7xToOx
RgviMGpkk8OpXxPV1dw3Pjdg7IWQh1Gk4bmhBFJY1JGKlGOOFaN0qhQK3mT7WP+y
Buowzo16o4FWenolEOJ8NH1GqdO2HOZ80VDcTmr0xJ9orJTpOqAjQeA/cJo9XwtF
W/FaBeIEPA0ZiyMx+Mi51efDKJzROr7NgLqRlf3eigubPdVOFq35nzRsZ0dHqOBY
5o6rSuyg3v+V1N+7tRb87qj1raiVYpFHz0ZAnWZVm1rkSYDN8cwegXsHVqijYkRL
l46BPew1XeR8OfnbZUb9sNtn/37vf/aVs5I/jFH4WsovSz2OrbdYWCVIivzZpqVH
IKUVJvXioV9HmGk6r0Wyxh09PX1PWXMoZc2YZzCsm2PELczhDYHWSPWZHeQr8mwm
pzZXIREP7cuT392ZZsGLKA==
`protect end_protected