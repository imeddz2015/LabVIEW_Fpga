`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 30624 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/59UwEX+aE7FohaWu0/8IpTj7mav863zUNIsgIH2BWb
Abd9opeuBjbGF/waQMI2vMJTwD1ie1YueHc3nSNpEh4OXp8P5ybZFY89uyGz3ztU
W1EsuUnchJoQgbHZ/sLbgtGRgsrAFn+ZoIeGN1d6RAF2wAESJmYP8zw+p00RvjZ5
pBGEHX7wooDexzkaqKS5G5YT6K9EPU1+brp0Qt7+0b7vO+CVS7UXBOI65MN38aBn
uxpxjYNVHdG7MhGljirztFkIBp1EViatpMJHRpndSk8qr57WDsn0IX9uTYfhUsYb
ERn9mV8flthqnFmCeD7IHXHAfmzozV1GeqX3RxgLh8QuNSxt4qr36qFmAvmQfq73
GPUWaoiYU5GQAwUZ7tcy6C96Atzs5ATWLg2keTXmkYPlv4b7XL6tN9UWnhC5KdTg
dvS8Kll6NE29UuFJF19gPyjXriclYsGA0ddhRkwtaZHeo548sKIt94Hb6haOEMfY
eoG/xLMHXTAK8C8/whBxQwO61JSGRzo52gbcdkDtJu1pK1drvYRfWnC2KHY5DmPk
M3x8NCVQTCYJC5E5dv8khK+ovv1BGYM3rXmCJKzSunsio6dla+/p3lLls7vL8ZHo
HU91Y3jcNHwRCa0dbdSLeaOP9zaiUytxRGrhde40i9cEbqAYeNeZmhtrdw0gtEVS
p1Evd3r8O87lDlesh8a6mGQocvfUWfixiD4rtgXlfL9fHI3vHD45qYiqbdEgFTTH
w+VI2XBtMtwjhhsSEbyXUr4sDUjICZY2VvV1n+Xl2U+NXpkxQK45IGCM0NSzw/5K
jiHMVMD0MTE8E6tDGIcn6P+ypHdEiNzXiQ3G1RTWxoFpooi/MgIB8pw5lsKGyKj1
DfbvIKOhlAZ4RX+GXk7HLGfBlQv8Who6JMYa7QFVl4w2U5R67J2PDf6M+C+a2Doy
D4F7Q7OoSR00LLK58aYd7KSExg50lcn/dGkvzuF338E+8C19UWin9lMa6lqww9jS
V4WS2uyPpmVyyAAWomvk5lQc/iDYFafqH2zwrxdmxeAAqbbdGjxzmHomWFM0vW+B
AVjYCtMHAuQecm72s83nq/stnKtWbF46jsm5a/PvRdf97sRo7wXpHwdbCr1fSnyg
b0Q+fkQFqwMsTDVJWmj+RLBMCRBrSXCIqMePSh8TjwpTnF/WsYD0U+ZIPSGsCZdy
iYyHDEz4u+LrFPUChJWFdhaltWrqOQ/zdPUWG8EOF5VYpK9JVYWkUu05ZtgEAb+1
85stF36QmOTTC7cf97DapK2WBbDnkha9KxzcggKbKBp5z52s4zYBdeWeA0E1QggK
nfIXM8cdtAC9kZQWXgDD/pspPKBN8iEHk6VitBmLiIik3n8gOSXn7pRG7I2FXPGN
oGuWAxDagumY64mgH6PUiyjD860OrCdGOj8oLF8/9RnIJcdhHdoFSdPNroi4fMNo
tjbCas+/98FDfA8LTtZZij3H1E287jxJnK35sOgB6nHwKOnqivtRYxF0JSmijAT3
UJmKvjwdIyYBDmbJiSOf9MWt+IQFvATsN1Lsq//tCssMLZbq00bizJhIrNPz/sGI
rllotQFvd5GmNTZmygchSKPfOj8GAOWI1wWkaIVofk/eKKReqUIqfSifhbqcPBrr
HAwrWAfYhz20389E+GM8+VQoIfHZtESySz6OdQKJd+M39fvwJvGVjGa4pAgHftht
3cYBFPh5dz4xSs3RqdSVzV+A+u6q2Jm2BcLYnQGf/TbNSBn+2tCN8/e4POOMNpkE
yG/u3S5f9iBlhottJ4YONAxpPMLwJdQUqCQY41gsqdQxNklfT3fkP/gQNN8Yr+yo
q6CLll1vsUSGPUADD01zUirFS3jYoIxCvprNY2q69y3OCziLlBAydc263zY+pHHi
EufNW0bYEA1wgTnH+CRO7v620Dlh4xaITa6kHfRc4dL7Testph8gQ6PK5ixWmiyO
ePQiOcN2jI1JmtzKHvaFieX8YQbzVR0Js6yP0dy9K5Pt/tx7FxCr8djmO2EsRDNy
7sY8ydhGaH/pyRvxpmIIXZTVa9uyFneMnXw46aH/a2KCQ0X+fknoKpPV8xtpCabM
zk0Hf1tEtHSMOp9vSx+OytQmeES6idUb43wtljvz1nLYYSApBKNld3Er0C0SCIuZ
OSJKsxMKXcrda/LpKApEkglaPsQaxKkGVGBDMNMg0zca0qUWQuSR1bU3IAEBYNsZ
iApcid2ciHPZGk92Q4S3GlbyAy8ysmQEH2Dqnfww8SO6fTscuJ4nD1TlSizpG+UG
mRG/fh07TJj44nLuTPuoJIlxNi29XHiqJXJIlMAz23ZSqcYcIfOuKIOAOhjF6rcK
8/Or/X+/GH6BpDgqvqoavGpJILQyYIc7VoWqP8umo6jP4UrTfWCQoQbuJBO0VYFP
o8oVVAnMCROCRv8haRaE7NXn3Nt368E8zq6VXxWkX1VY38G9AWoPni4uc3Dspkhs
zn6c53jK1e0vs0VM6KUmGgkcCM4v/+C74ZJ6eN1Fk/AXK4nIFRhAPKcsWg9PvmKo
4oD40ZE9Q2fuDoYWV317PKI5pEuOHTC35sPPnEfSrAhE7ZyMF03LpKtKvISOTcVu
aKIAc9SYSCVDxFkzdpQdJjsBPFZX4y48b/Zm46dWPscYZv67Gf/267UanJtBjdHL
4xgzJlImg9hjluwDiwOlNSrv4ZBRdivYEPDis5R1BjCUj3jNSv58J1/L2zyQDRrs
a1HJ4A6jmrXmX05CGGdTDhRiZMh0wZ+vbxe8/fpyenFDl5I9xjbJ2vUDgDEwB14U
+yRGPhyapmLbY+tVukxGdqG2jdZWzvKSrJzIt6h+AvgqQzhZUy/llo6pgPhSOxXH
0Ye/GBaDqSuC2z+Nhi10Cbm7ig2U769zzOQSECbu4f3VkALaSdh/hkSuKO0P2xjc
L3u9m82lF1VzVTbbijgrK1TRRXy1KPkMybQw3GHv8smQb2N5DxYcmWLg0+CFVYH2
ur0KfxecelLlqIcV7jTG+LNTbFt/RDZtxlaWHhHcWbWv1x3/79gG48PpVafqIF2m
6jCALd6OW1+vSyG293wjCYoIb29j8zM00FsE3TImXkmXrfgCD2otN9doOCmCKxYT
5wrsYywmlf6amIvlX6peMy6dvg/yDlL/XtAXPdel7yBcvQ2cN/AjmNFxYTF09koD
K7a8aox6XYzRXmyvwlhyqgpyqPjXo83xnaVIcKri2NhrJmCpH+xm1Zu5CgnjkRSB
dkqrwVmnknkRPGzDAGHVPa7cCb57r03anTxMj2h/GgbvrXP/Hp5gmNIrZyFZWsiG
oHWKQV5LBbIV5hgNy2XM8Jkr40hC/Hs/Hr2LOBtAbPsQ3/0VhDsmMLYfosB0asVS
IXNwpbd7ifLDy//yAVGY+EEY3RY/Mh2QXBgriMOUjPZRadka7cVPHwY8coXejmF4
h8VheLwHz7RQSqn5tOBOawjQuSo3kvk9DDRfypLr0yuyrsUh3IwJgVLLRGAJXsKN
+PGHcrK5n5iJh9v3gtOPbGdEg81hbWlFJFCENCvKGj1xmCfR3lZk82WlmGnlc57g
6rRAgivXmcpaEfdlBonxUUwRq6qdW8beHQ9ReFn28H34PfYSHlUaA3QaqHAvONS9
GmwiGrd+h0uLMjF4Gi4b6KXA1Cqsm/BLai1ekgaRYdGUDy2hm9GzbqYIue1Yp7Wc
Cf4CUuseT8pAsrAUVbGjpkbALVHJQ+PQ846LKZtVofUlHNJbmYUv/hTmggncBqrE
OFpnRx55bwS6tLXNi33ylCEucmQpMcmc/9s80c3mB5mLbbpqEglZ9lcgWEwTYJDy
oFFW2jTta12oWTDcZKbaAahUhAWmDuM36WPHsjOJ9BogAISI9BuJZm5IYX6new07
S9L1pmd5SHO4GQRloPJtLFROOpY76KHvlZDxXNiFskKOnVw/Z9babBSrLfnnpAlr
UDDly+HXRROWLiucD98PS9Om6pCMsYUpBOf2fFs++Hayfauu454729mJkRVg1358
letBRtWCqO2uSFVCtK4PuF6bbkDaTQaSnGQrJfTyYBiN2AvPVsPN4CnAdLzbO0Jq
7CPUZOZmumiSCq170uRiTBNBd0kqU8fVUWtfFUcCa70ZLP9UbyhbyyuSfL1vpY4j
j+DaXvn1u2kHBX9FQjItKxJKZi0xR3tkoiEr3ZLK95pbFSm5gMaZi4Z34ujE9uAb
usPwuHK9/tiwkw8qy9cOPdnMms7qKrc2fwaswhl7eaw/mY5DVS+cWav4/sFQ0uSK
S8PVxSE6IBE8whhiPGkKhGqHr4pFtDnndRASONn4Mn9serePumTXGK4cbtn9hjwa
zxUm08Srs8jpRb71IYbpSu6UtbvQHkiPwbTEo7aYVLS5wvt5DQ7Ix4uVz2DrbGRO
0dQJZySu276vkuAhlhmnVOqxX6JPzj/sUrp4Pw5OtmR7Tg/YZ8Tq3yPWzHp9a/oZ
+BV0P0Ghnf2mZoPyxHUKUnCfZS7tcNf0+z/glkvcwBKMrBZq0tV1H37pgp5YAinF
rCNJFnbRTNtEosg7Xk9J+yoBm4HXF4L6Aak8TO0lcC2xxtKfJtTohexrsuAF4XoK
fcPhhq4nXLJ2vQcVdjp0buGdvCiCp826HvSdN1fEfwPB9moILVvvJ/JoWcXv8yHH
XTds5oiQjrR0kohTym39cVG4sGDFskQNM9RdgZ1SQ0RjBhAaWMdcGdL4SOn4njlS
LBp0aQ2aMcQFFvUxdVy9jC07qBgC8VksaEPTfboA5nL78hePYIsnbVgFRLY7dXCf
WFkNRZbDK+ZPhula7M0QH1ZhICHg4H12XdGJDubiF+0341QfZ4ch/8PIJS8T5NGy
6WXVAu2m7et+fMsvV79hXqodhIJ9QC4N8W9gqJXEVYV5Wfqt5ItX4CYJekq0bQCz
Z22AZdRRVeGLO2M4DwgHsYmvc21+42smXkXHGzJVM4eF0UBoXd4hU31OBo8eEE1b
n8kqtbJDBBkj/Hy4k795z9Hfzh2DPOj5uc4hAXJCREfCBvRDGm2i6cX9DKm0ZkJR
HHEIrdArEXkxy56863q3p6e4zMSTirJLF5PbnH+qSrZ+FYCvR/e+rU8qlay9s0Kt
Fjqp8poE8yel5TqaLgswN1tKqilyfUIlLIfvxHZBh5StKbxZy+zyZ/cu0Bc/6JsS
ST3IQ75WlGiysfl7H4v5c8e2Izu+BomuH605jofz06iMJBJW4Y3RVqFaNNT8QSNI
O5GCbBPdA+dZsl3AqeZMFQJUU264sbIiCIgOB04l82MMf+bNdZOYeb1/kybG+SlI
XAwBqrKvflzNKX8ZjFZ6xzbLySgG6qfLJdFiK1lfLrMr09fM+YWuaFdcd1Yrwsip
v3Y9zz3w/6aMSD8weN8WbTPjY2aPU53XZPSi/uxqvQtVT5u0V2sfk/maahmbAvBu
bwo+3s1Br5LtApvKgD4kxVuhab9Wpy5tTdFCHcjEeeLw58Cn+OnRSBxbILzyNO28
M8qGzoScLOKCpru4lS2cJKG2f45idujlIx9irJjGtyy2avpkSrQ5d3n15Dth/G1+
OWZ0Um6tXH7UmBt9NRqmzKWl90uLR1Jy0JNip2MZqMI7RoUxobVWvRQh8GVvoDcY
fxwN8/uxHoZxc2sBYzO0c4tBEPWM7RtcbbNvqHLMvdRpbLJwx4YpcRc94E7N3xDG
luSDfqwWDtnz0uPnDVNrWBfmSFvn5vUc5KaDwO+C/TuZVoOPh+6j9kZn2bVkEVuO
oZqX2AmOGD7nK4uTB1ruJ2r1oQfMNOtTPstXuDljYuamBNzMXSBSzrZRLogO5UtW
HRIgfVApO+cnTTPn01UxHS9+LH9Dhj7jHihY/nj10DDAd0NwoeeA1FexDa+cwcoY
yVAEt+K5ofhM7d9yRu9RMlTcw1e9dkJLfpXAfgqDVIQbR8xr9J4pmcWp6ubBgKJK
rVoeGrKNSp7gkkuwsfnWhRXTQyjD8NR5gTCep8ubfKjhFbIm2ZfSFOcdZijSEibh
n3TVB9q8VnsA0RtK25ST+eoFvj6qt7CRMFKbE7hb6P4cMeHp14MymmSBgQFQ20q/
jbcTpz4QNqnlFmOb7YObdYoLWHqmArqx5evhytHMwxTu7+O0dZsA9vEr7CoiBfyW
R67FR9XZ0Urbi/9sjO8dESybTHuMhTnz7F7uM+3m6xp8isVNYWbs0CiQSvmLe83v
D0HhtZFlWd+1Ssn52uSyjk/p8Sr1S3u++K1/KWlOiqi7kmydxQmaniHwz5Lkemz5
Qm9jIRj7O2IelmhikkXUKAGIgQffbePL5M5tEFvYnV7uWGFEx80xz4kaCshav4TT
6z0sqm27njkhohOzaYBvcXwAo8kbJiiLGwDWYChsPgLV8kZ/7XL9eINwKnMvlZq9
B7ddak2p1hPxlos9bQouKnSxChUZRxQ5VlbERCvxua7pBWmKS5vgOUJboC0+DovF
CjQssciH8GkJQdD9ZrbhCeT+oS+ALj17m58gr9RdFEk6OdWDf2ZJsk3C80L+bwno
ftJEIbJkJWtxVFUxz+N+1K080F/O2ZiKmOJA52pY1fJw/fhf9VLxIK8AkJFFga87
lgLXFCuf5KopAHRwIQn/GVOsEkGvxeWTAj0F45g9Ci2cIHtkbWDSKOXFoqrDFBGK
ckmr/kAgzk7eba1eO44hztdJfT/qqxLBwEtijfWmteJjML5n4GsuYX+GfEC8Bt7G
99NG2BgIW0npZucIbLORV4bOGb1D/fJ4XFnM8lqgHZJOrIp2h51O9Gmj+slWnRjX
mQczfTN7bq02Z98fjQK7uhwKkDDsVtMjjSDQOwVt/giLAByvLHdadDxxpmoKUA+Z
wY21zQkJYgBXmsI42inh+fnSqFEbyyQq12ekfgeaZoDWixzPJmdoc0+Alen+USov
maFSF84tfmg3SgdRiemzOL8COEdZe7lZwOtITSjMIZ8AsqSOAdtiLcNQ9dr+wBw2
VRYyWGJ4yx3gleoHaLYNuAgBW2vHKe3LzDs436SV2M2MZbFFxCpa1i4j0YLjNpSn
P1enZgFBvFoHvZFrIGlLVU3z6b7hwM0laxFK4Xq29gfwiM8E5GndWHSMj0RzooeG
CToW0XoYIQugNJeOL/UxrJuDR0Zutoo6d42DIuuwH9HPlFp0ZsfWiM85gUMMBn9o
3MZT09JKXqNHODvINQtuudqytTfxrlL5H75tWR4cUvUkG9YjIf2OP8AcNZ/RyjXV
2oaC6k3e05vhzLSoLkFKlJSNfFowYHr/RUFs2ZXHfkYFxdsvTcHdUpZLISRZgs1z
9PJyRDxbyG5QdmCytSaypMcod3H0BT8SDsXb/RZoEiwPQ3E1UCIOMb80H7FaVeY3
zxgn7RnjNPcAzP/tdLXyp2UKz99HPqLZQmwPPF8Xu7ksoiC8xhrAfX6RPomTVlKT
CshABEAWouYZ6DFLaK8cM+6Q+EO2Gk2zkoVGC0QJT/ZZzVK2jAoKyTKGU4+azyIu
t/NOcjQ2X0hJF5QaeDRiytkXC49JZlPOpki/q6S0ZPdZUwVqI7CN0/abdUA4cE2u
87oSa39HoJzYGod8U3TyyWgiNsqswHaQef8tJC6G1p1ZOJw9WnFPqBzcoYeev1IK
iioSxxzlA9/o3zIWA5qpDhIh6aWnUf+bt2vHcMTPpdYNzTvJijxeV9n+gv0o69En
5t+oMZjM/AOfRqFYnxxyVEAW6Loinc4u97xHixxxmFD2ZN55V6mZnT16Kbx+51hV
mwWDAxvAmcyBA34eiDDB5FfcKVWzaGy418dfr1IXiC1o48riKTCPg+O5e+jT+Kdp
FDLfo88AC7H+CNoHLs9BnUU35IKFvZ7K5JXRqL2lIgnms9AOyKvsbtFWZ1dELMfT
Uvj9FEoAYhJrGqm7GyClxZLJTgdvzxz9N6Su4p05nQs1Si8BkhEUUPOiKXj3o5V0
OUKglW8ua41HiVFCtCeuJOG9GTyrf6PloIKhJMgNys1eAfnnMYA0Z7QyHMASY19x
QMWIXlt83LqvTHO+eCKzkPcPZy5y9yApKq+4T0OnLdaEoIWLYyCEa3c67GSBk4+m
ygfl8q0xFbU0DHlp+mwjzj036cgLLjlp1mwaCcmwNGgD6im/VCEoOm6kP4W05za6
sSsa5DjKvZLLY/9Un5g6UuWIC1Y54F+IMIloZQpX87WM9pg7ahrJfZJL37WGmYEr
o0o3k15ob1dtVbW9kwPjr/XcNlDPU3+iQf+W6ZLDVkHIF6G0INDJNtZxNIH4G3uH
r39DBPhEjZvPYjpYHKKXAb7dcEjqFcKaMnw7idGPPk4Fwd7oLJBn91+8ZkTxNG+U
ScZAgqEZjT/nYZqXbHmjkTk1HZ9O8PixLxqdJSAWnZF3Q68bwzGG6khVz99RVC7C
mzFrpnOokCs0kUOAIjK5FpXDdbDptjM4FfRn3zSFDu9ZLSwCn58TPpSqqijVRXUT
yX657wTL9MsO7D+l7N+x4ZtHO/dQsDozcHSOBOAzhpOOoqj+DsxM9IdYbPsnuXFV
KYa4vZpySdsEBOgtiRMTtmSxT/BSyoW1+Ju4N9neHXDfw9aHdMrjgJSVFobLKCYl
fd/QNAoMNnow58UInjIsR/npktxs3CI2+7tnaQ1+kgWdcVywEwCMtMwoE+zeZfQq
PrdV6rdjxmr/o0FHAsNP+xytmmTR945DNcaRjF1w4uXJNHIIDjfV7HtwJR3r++Ga
nRA2Z/mOdp5pmNZFjt4ZU8/PlDmLXQqqpzuCsG/Seg9jHbjZx2MiGMtjEv7tZ/eU
SUpdR9UMRp0Z3O9tzgD63NvM7goaByZY6BE3sHVBYLuJqOpeIOPPuVJHL5X9Gec2
nJGOLmsGN15CBw/Yd/wySbFidVM0/P6WbB5X/F4efrQkrxuPqaxA2ERnjrZMF9hD
sFFipOXbLeomgcumIpaWEjOH65wHCpcfd6O00cM092y1sfwHVPThH5yANSPuP5BF
4WDyjd+0chzvS8kqp1WS400/IwZqgjRi8B1Q2E1vPEnJrFDV8VKmjj7DjSmf9WNS
ojscoEux68vR8OEEXVsXAb/gEt9Th1uEgB+RcP62hP1cvAGwh6nyLlLPuK7lQl3R
YILKaL24n2uLdb/dWxR8G+HQQEvVLveX5OKVsOeg1TRutXy0RdBrqL56ynGZzJXy
dZq+K3T7/E4rK4+b6zpUSINF4azhsjSOx37WK6T641nA901txAFZzcvuFDmM0t3o
0AxfNkybzSw8zd0Ni/UrCVKmqF0cDLR+DLkrapIq52ClE0VX2wtpUbBFVcwHfpj7
Hyf2/1PtCvM0E9zcbRuNy/pSrTT+MkmIz3yx0ajgmR4/fP0AJfTT4y2Fl7j5/KIu
yHcLua+B26qTJFjv8AdT+NZ1IaRDZ8bD/0cDZYgKNysFNyKpvRkk0BVgUvg+N4hA
5q2rSOqvKDSknTroZfbJc2/URohaUQ75R+YTX3MpXu33wAjYSugeWZL5uTbpUYpy
T3oE1qLD7Lq7yareudTJLXifcIhPqdmWtImmMPxYHRtR2lwJ0R7PlAD4jM2F2ILe
B+w/8QWYQlWvVMoj92dvklrqk8F92UBUUgbafnbyAmDRQEX7zwba1ij3Qat5+gRF
QIxHRQqBsatnRNEoQZJFTQaYnJMErGCpcZmJnDRmCX4rcOn9bwXS2aS35zfN9ohj
JWdJWmKRmDbXmwJqNURqqd1X1BPzeyCcya0qTlvp2QflUomMIkqxUIhAXRY+v8Fr
bwg7nGUDNZftDdAxlAKVxzE1GJGfr8tWObafPAGOr4VajSzAPGYiHslDrOLBaP6V
rh15W4o/1HSD4GqQWDrHpeRVqSAKFbpiIvmXiS56aFyIETZoBo/qpKJ1IDh8B1IC
RkIBwDYp88MTiPqfMEULm6XdeQPmGCoY6t5FQf2YzHaSAp87ryvtmWi+n9WSizJS
fKsQghmuUy51Q9T1VciGRVqxpPCBr0Fa3mQC6C1UZ+CiqTAZzvdm1Ljmqqvp+6GI
yJZB4ZLutmpG5R8HVmvcbQ+w3f0n5CkgC8xSUrnWeaoQrnu23BlOJWUFBYB6f1ik
5T7VA6Dj2MlVWJixucqEx3O8wrqVwWWE5K871Zev+fIYiPQBrKvKW/ULq4m+zeMG
10nOI5QvYgIij1hi7gAOCrlzuBVRLqEQ9kOqJgEaDf0sDf7FC0JAzkkh4TZ5kJV4
QuQnPgninp5K1u43DEwoENJFU3hDJAU7MtBarQIZesqy87Gxv10bHZIeYEHE89GD
waT/GXV6kaBklHGaQhdAioafIFslPwnEOXNiozAKcAacEEZFazQggYyHNgwu0kvI
gG6IU1618uldGvgnOQHnjY3BQ19GaGchPBvPRoGULMkLeysyb7CAI+xj3dcpbnpZ
lt8BpZJEWQiF/tZB1Cpv+9NzfAe6KfEdXdn2MAgmmgDqFDUOPHYfWq+F1kt+iDyR
8JxhHdk21vV52wHiqnNeDm2w7nqYZSamWKGP58a2+h+kIPKUHdhO/VpunT33lFa7
8doBorA3/y5052dQYyPvpdpIDEm/S3zbnSvCiI5Etegz9vznqwf6Mq/07zJKkKOa
2xsTQoxNbTM9x+ZCpr9hqa+A86TFyobbpHVRajLjqEZhj2gpNiU4irMsaGVD/wHb
aW33i4n2VKCp/GiDRr7PQXsAobXldNUKuuAc6GP0QR2WTmleLcIQNNL0TeB54Bgl
DuXe9s2tisFYxcEfcpKQRIFF1m7Z3QKexCAuds/N5llmBE2MNVloRSPhAVK4tshT
tEXG7QfzmwSjAsM+OqK5wbul1yP0X5j25rJtd1J4fQLLJR/X2eKoh/KNMx/N+JoE
9wWFmkNrl+mal8sH8MLH7Qr+RwMyBO1r3iGUqzczyRxr7jyfP2aK0lsvROR254w8
Vf9dDo203iB4ZQRtZU5+E+C4hhs2O3XHO+ZfoU5hDLwsHTLwhOyyvRJOxqxE6goo
33QV3cTPCbvDbOXwqkvpFCOnWuXiCa5Y3kPPG9MjW21sI5CWcPVo/s21NLkVAdq6
u27Z5xISm7by/RpNh4qGB+4ySgiTWK7gO9MNXRzRDe+DdqHDrqhFhkldebuStJP4
QztUtd/PxgsTuAg0HT0YVDWJg/+H6PnWC/973ymu5I7vYtv/P0LpwZJeH0OuJAtK
ePjfsJrD/ykCuGGmdd2YruXF3BtABiS/Se1MTGBHjPhZ+B8VQ187ZlualXKt98Dk
oWdDmQXKCParZZ/VZ3aB9Plev8ZmKkaZYcLyM3/3380n0pumMSTbqvWe2uKdoqwQ
H8B/JYnkYpNbQPlrxZHq9ic5kNFAEoZhtWI5dCDlJE6DJyTxuMQzNkimLziscFAf
9zDvYNusyZvRKST+ugY4bmLLrklHcsAryCxRFGbgQPTvJoYkPwLaB2qRVw8P/KYI
s9ETj2Uaf896iXv/dehk4RxEPmIT9tZ0OfAz3SZt231RET9WJgZYjmw+kEinpyfp
UhJ4m3B2GzSX9THdYje5CVPQQpVO6fNsDUosf1z+762ngOZfGmjQeDoXw0QUrpa/
P+5l9I9u+60eyZs8hfplyVS/55jKOYdga5sq6jYd24CF/d4Th8Utt96plfUrdIWm
WlICsDny9E0qXnzR5fTNbyr2jlWA/b2jnbki+2SsLH8RXuQwsbd6DI93FiW/0tHK
V6mQqQR7pOPV13/JwwASj0VTrKzy3y1kgj3d5ueJiGSk1zrBikrgS/JHjyb01PPr
pM7Ee+66d1dwpBsVIX79UH27Ey3Fw3NUjICB1i4SYO2cmsRpjnUwuOlPtDaT6tFl
0pnwtpCjtrZrXropIAynspi7wfOlDtcxZa6hoLRfGSY1r9I+B0gCIRCaxlM+tuG2
VBuUs3TntqTSXEOkDnGLZvCKBKS0jP26OnNCSuNeUiTSMRe30tZvA0dYX9M5Hsly
OeCT3WbcYkvvbstLucXp7SUjUr8rcJkmm2sVudffiDwbm5v45N8TBfRGIiY4A0Cg
kDdrdyCIbIF8woUuUu7KSR3WjVdSg2isBcmqzDILr19sL9pO6bB5uTtSIcJtMyPz
2j79t9syT2nYSbHyzD1Z73yZ+hys5P4epNbnp+MsZtc3th2jb6V3YZK/NZYydhX1
6yOz2OUxQvSV1Pe3u43qbiUIWjbvOzGghqDx7QfVBG4IsaDFnqLsCl66P/sFSEqd
wtpOw+bcz2uJP65ADIaXdb/7eSZ2XzOdfhjgpcyD0LJl2XrNN3W2Ee9opkfSGt8j
AH3Fsygl1OBsdCGnlxFpyZ5fd7CWFfXxklcoyWDy2WvB+gA18c5WRO7FvDckhKY9
VSnigBDeyvp50VadlvOb5i0cEO8+qCaRmAiQUeAVLbSN7OnmRaAmDi7BMZCEdXxW
F/XsNrZONWJppByt8V0QI22GUYYDYYUeCfLzuMLg6RaFDWgomcrYGhRZx5EVHsSO
5S7XtOFL9r0lW43MNJkt5dY7GgXvcmTCIfVVhBOmr6WiOE1/d2E/mIBGK9dFOCAg
9jXOWb/YtqS5kC2Mmg97p21mxd+tndy8+7IjVt11PVw409yVRoT3aXUGehhOaEDd
SVd63fqVR1rpxPWDXZLIle0qCSNMQyUNShIJxwl967x7dyLUV5l7hZQIxIHA7TZs
K0U5OsnP6q0YDwhz3N10cwDA6OsfYEhU9X4kq0ucQbmAj+U1G3vKBuRfsBkTxKUc
ChxNGOdoxPc8sOFvLVjBDkxmTxrOQAc5u+TL9VGX3WwZw4y2DQFOuA/Wl66IW3ig
sYoXWFP7eRA4snr1Pf23H10b1gyG3VfSxwUuJzJnZsAxo6pfAfprQI63FAK83kE1
6eEtBMzKAE3u4J2j/zF0fxFvnCt2LVTvC+BE0VhhbfgUDCrLdcbeTb7CC+EK4PDN
AbzDbCvZv3v9jXUpMwUBA4eKzyvn6SdMDaR9LDQrwyBo0LDIX7rfhdtiGVxqVYkG
7rRBgW9tXlYAMuD0DKp61NAwu4xvsbaMDqYVZ9e4/ArILgMx/TNKL+0lMBzLVeJK
M1HEe+ZPwld9PT2TXSnZiwSrKMKCk+vBaNVLsF9i8Is3nvt/VVK6ARSVe09LiD/k
TbZIw89fH0k0fVRjdg/DY4WioS/l43Rh+mwD7TtQ9nD7/i89Cj3+pA7j0QDAtLMS
k1648nQ/319VZ6k9n7aHBrqMht0seg4Qt/80IEPvU1IgTY2pz3UuUnWocIYYVbAd
I4Tpomn66dC8FnYdsYk75g4HynIe3iZSq9+rLfWp5pdI50Mr40un7N2PPhFFExkR
PP0Yy4S6N2EOHK+hOhzORK8IvLcNVJY7N2c/BLiDHXHTFBbWWdtdwNBJGZyr3Ps/
Nxr3ZrhZiy/zy6FBIQ4hkR23I6CJoUdwLAyseNWc1OOW8+9jM62FmeYsxcFu9chi
E6v39dH40r8IIjaePeMcctcxjbcAd5lfjjpSp6nqscInCEl1arEHVdW6oeL5vVpL
OP3dkBWCEYesUVAuUYIieTKX0y3Xu7DV+U2DWDmLwXhg7TvGizsXRRpL5SIqxiXz
DxiEPzLWa3AgkCgUuPSRmAI53aj3dhiv90NbZ0FjTS1YRJenijVlNBsKzz0qO+9Z
2u9JpJQu1kce/0pyUcFFq9LnD3vS7WKL8vo6528uQyqA48njGOu4Yh+Kw6GDn3BK
tsfm/5bIy6CzGQWmnJ3i1DjnsYODMzQxKkyaQhWy7S9/dQ1AMMiL6UVOfDAv09L5
8kEJZtBtIoiF0g0tNCpzzL22JoikbtmkTcRYBopbAKNTKEhPUkvazp2DGa/0wT9b
ycY415ILJh6GRG3tGJ+3MQ0WOZCkNcIWn0onjFUMkkXCGtZxK+pTiC0mt6n+hQ+H
tZiYak43aLC9YE3NhvX4HN/JBYW6V+zGqRGSVLagvEyq8kWLlLt0TIoll1xlX1pi
KriJTU8PbRdcaJ3cDIPiMqBAEwTBgwPbIAyvHOHOnaAWgi56lJ4jJAATPAs0856G
Jx2VfW/6ZCPmSZHEtO2Hg7FhoJDzVtCUrnmGdJ/c4r3UXYIpDaxYeEA5dvNY8BfK
viEp4oyuSJBojm2ByTj5FiaYD1sd6QVA/MC+T+TN4os8MX4HBTrIQ6uN2MwmUIxU
w0Hus1SK3F15bkDK4IA5bDhxrA/+8YIBhzwum4BngBftc8EdLJidwtPkqZd5SyU2
Ir4M8Ct3BpPZSwRsmojvy5yT1MsPvPdtt3Tt4gJ68/dFSH2heCJ11+hVTjX7RHFO
QS+1UVDFX5mqvJMsxWJqu5k4MTK+eZfuc4s2ANFKZsQCd+xuvbcv6AEUQClmsZzk
9nspUtu/KeNICNhuFuarHBf6bA66Dan+/JsDgfRhCeAxbH16NDENOcSINqDhu+Qf
FzIJ5FrgqrvtQTZIvALqMCb5pzRcCl0/fdj6aCQH0iJ62WzZcIJskQsE/iFEymWL
EO9fPRRyrZ+JBSYBPtNsOss5z5CzZ/5xHK1AUo8HgnRucCtWIhx8yWKzPExX/Ozh
NrEmVGM+uHWcHeXThROCYAadzpIkqwaIPzlSckylKrTmQKYFfTptDYt5a2PK6OlC
y5Y5oPulq26T86TO/SbUyjqe8ph3ZzBhcfw1ZSAxpExA5+tDU6O+GL5JOd3rMJuu
0Dwwy1gLl19wRmBtTPZPdyrk7KxyrKZ1wF7/KpfMuhimmxFGviOBY3RmTFf0f7a3
t81KunqFSkyuFjr6KLcGgBX0NKOV0GB8qJgpyG5aw78IpYFFFcc4FPN4ySdZCtDh
OrF2ng2fpUHhE19Y7flmrRJDJid49/llD4LJ3PCL3evmcoZnT7AwwqbjBCCpOIgT
p5pFDpUInIp98rSHaLVoJcnfA9Ip1TqkI/cRsa/tCIZmTepkk8ISSc9ktM6O87lS
Xat41i0RSoIrkR/C4IhBKFrXgOInkOigzsLbPEFFToWFOqF1shNjdifKeI04z0Q6
V7ZmeqP5DGJyCT6WYgxZJcdrMCd/HmO0zKJkty8ZRZgFS94KxtOTNNOcSzyXzgvQ
4wVdTJND5LPkDURcUazFEnhqFz35yQr7WD8THl3HmDgT+dgWgjtRVBqrZdCixgY5
Nd72+FbsuRbRUQgvnZOeHNap9dSL2bPNSTUMBzmuvh+Oani7zkBR/k6gsCvSS+Hx
EI5pVnL3UVHLkPqavN5Ph6MtBjuJv406yurzpzkPwXkKdvFmcSFLF8AtnxTgbsCh
NAW/WDWwP67MVs26yf1xVsho24In4mLd82Yza7396zxnGWMR/NUXo12pfD7yiYNN
oOyVXA7aIKYQ3FikkHK5rYhg87YIjrT41s3NS/hOOzvF4XqHpbUrsf3QKfsBTQtN
baFsuSwPlR03BUJnvtl+nqJTCWHwWRAP4TfpQ6f2C0BFpN2cvD4PQde4cRiH4GtH
ACj/IvRelLHuqmLoIfR9FJrSJzmJgX/xP3tUnNxQ1+3FKZ7mDeDygFVscEinQxKt
set2lbCKy4/jRZcui5zkj6nSL90rqdzwo8UC8D8zbcXsFQM2Tq8xE2B9hGobg/nk
8IMJfT9bsHhcIqEY/l7aAqbwVKvXNTkgj7thhmJT/sctP7XuUNffiHLGq/C+nj4N
7+nTwEAmRcShnA1mMwaCatJth/Rmk5ONnN92bgehhp1wqKeGwtLC7XgztNqhnVvV
ktSgOw3RFCGqt/otK8FXwqcXqbp0zZ0aZsbYu4vsNTM51dW83vMzngJMnA2/ROPu
tqWeXdoIrd+aC2D4p57hc7QTkLwZyAybXJ+m3qJioIl6vjvV6ZjPHoNjM45Ekq2k
FFU+rf3NNP+CDPfVhxgrRywST0Fgw9M+CPyFVqioB3xG3q4EGDaYGeHsjwl047ni
9fzMQ8LyBpRtBcx76rW1N0FhCR1bdJtmuHDV/D957uGjrFE0gemvEpuL9zKHSjzR
+o5ewQMgvkj78tRVT5/hv81kAAgqT0epLcNHrapxg68DHuuycIBacpVVpdP3edw2
8RLMkzRFfTVEAT8xqTE0R8BM49NBVibaV/yYOekmSINMD8aXxEET2wF/GVnsV8fV
XDM9A8nuD15bGn6qp7TGrjBJE+leUAcpmyWpMZO1RxDZHuQ8WQoCbPQhB/BOnRH7
E4/3t8cIVEdOMllJXW2vPIU3KKGnYViIVEvZS0hPyVG+vcm8G8YFhe7gvVnIMlKF
Ly3EnenG8u3jPrpuiBqQ62xFCXp3fF8pC9ZohqzWxBtZPxbXYfuxs5meazbQqKQw
tgGw5R4hHi7Qeo4OyK3CfvY4awZ9I5HNdwimAgpbClOj5eNAkic9y4MIXEWB0CME
tTYTq19ZAPg/IpL/TYG4RQHh/NnD4u+Z0+aGId72jv7o2HoUbZ4FUijnQSlqfmDI
Z1/di97Y64oS/QXcIHd0ngNbyRyH7Kf5IGHjNdEdr1I8GjiCiqFEEuo5LZsNXXFa
1dZ8Wf/erpxxw1cBO8g/tt801X/ctWM3bd8CIA5E1x+yLxakcIbMX1KSwp4/jqg1
Iup1C8KlD6PX4krQwC/7/VDEEY6r2ReiEi3le3qn6sBmJVJie74+QqB4z0vjLH+W
63HrmnTFwaCph0n8zA9WtExlli4cdjcTz0KuN5iLIoh8SKNzf8eg0FCBTDX4qvEi
URXaJD+5YGEM4GKhm37/axFza1db8FZj/xmNeH4sT27ZLBGWedM1Yd7iousTMhys
PlPV8zbw9lvKtmpjZrKhlT5gkhnTVieiExOHoKIiuCboIJW5qHyoI1DiTyob5J6X
PlMUTPKnDdkVYm8aUSWX6NmYBocchhE710C6yhZlVg4oGc82quB0oF0UOQYrXhSg
Yara9xAA4nwrrmDqGHtrtasE1jH1j4qPSUilvYA0xwUoAivcIVT56cbloM3jnl+e
PJU22jMPnwirtofRCbKl7ulJFKDAg32n48x2Kobic0LNnK5UA8nIE6eWeRImIVjb
LuJ9WGKC57ap8h59vm5P0bBYJwk/N9hRIcF1+A+ngVjAx2kW67AKMJKJgjM6/zVU
7bSokLaBCZzrpujjd0SZBna4jGtY22kFtBz9FjHWRgsck8FHErFI/Nb9ek2LuP87
Ol1cwuqo54v6EP/vJGm7z1w+t9+8k4aSQIIJhQSxHKJqkt+KlMvRFshnOdVEZKMt
UFPka/TrqIsuZLJo9gxYlW79SdfbCXpp2vUHvVrXRfhttX1rCZLEqdrk6eGnxBOK
Hp5sexnJZCHbDOUllLaXEOLCnvo12LYTSu0NtjhoDUvCbUvRd7TSG1knb1DNZ9gv
OYoW6bkAI6c1r7VXQGN9pnCruksmWJ8UcsEyaTIP+95t2ocsA+GdSf+3pPYkmmgg
Cb5wUJ+WaFLPTW62vDaME1Zz1ztDaQWLQimZR4zCArit0G0TvXZRl8k0f+sIGJnw
V2iQt5eL881f5f+z7eZjQ+gSuZgG0AxvZzuMKFnokTCepkiIHCppPB5WbN407UGA
ADiDHLhGKKOWxk5jSoPiIaWE4X+u4RyhGyVrVnO89eGXBqLUmT2lryEu1egpqTWu
/PZ/B5DiQ32uruSYUDQVH7sK6cqZmnAPK82Dvv6ulTCcqvs+QfQB9k7ycddpJeff
zqteApBNRL/s6irkhOTdwf548O5CjOULyExQPh/5lhdw5+gJ5gbBxFScAkV12IG0
LJyQ0wETTpFm6CUemfh0sX/2/bJu+cS4fI+zc4COeX3bIKDH9vVNYhMGFHSAsmnW
rCQsliu3e3kPfBRqdWOb3UaXXmwO3lxz0vKt2aKHHWQd3jG9zLdJRZvrYxVV/Gs9
gQoSZDQZ6L8bjzr24WnLR5x4XNF2L+NGb+4SjaFdSq4p2Ru09+rgJKBmii0KkNkf
G4/rZbIO1k0/G6uqJgk0W7K7KmORYxNIBlXEdvwox2Z91+ijPbKqUvT3/Z8P+tPW
skq8Q4GOFZGJ0PBlj8DVgQZRPv3oFQWZrJz4HAw6JsfOtoGpKEttH4NtG1atjlzo
z0KWlJvRAOOCQq5SDQVD7DA1HuBIgxvuZGlvGP0B4oleblnD8bhHCx1huRGJSkUZ
M8Fuo84pZMycQ72kstmi42OdvJmeLUUxkh7bXN7UXWHWL/zfH1XPuWbcnaO6Omod
UUBzu44tT25v5j4iGfWAzeIoep7Xg3AMnvuoNQgibkkwRmhTNkbiGDUah6cs9ujC
XBk6R7DsHz25hqFF8hjEhEWuduYv3SOq03oPyUluimpQ6LH/XX7tD4S49idjzoRC
6pZCurMN07rpVJ2CMBbm3j0OIu2lQCKvBDMHBJVViBnIfEZkcz1b8S6KY2iO9bW2
Pf2dvTL/cwibg8sy3/ilGs7a5jw/xl2mJNshNh6IanUl8KYrl+j5/n8anhhbkjaI
f7067kJvYRHhjIHftvrKSfMPBK7GHy+CB7yHoNHumReYcNmDMtYDLUx41DuLfo1V
kxbKQnzqMQoJx/OA7A+3nnwjdI6CC4unyBKBV0iTcwN+RygABbh7rmGW2LSXq3kg
lu6XJoJQGs149ln9Nb0+0Q2t2L74rMz6AjUDGlL9aEaZnHiUbSSC8KCV7eZUZ+Gx
/tC/nYNBHQxs2WmsgyW3Q61r9T5jvYLPFNFxhXphvVBuyw2zQEFI1+RLppPxiXAE
4olXF9QXS2y91zNG0DH5SdU/5h5kd2jBY87AQv1xLLYhGTH2mt/yRfjLDGUp4pc5
rlMNDQ1mTe8WVfLbJ/E3QTbY1Llr277JoNNytl3W1L6xY27+ZlLmdZ7zihBOgxJ4
1rjxiripMkRlJhYfz2vKI0j0HajFbaKi+f5PYefk8Pv9u3fm7frpAJG8cqBUm72W
pmG41tSvsBt31WgFnDAWgTHmaDNd7+xED5RXFirQSRZ1l76gA40dFvUPyI9g1ptK
TQhsXp09bWRCu3Q6+sU8oSRIuHbpiEj8xf+dG2+9F8El/dQcWJnuerXZ8sUi4uxs
GEsp96T7u56CBgFENLr0VQDwzjfJiMdoi4kx/nGfzu/JVB59E8a1NO10cSOtaCof
bA0bHJJT0Gjo+ZzmxhH7baqLvEoGVudrsxuSBmZqLTd1Lv2/+pby9fSLqmnkcO6z
1YevqYqtYHePgYpcVnFZuQoDwuInDxt0bYOH+nhOFfk1BKCnpQ5IVs1+M1PSy+WF
Z6bPhTDeiuudfB69ahce9VXch4hcPc4fDbI4NzYGiwYCyQ+RHBK0bd5+rh4sCbpF
uPsUHzHavewH41snCpjCO+ExPaSde/QUYL4JUDVkVkhh0G4zEFow/EbirK+W1dwz
hlTy0CW/TvSxL+p2TEz5NnBWqCCkEMRsjQ9sBcrcBGXqvPbwcLyJldpHOopXYNTu
kmokGn2JWqL6IHYJH2vLUDW/9OoDnKSEfKQTKAJ9dDWUJ2ojYsNRZv9t4boTlkn9
MucAqCYlnQ1HP6LHuG+kvlYjjw9bStVtVTSE8BCVRiE7Qqtnnir9rvG8XivzbpBJ
Mw9k3SizpCWxJyOeMgKeJs0prPJvVdT/GsRsTjY+jXTREfNBz1deMy33JLAud8Rr
kD/6Tn9R3QH3kdI04iNj6P8T3ryj7r7H9mVtimzHm/cGklQkcd8xw714YagBnuCc
+Rn352dx4N5cbwFIADm4H3sJWZbfLGjaJBDoMC+eqIDdjLPsaN3cJCZBVM1ibCc1
8fCcvf+9fhum8dqJF63wpjcWk9QvYoqkX7qYE004uB5irrNZ6ewbzT66i7yRepQx
8KtYNCasHuwT+Pfg9yTnHRajRmF2Urp9OC4S1PyGoaNjfpVKTIrzytyzkVQJoeVj
USKvkJDlczjD9d28dvHQ4Tg96oigYARWeIkpOwBaHCU0y2dn8voZt66lqn+AEQVI
Gqn+uZenb5j73Y1Bn+haxlxl87iKEC9IXmwnAWWM7XA4RAJPWcbmUHllm5AudN3U
o9bnGFYhDl3VY9pOf8oEe92tpp1fnV6bFgrPId0oEObvqU3xv5zq4hcG2yFRoBr3
LJFfusAles1jpLyX8PIZwgvVBS/FKUFt4DBRTUY+lcbJpJXk373cKiuvP7PZPGPs
G0i+zxWc3zLQu6c5h6KE9NHS6pslEpBw8E+QuxWShSLFnxqtLf0IHyndApLhuFkL
yWLwPtNSdKh7+lRaKvmmjiFL1Mf1IZtG/PqwnXQaYvO+uI7LMXk6Bh0fSTFD0kIi
M0FrbZ6JaAmzx1snK+UFRktmsFrhtOX3oIDE7ZuEnYeFmzDLIZGVd8osdpOulBxM
dGimknB1R/peMechUb3AVv7GpbM+a9+Jh9rxTeq59vKZHptJWlocRWCYmDo5QrL9
AGISIH3uk3vMnKS6ENAvWBsKFqXhTyJn/tREg8W+vSKEqypLihBwQsrpcmsw4iX3
Naf6x28pNNTXR2XsB9ieUbGiwZeqcma0bt0njLl5d7lNIhA6a+NWp7PT8m5HFmdQ
AYRvHUnsGoXPAhBRjhjMyVLTaMXS5rwbf8ZdU58gLutYIAUQAOSOk93c0ZQM8H/X
enDXltMA7HoB+CRG4XbThkzByLPQ8QCJIDQ6LItfS0fVVAW9Usz/toSAQ5ED5LTQ
RZQVaESp/WibbV0YMbH05gIsHLnVSnurjRACqfRwdBCBovos+1O0mlvkVTpzWA8H
SQnA2/GApYMULywJuARDE+AuPLOxDjwR/GS6JG3tViJsM9YycCOtKb4yrZmtysHI
I8g8+Yn6ydwdSw3R6Q18LpCrp7NbMLiEQEwuMscXwUrXrmBkiXgQPy0+CZv2OP+Q
ZueYA8PfRZ/2B2bM8E+QI2agR2lnuNpi3RU/YlroCokCLufrVwc9FeJ9W6+I89i9
ZHVIeEy5r+5Kt9ENB0jGN8RQcokb7ABwlC75goLE6wwbFe/KV48Dt25yHLyQpVEq
JoVi1ZzAjfIcJBxo2FjQE8QSldRf7WxkgKIX31UB+GRMtbUZHLTiE/t7gOqeaIhZ
hiFGcLHJp1/G2iKG+rO4M8b6eMVeRw+SveS9mYLxM+fs73FcguZxcDWcgIDtAMgR
Q+l5/qpmyNKrL5dlPSM1JxHeMzLZSJiq+TQ5dqXzR4oMZnm0+7Syz9GxilR8XUKC
PfMYYLnVrmO9QbQ99eu4LSrtzDzhEX2jOh+5c/9EKWXvZ6rorGAmWONohgWd45OP
GC3RynTfM8NBF5RTaZ7mmsmq3K20ei6+ExryxHdE2YTY7GRRz6tkT+qWz0CWadky
Vfr9Mvm8ny5+1J3PlRK/jRuI+RbQVoHWqGYvL8epCHEKosnR5NFWUotoSVRsbgaD
Nxl9LqSXkNuv/EeMr4JGNhCkGoGUp3ozrNJgEoHECSYN+GyKL2JIOXfUExEGZvJW
46kfmXJY6Y8aHZTWzC1XWkY3a3EGtgiCzQbH9XVCZ170okRXhXLrjNgAak+y2sbo
dLSwb//AWGZHuT01+v3izdgA6h92sIVUO3xHkHZVZzYXByH+7HphuGc4j102nbk3
xFIbt5G/ogI1iwMVoqcPXgo+o2FxtlvPnzi4mwAnFmximLVJ+g33GtEy/BWBobYs
GjyQBp9VORJoVfUYbgYpAEeeHcmS8A4iLBNdYDNL7V6kuRBXdNnZ1Qk/G2jC+Yom
l/pPFWF/Ixr1afLqJg4E3QQA1Qvu07MbDxkPeYgL1HOkE65md78ccMm5MK8biGVv
qyR7JkyPnDmJrAIcy5Kr4Uh4DAaFhGfwNxjgi2MC++liTnIN+BTMNKRAncnNdZlc
H5iZFnVmog41XCJMDOT9cz1elFnby3wPBRgw4pNmeL4fRwGQZMIFq/TUEw8ajDUi
mPXTJJuNpQmosScSy/8YBXThRMpwyPToV3OB60FxipTn1phGL/KI3AdE+nWN7A6s
8wL9oQjOziQGjXnytO73aKmg/XVh1TSs4DL50rQRZhzL3UsQRw/M90LMJo8u24ZC
Q8EwGH+QziluCVe39hA27pWY1FjjgvLQRBtoszzqtgxygRzTqTTVb/ojO5usKn6E
MSXvq8AcI5mO/j2gfIFLKhojqyeoF8bydx6jQxgPXqS/G6bm82UAwPzPyCF4bwuH
pfCU+AIUzYT2KRNN3RPhjUCFLsvFWMDZc8439Xk6PF8cQPxscgYUX1aofzAv5dU9
I5czURKc89JKYJbhprbYbQq0PvII8WsnYR7dnw3+mnw2WFfgi7/xUaTRdUpIkZcZ
L8SqhLnVPAbFk8iAKZA5E3eGvquK7YlQAbtAXzIN0x0uNobYmpD5WBuCNZzjO5q5
17jyDR5AlbBdozPehKv1Cu3aby/kNLm/pdDlMIbzPXlp1+FJq5XeedvvQ3isZuF4
ml5pLSV/uPSUurRdakHOULb3VJs+URMKG45njbMkW8sJ8lRsOCxBHy9Nokgc7FDd
gsmYqiDfBd0//5FEXIeRLaWSpiamGqaXBHUkOO6b247yy8HLNclP/DgPEjnc6b2p
m/7iKHchllfmAL1hWm1mU1ho0+lAJVKYS21emBNp3CPSc0Zy7CDBM20G0EB+gUBK
sk4/W2Sh/sXH1hH7g8rN5Sm3zao9+Oi1iioq668x4I5CHhPDPPvJFEhcx4xrED8e
XZ8HG2SM++iTNaVq3zGySskhhqBTKa9ftjWrM0LwJOD7qxtjKav02SvZLqXGx2Ft
tp862I18+EdvPb+Wf0CY0G8ahTj4WKpPzurgf9of+rDqfTc31Cfm1pJZw/sXtfBF
NoNNsbdbaf9uo6n5FK0NeSQ+FP/NSRqJ+F5Q20NVAZvt8IyXekHi98lnFuffW0Li
+hdgtZ7eacPGKDMsTfng9Z/eU004cFjb0XgyPQlWrSe/iMdZkqGyiOIW8PH8fKyE
s+B0F1PBeYraAOALP1GgC1Aihmlo93wPExXBjDxYNffElwDPeuegooko3gAnU1xl
zuMoa13Sm+YjiR2v9yQBqGLtarSkiAKWSdG5cILPZhiU1PoGA965IM5WZHjc7WFI
nmtilTTiJ/RhmwOlTs9ZrLaK4N+5J/rEHRkyreM0JxahpNjyDsWKtdWwugBw5kh2
fVbROtXvppkiHi+/Mhxt8lPbRKA5DNylsClqbj0V2fqLr+/ZGvgFnsm4HxFNMO9y
jo5nKEafZfrbMJGq3Cz+zCWWNeIwqpfiTanGGIDkuQpVdNSAbnbi2ThrmSEfy4As
dNGJNUtSjNzg8ECjgEY4vyNn1wnj6Pq7nUQ0Ot1PB3gSPA8GrdyOTZvOSNgFPZ2o
cPwfBtZLcndoH7SVpseXFNXPm4oLPki9wIjNDrqWuXOZN4TEcjB1zAMEn9io8Xi/
sz1qxYGPhpdbfyzAoNBbG+n0DJ8xcuO7sqfU3bMBGmSghSiDCBxUUQxEoyDvXWMv
8tYm9ogGra5sOpt4b7LJUbr49L3u74M/AI0YI+XVtYTCU8zWsAfgcZCBqnlWMdl3
pEskB3fn/lrtlbyrR+aYR34K1LSp9bvCs0u1QNqRDuthHKuYo6d9M5Dm5KgeDCwx
I57S+OLYPZPGyc09D7w9k+x7gE9sD9MWKmdjlBfClPsACNpgF82K6D3pSCOQIPaO
auxYcyFMeKAeAtgfA4/KC1+Z8sCQC+YMcrs9fPOFLnb7QEI8BrOpJUhFb7mT9Ujl
V5GfZdkMxhS2MMyzfE8PiWwlxDGrcc8hHRUKg08QzL7x+6VxTtmJzdXma4Kz5eBQ
JmgSxyoxpSRM3wqr6jPYCZ3klQFxi18DhIczbGLCj694JGE3b6V8kbRNKgglNLFW
LVAkae+4dq/VCSICrG6r1UL4j6pTDvOLUaV+y8IzVGPsDK4zobamGzRnZFdKAlXC
LgpfYcI9xCTD3pHmZqg7QfNTLVDgzf4T4iBcWGp9NsliDefQYuHhhzG9KrMqsUDm
ySCpHeNw6H9+x2qO9aNwbMqpMLKxay9r1qnMui95rxEjKNX27OPcabJuBDq/otHr
igew2k1ZAPuCKgXDD/p8Zv4BvwNflvrkeNXkJQtUzf8d2i6zQUFI1fQdUDqMZyq4
rAL71O2IhsRWP48jysjdYAJe5PgIojXpYSgxtthVfjVqqwJoH4ojYZ4GYoM1sON2
VP6hx55Hp9hHYZF0OoNX0fDPCArVkFSoz+9lFXH427yXOefe55qlX8W7ubkXNdgA
WSoLknuhp0fhSzCO1BoM7fUobRrBOzliuFmQpydutmqNi8I0RlHGdVFb1bYfcDyA
5AuXfrKCAYfgMKrXXtHibTx/Ez14fb0Xfav6VRJ/hl4sXd/e1URhqjvaaYEkPtT/
VEgalwBH6/H34OYwjAoH0DtOKk81X/bxU1rGEcCs/RLYxGLaAuov9D/9XbMKk+hD
/ULG+wyrwYjt7sZ6ShAjRvJTS//wLE7Uy26tlpjKKmzWsoEyixkj6DHJOvea94GS
KCyX2+PjReDfzqdaeSBUcaNIHF9ZujNFTG3lqG7IhcAq3X62uL9gY7+5EZbQythU
NZyNPup8c9ohjwUnV2oVZ7gDnu8qNBAFdKxyUF813NWRys1R+i3MmrHD2WeCsY7N
q4nmqOHN6y/LqtKGAm6bo1Ym1TNfH11kUA2iBtAr/ehATyXVdCLIdLzT+ly1wUvf
k68Wtx9A8jCKxBEvL85Mz4ni5IIkKjD03NpMzMp7+HbUzD38VzMO0OvwGVI8lZ4V
tO8dH3XUlY1SFHm1Mve47Yi2YWldMdgcauAEdc3Ws5XPTLsASlvbvlFds6Qda073
bus7WqxYTwcRkEDHGklxt8Kf30NAOO0uSy0fT9QNuWWUBF+ubGdv2yBpWCkCY0m4
3lPURN8PfUL3rzO+t1WKrBGTDP59cgIQbA21N25eV4bB7fmmLpsgoQmh3DJV6pSz
nZXZRtHNzFyeLWmffZBy35hoxsIkl9q7Fm+J4WRhZy5+bS7eKhqE6relVi8i+kZX
Gj/LPx2QlezqHpvbfAX+Dx1pBTeUUiDb6quPy1meokQ5GbV5ZySOlDZqHTdkv4J6
uxDa1XnzjsBNyFTzReRYLwxfbaZuhgnWPnQpJqLwSZmRwtL/QaW5mi20vT0aAv06
XL2FuiQufgOzQINtnRihI+qRC1mL0RiEPXpnHR/eDR6Jz6FIURVG2vZ70SsWhHM7
jA67uhilSICoP/0/eFD/uoonHrCO3pb3fzvgIfAl5zPali9vpz8BYvOELaJmq4yW
0lUBGxuFhABKI+h9Iy4dsn3BWzPIJt3CEoKpUvHRZVOuJlrUPRIrNmrMPJSzvjoB
LEfvuP2xh2+qrtZX9cf+LyOMJuQvEPEZrlpyEvHPfhtsVCg07GU2mLOPQ/aUAwnb
7HTtmeak5y7DVeqpjwmTktnd8K5HVC8LsZOmUEIrIp0RRK3ZHiUvVCEwVCYOR1ll
e33+BPpmeo6SyiKmMp5N+ooKJy5zRKJxhkQNJMa6a5F3q4CxGklRlvBud0V1XCtm
fO0DnV1jKoa+1mYa2M5QnuuLLy+4qyvMY5sg72dWd2kav23pntzzyuUUrhs6MZvh
AAbmTquxwtIeoikbGxRbmOAkm8enahRndEl6grPxsipdzXRdYMKAvM5qFmHTqDKW
4SHEk7qyy27hThyQ0a7+sfG48Q6sSKC7c+pfGIKSsSv56NmQBg1Xl3Y+OOehsbyr
fTzteH5OQF0NjVkhY8oljuClZ4vvInashyVdrTjlFNc9rRuLoFLfbFfASZg/nlhZ
56pMmN5ZnqXKa0lvNjSELS7mUzIGvKKrK2owswJxQa4SzTa1vXEAPCNdk+UiFJ+X
HemnvwUuW/YPG66M0eH1mz8jQhgSxo7ca/sYyfsc0P3GQRpuUnxkk2zK/DiWCW0w
fbMFVUqj6zI21kbKsayw2bcxqn4sXKTE0bot6NuS8lHB9Az4LMDItaPaqxIJKcY4
hR0Ts4unhCyFaAKNihLW+Jl0m0SXHq09xJb98MI3VQVdZqnMfU/MDL9mAPkC9y+m
CT4efwzIZo+2oEevsL6pExCNCxkHUd3JK7OlIUr9UvLxOao3YEP4zB1gy8taTMW9
P3QySO5sLd7R84P1oIVnqWqxNDeyGFawUReHA9wB6QlxQjlhJlLLbmR8kNCzAe4g
LZfulnUtGVBQfmuRLpsTLrNqCsrYh0NkPl+6/7GKZISg35tPCCkUoOaBnq5ankp0
xsPNsvdCdvyloNYIUAYx/Gom4QxL2tbumbJT5fCF9JcUgkN0sSqBHQZHXBYClSCX
lrgWBwv5rZgKYjSbAEU2eRPh1kZObkHYmAfrBuyvZEu+TKNWK8TdwpKh54pqXKMa
jRgVD2erTAdW0mK6SXs2EYK2FVEp14wFNyl5OhgXtfz2Ox/F0QZTDvcD8dQyM7y/
X4GM8ubzuw7DFUiQLrCuQWmJJDzb2J1o02mzZz2aaK0NbmRie34t50LzXFYDkZod
Q8KJxaiKJttNNYa86WYm7YlkEiyQZk3wBWwkaCnVjtEKlKt+vHTyE700mPYKwafb
reddbZEyYqIYMtJifLd7MwYR3rQ7zH7smOneckrSpQWuswNEcowbH/Rn/6aG7pxo
MCsrPmXX3deBU650jHgoEx9vXxDpe1qOyz8dhjfUNT2nomDMPMlXW+kgYQUdR0aZ
75xLhnE0SYU+ZXHejOcf5SjjWP7T67g3n6RQV6VAgumbugWMjXtXFblx+OSE8vP2
j2LIU8ER2EnJgEuE+TFMBmLWwvnOkgglysxHOInLLgjOniotGBkTDuFavH+Cw1Dl
VGznODjNOJJSd+qanlXEZuRskzGDJKUh30mLm8r2yL0f8Y24z2ByiNx5Nohrjj/w
mq1kHEwK16LFp+CtoUTRbvxbuOLICa3yla5oLr2qdLfagR+HgD5mW3NLSW59ODbI
pvZ13Jn6MSVN2qDzSyAcQnEvR/tndXKUVfzhYq/9yioik6RWmFHFp86q2ySCctJ4
K175+Wmtt6H1jocwz8zJv9Mva9hHkVHZUpN4s4DSLD4bsWZ+kQ4oHg5IeWElGvaD
s9dKnb2Bw9LdfdzRAgroiuOf4FEERI05mgqhhxtTw/lj7IcDFmPjbiq69kho3XmY
nNPVVO4okzNqOPa1lJC8GKx3yZlNY5uMQDLg3gQiKUvwJniBB86kD5XCnghnrP7p
kNxRACsFtZzCq9Ar+d+Vz3RkZuIdSVrNS2pSJJIdj3arIase54agO1c0qST++Lgx
NjVVpn2lLCt5PIwJb8MBq21qPiydN6WtrUwk6E3echPVcV779Br8P+tesN6LBFzh
YFXlC1nDwa/z/w594fd0u4GKfnaZ0NDZc6OCYucpzdqirbsWbuvq0LlF5Z0/F03g
DHcm1A+8gh9lEXFTeRr98javpz1ubfaWjrIr6oX4uz3aVS2ET8y0mKpGsLG7C14h
40wvVhwwDLaT9QdHKtX4od7Qd3ZWKwAvZLUpBMsNRRd7+bxGbra/6sbrn2rZ+6Uw
/x604rQOUE5EhIoZ6dIbO5mOpe71EdfTXYXmf7aih1TTXjySHaCwWuu7nYy86bWT
ja9PynP3KdOR431djQitoj2ZUurJ8igXU9TgJkWNW37TXJiWkHvQnSDiSYo2Ic1R
VuFFafm8zuOQ+l9tcY0iegLii87nURVK2gTso5ZPBkr3dBkvmi9YbACT+HU2gcjI
pCVlbgfFgYs4Eo+tRxt80IUFiluFOYT9/vgliRafkV6PTcS4lWygDO5Z8und4r0I
shgxtbI4AoezNpHCyuJ+ZeVNDNqV82IMMN8KOLcQTuM+BjpwzwRCYY9MRB14wfE9
ajILFj8o1Kvg91eD5+uIEXV7ALcoVXcYQ3iJmAjNR4bxHVGyo9hVsRWgbHRnJbGD
c0pg8SDVSdDqxdGl08lwWD0WBUhmInlLHmjc45EwHtLI8isqKNptigPTAFzTT8Hi
xLXQ7yFiGOleyh2D7AyulR86DlnBaoHh8NzkxhGy86dydV2rnc0dP03MvN2tbNvZ
M/piRs7oHxO8h4/iwM2BKNRfj996QpUaiPJL025rupnHgCTbKzPOcdU/of8ot4Zj
Zl1eFSqkFh5DHbJOiGAVjSi9u8QDnnXlzSjO02hw4ioMsGxiN2+p5KrkyhiIcZJ1
q+kW6wuLBxQZHLnlrQEbEd5IVY3rVYRmnoQbltc8gs8IuiPq/aShgd80ZUV1xqfQ
GG7ctWSQLf92sDYJPuQ/YawTM3/Ic0eVcpj/hWK1MR099iRphf6PzdyAklND4G7R
vbsYnHc9rpkMyVx81/RPhFmLY4e8JFVwsNIu5Bl8/nCZMRa/uZrVILTZaOYPRg+2
qkR6yAAPnQYGqLdDTh9AkMkNeuYuFpylcT+Qr7qZ7Z0vtBQ9vMefaGXrJYaSE3Ba
yh5Bx79g3XnyTnyRN9osPcCy7aorKWx/N925P9BtlOxWnbAA9IVsx3h9qj+SbRri
joiTArIFRyROP+kAzUvTsHWxAcif33rFBuFUnIvUxilkinF8lwGTyamRkAxiQAbt
KKpI57mCsEjisjnnTP9pW/ocaCkN4u896XOIW5nH3Vs/seh9zp5LszCLzPsN33MG
UmNiSF88MxoSrCc3W6vHabSIAQYNzdmqFmrdbeSs+kkXS6/eRHPSP+ooT1nRS2Jc
mpapltBdSDfjhh0F0cj4psrWzEtT++OPx/kHGVj1nsqKpQGqYv906AlObsfXSxQL
/f/5DZY7nezWTQsQue6MWb8Y599znXoD3GIdUqlDB+NjEoiPCq6lXZiHi6l96E3n
kL6/0l+UmJj0xXCDgtyx/1apPJXFsIiEUxlmNr1zK8dPDzNIRrIEZorHQ0ZMg3AV
Qqx4Hq1OLrJTx6rjK0JAcobMBH5A/24c2ca27bnbilW4XFy84Ze5MIlmVoAyeCMr
8gxknaboc9loBJMXdOikVNoxsyPxf4nNIn0aZ+MVhAi2YAxTlnw2hnqL1gti1FUi
BCchz5s75qw+rUXsya11q6h/mD1IwLxOVZVaAeYlndbBhhVgV9P8fvQaNSgcua5m
pemdgLkqne8m+e90hjobOT7M3dfxnfAEXD6paU3wGVcoydmnZ19+KJ6Zghx/edDH
xHYlg5rAWdBk3dk2FtX9POuFWmuwJe2ZLHy+j02nHlfdNtpuYJo6uUDC3UeGse0B
hbAXevWRrnnaJcvr76lJzfznQJP5MHUrzdnH0N3VBMMYobLmDTZum5NekNiQjfgV
ExoOqTcSQa//Pe7ucaoc1TVEP062ZcbbuXun2ysJ/2k9VpvOBOl3NaqGG2UO1dAZ
5bEyyzRFlJzNxkeDFzCGtvIV2GtzOc8I04zZz1Xt6UuDnCvJGtBOnUs6csDXiMfg
NEXDKtn1UJmXZk9nx5ftmxKeB923S/JRhTupfQ4Dk7+lvPb8NZwnENTqStGENWWp
CYu/wLJSlBGULCdZIx6J/D4NRzIIjimzkjAvv7PPAeTLS6i8eqtYo7k9MPJaOwrb
b/4c/vzaEU/Si+alC78o3uq35+eKdX3/E8RZdsBwTQTaSgsRukZuXqxN9SeovgBc
e+LSVFAat9O8h2xM3eRU1Zo+6UqDTGoNY5w4mk2ukLkvVYpI1b4DdsoXpqf6lY+L
cLvrisLo2zgwzF9OdeZceU03ly1IChM3w/OB+MjwbMMtTtUhjHgSuNuKqeIlpaSS
Vkq/05yCPuGP9HxuwGtM/efRkcpX+9onAcabbHf2HXdSWZwWA/8RFSlnSTkiGzP8
1pOqIHphQ6ntPklVzDR84Bfl6FiBuwNbX1kuoO359q0UQphBhlFLqqebzmRzMF7E
9fjuaw5/Y55hwPv38Fg1QgyvXsx9BO1v28oDqpOmFgQb29iE8B8+I7INrnYHvzQu
KxHgfZjCFDUX9DsviLSNn/nflFdA01msXMd4zkAho/PGr8DML0SmKgpNrmd19VGP
M3pl4+lOxT7xk8mcF6/0Anvw+XKZqTpfa3rq7OTYfthwAYTrGKmfvgtkiVK89Nzc
QWoqO/E0JI2eu+tRcU6uVFyJn6N8SHdko2hsSR9ASJdA1+Wo7Ngv0F7hYXv191Jq
vYw+1cYV37uGAOYnXTC9AzjfRXA6h3KI8IxYi3q9QplEGKAGkF/S5ccE+cPc+GNM
2MLRfP3eIpytM3tyx4ESaxuArv3MuBFajeKOZN1U3OXUakKen+PlQlRQdIJ1bzqm
bn5oX0Gv+NtO+/IYdBDPMvmAyGNqs0Mx5J2i8GLve6HPsukBaI/lLPESkau13t03
4uJf8HeMJnED2EEiMOma4gM5G3945pF7NGb3FxW7SiKieY5iKNOtwYa+DuOtdS0x
7zcJwnbZqF5Vccx9qQo6KQlsDqjowCfNjIUoROc38Wt9xAt6+G9Lv5oHAxa6BNVA
nzQmRhzQzSdTUVW9BH6VZvZNsA8i7gKjwOVQ99skp3XdYTgxmxFWkEY+6q4BQxpA
El5fmU8EN07EHSXHe9zVU0CGJmBkaMJqVVn51bBKhsuahLAK+2inPiPLhj3Lz3yL
dJfd2jmxHqp7rinSlUJUS/wZlkXzwbVOH7HEnIw8z722EZGuE+1smjc6CZ7OU6BE
fwlHp6DyUS5I5mx3Erg2z+HGUQCNX0iJr5p+JwaeLnkkeuD5Z6uQrmhpr7keRajy
T6bYw/VH+lLl53vL7k+1f72CHZaIPw6aZCh3GVHAOr12XZdNjgXdRIQSqwwGp/nk
UDrKoBOyuQIshv3AusE/C6KMnMASwXIgNK7G19Ca6eoUiR4pyIRMCdAZu7pQ/xPk
mJqtKb5YQuxYmJzC2YXS376pnuG/aUAsYafG4BWWKLaqnx/3BgW6phPfpXG+eykH
x4hcEw7acTY0MsK/DN9zoSGuQ3/9fJOPYaj50q0Y0/ipzMCInwB3/NeP9ld5o7aN
DoGk+/KpIAzj260wUJvjjGgwxlr4N8lJzL42IqgMpCrvhPsu3szw3rLlxk3NMvLe
yEDFMcbNlHQvNvXMXrEPr7nupvHkXlH81XFa/dwqAky+TgsaAq+jepqR9aH1/Wwl
jniXhJj/rsayw0dg9LwHAAekHjz5aUdrr93MT8DLXQNd2uCuUHP0eRGWDwLvNTgf
hHefxJGaP6eNPa46/WMcel9pocir2Ypjeiv/laPNOBiFdvCeK6o6phCST8Jl3ZdA
KxqNmd6CPxUbIfjT1Eh3QulxHJWdzx7nVVKxa7ZysqATWj0nuhYf7MAIVNFfHiN6
cke9Cjp774vdvTSuIs/jAG+3Y8tOA7SRpqGEV1LfBfh4Dyf4mATXtFPFVKLZHDi2
aRIsItqZ+yQvU2LMzodnF7zuzbJOVMn2B+9Egx04DMeqnfaMMXrKjtKOPkZfsado
LSQMSWFEmSL6z+SUsWeLhQSmfyjGEzjUem/rIg9GH4OQDqV8ABgXsy7JvBBOSG7+
lO1xFYoIdtFe2JUNTCmStlS6foT0VwjqJL87RGaie5+D+vnjYL+vUekRIxB+AcHh
RcJoSFLZddE4NwuU8dfUPrv13TZUi0xpD7L6YrlTw2ZLrsr8e8Pzh8/NsbmJiBsP
n0ZHHh3/SHf1r0r02bUudR//SmgAttQnkUIJbRDzwUUJxExDunjUhum9qQ+eyLEd
qI4KGDRJkKP+/iEnCAh+jJa7LNSeoRmSEIEF03QHGWxG5COnXSoKVnkX3cQDAQuC
M8eCX6CkS2xiXJfegMKMDqKM+5jzLBI84ZJ8RbMdN42OI7EKK/z6ZzvZVx0s9hZe
JWMvtbphnaA+FvbsGLEOMuFd37mOAUSuIXUeyRz9UxDN3ZCp/KQYHJv1lk4FAjWR
+gpkpkEfD8N6bwcHcii2SnfX+xQmFR2oxhcxT9xa2VHOVDuT5bEsWgXDz/YG2HV4
RrXQIkUtsQc+1yg+CS8nf6qxLpYRdHH36zoUJMDp+0Bd7fyuTRvCRuybFDwuXeoe
EV1n1b6aoLvFXhdAwOPSBZALyxEPPjqAdGDW+hcfdI5A0Srfurs4CogETC2S/JRG
O5Fmk1Dszcu2sEsgwCh2d2XepymjKXxE04nnu6z18hwC/gF1QAKvUiVNCJWbIFwi
XZvLC6IXQ7FjyqyH9Qea61LIFXSCMY5Da6t1tn+HPnp149ohHea1XKyk3ouznAL4
bWIQdW/JOQxZP8PbSvLVPYhs37ICT0ofBo21+Zx3NbYuo4m4zewAVdfc/9vvZoS3
Gww2hQmCmilCihvfK5XsOJeoMNqsqSKJQ3U/2l8H2dzhuIECByON/EHGUqRnay9P
xVKwjsDYOD2t0yR8ipURi1AijRk8M1v1VBsMyL/egrSg/Y2ijgOZRUgwNkVxj4l7
VLiOWUKiOIcf318P57KXiIhbRF6dYRUXSNZTKQcf9BLIKWNWO3kCfrM7hUIb2Njh
qUUp4LZLEB3pyuvB8ikU3XfTuaWIJvfRF0jCi37uBvvmcqqkJHsst+o/9C1CRAzk
P+prMJFll2i1WL2kkFgRWLs5ktR747XidzxnuqfzOkp9lepLmY/IVomjAdY1E1bP
aLh1iNCF42y6hAhOYO22PDcYHUQg9Y5ODLLqiPVvbd2Mr8w07aTYvoAe+n484cxm
uzGjxjsjY67QS9QtYpsMZ2ZbuuxVGlueRnbz1HDvpb66WSpY/3qrne3PCMLruqoB
5XG3JCkhpbeirprH44wY/5roJZhdIAbJa1fXdj3IRVsYEjipbIqspfpu1d851FDy
6qq9OaUsqT3o0P/9X9oJLIWuuurPT2a/z5w1W6INBEmGUQmWT+UJgRwps/GIHGI1
yO76Z/iJqURFG1b89xiNOM3VjwdbEACkOZ4JHICKU5W8pzWIPMYx2aXF6ufE5f8w
41DFMg5Oq7GzZKtSSQZlZMFRUW8Vaq7q9/41o25/p8PQo9O2jJF8/oSeojt+KPQ0
JThh/ysAu8gYUfPdLX+J78WNXjjXsFwDjNSbkr0IwjPLOZ5UAvGSrjzt3r7VWjAb
neKaVp+B8GuRpnL47b2OG7b8Fgfflb+y5febNfgHy7Pwv/IQzL/RWBxatNpbFf10
YUu835p9xy9sXoL1mF+pLAN3ZQdRNViFhsXGDfbH/In2DF2nBMLvTSMsdkxj3uim
6a2jqE4xWjZCuygirxS7NuN3CevfCiM6Wv2R/dTulgiBqbmempkgXxw+JmA11i/2
NjyXxWkUW1Ndm12oHX1/Sd5LWlqxfp/k9muN1WODOcMYx/IW1hN06YlH6nvF+fQ1
PyE99vSMbjcL8dR4XOzAkwcxxp3UkCtpcFwyPvZTY4bm4ZOm7QJxzrH6c4MnlRMd
cY7aIL8xCc4DwFFbbm1DD2sbsPGYzqyPgCNmL1ZaXNLkNjrPmMOzcoKwDnWOk6Y2
Tmp9ntzzHRBE058OejTqE0nFOxMXfWpHAYvduNQeGKLowKNKkWIqMvorQLxfsWxN
243kg2RezHm1c68F9pKd7NWlAMCaOmw1/K7OOq+/LeuOoOw/mrkuuZRNqJ7dV9aJ
Eqjf2H3u259vScK4X1k3Uo2btX/GrU5W5z1tmYXCQrOQkUJQpecgVTyUGn4bGb7w
0i/zGCJPdxWsN4Zc18D0yoECYca0EaRb10zZquhEVymCFNxzOL1x1XwEmVz7SaL7
tTH1h44CtobiWDSHXPbbTQxLYkGOPJXRrzhxi0fa6Woo9UCfi8JMB41h+YHybpbs
iuLXUAYJlgTLvy1ZbcMmLwWcQa46MxRihkU81k7nR5TvHy99VyHTL72H1qcFcd3L
53LZ6EyYoXc52VKEZUhhMA5te92/We2LIvQiLveVekkajASzHARHsviunVbYGGPW
W5dyQH2o98srEmPdfKtoY9BKbpN77J+tjYIORYIA0Jqj0zwjdN1jigkONgvro55P
cF2EWWMpWf9L1dcKZyJ4quROArcDfEbCTWovNLzN69mQW6QCCWXxQvxvPv+MJnFq
1RlrUu+9LX5Id7gxjk3gyySB9+LySLvtmDYgebWSwK8pFXC64ZfKsxzlcWvRHVGZ
U5+I9AjOgMgEoktx0al9Fb71Ge5GfG+1IMutIfAH4zYQK8PXBzYI1Pj2tv+voR81
yqZL2FUaiqYNH79V3OvqsyhKcAkVOOajkt4fw/vSEnhUiaQfYwf2GJTFxnYMc+7D
QiREtZr08xvBNDEnjmNsdZZuUzsxMYVezmpsAoI/NLEKI7Sx7VdIZY2Wyk/Q8SRv
s7r/8X2Oz4r13mdMZdxogK4rexCWQh5vMx5arTAphKvx0vHNFXI01cVw1ZyafUrd
roW2m4tCWDWPZmd57nxIMTcH5gUKLn8ShTa2Jn5SRPxS6E3Gci3UpJ4qMVLws0q4
lYWim4kM4cjd+hv6Ib2rx5VeM1BekYb6tnfZ745VpQ/IEngE69W9A8Dj68tRLbX1
efOQ83u088Tyo2RtJvyeOrSi7FqmOo3ykNQBpLiYRNdu0Jcq+I4sb/wwXmRq7Zl0
ZzLpu4jwVvFYFG3MQTWDTmd/OUSW1ayF+z7ws56dxFKRabgqQhNhumOVMHYEcHVK
4/VdsSCnHBfogfBiGgbLa8jLh9qlpdhwCErZ8CRC9I5PvoPQ99aNCWMwbe3tPSVj
Fe3PaX7/+Kl+ZaQTlyfDXmcTQ2/dKVPrlruuVw2tdL5n0ijQ67o+hU+htfxTAaMu
pAdGWGRqz8khJhgij6L+D/DZrSeWUB6nJJl2jcri+iyo1WRs4lMB7SU3G6fOGHNK
qTzLvZbNcYCBykIx8PXOqrqDbUZ/pzW0IGayJT3x3c6TR9JiVGP7I8mXg61sxF7N
QQjzXdqGsLoO7cwAkV+iZ1LB4NWZCgllucpnu0whTyH75w7solymU0DtTO4x50b+
oWnNyb3OvOFu9n6d4SGYZt+PuL6Nz53OXoXBJ2e2+gw5iXBbjBWsEOwx6R+36qP1
5U9mg19gC8RkdDIO5uYE9ElcZUJh8N6c4mJfKYpMTsFShpmNC3F4apP+K2UsJmJE
Qggjh9nKznMlGBRBE2Agj4dIeN1tHiJ4BHfIVql6fgh0+fJGKxkUJ+gGEsYdrrt3
P64thQTkhxQXJwJ0K/UzLKOnc5lKEHt33VeFaYqOfJclZPZ1Vx+2ZUDXsgDpNjs2
S8VDtBJ+pf3FyCvvkGpJkd/9P+vhZHutIlfoLAJ2HfiRsySaGNPjNKgoCMp/DCn+
Bsor57H1kJUu1AX833+MYdtvORZKnaoW4mPsei+r0m3wKG1Tzfi2FEk+/TAuHju9
sHmG4FyI5ICskjg+PA5lZjy/k0fU0DE/uQyMiLw2rnUVnxS7e+tUpGvboOhugumW
QHG8kmDZyV8h9fvjOuAKgDsRHN7zsZsVirvCo2LuCs3RbgV/Q3vRYItMkK7mn/On
sDFl5zfSKO9agNmOHtLvOd/FYpy8r3+Z7ZnWgN+bO4zKYv3ubfchHo5/lamGANJ/
6NI2HFXlq0uYczAfzPwPILOiEgahM2wrnb2zXSmvRzvZ5UQY0iPFjnlMqkEfw5Vj
X/OeDlbFtxrOQzbjcLCmWXG+Ibh0ypggnBiCS6XUNqpcpCyaiwrE1iULWv30hFJz
p/GTAXAwSKgQuYAL30+Y+GIOpyghpuNdc9rMcWmojtGTa4+XEorGjmLMUg0ga73h
YEOWKniXN8UQf71G0Yep613vOFL9dTZPLduEbjhNPzKmzJCOng/VM2ekk9JsGaYQ
wjQo0WaSmzY9S9fmlHzcq/l4cTt5ylCG7WRyjVuA4qNazdUVuEJb7z2vD6M0pVdH
h4O/rtGMUJYkKh//FaL32VsA546V6PgEIpFqm0VUJCis2cuAb/a8BHdFMN4FAFn1
ctlVxPJy+NTcMz9F5LvjQrSN3sTs0zYiwAaUOS+NfHfoMljT+8BZqvvLFRPf+lqv
mFXiCdwZKRWu6HFEgvXo7MV1g9RG1Pua8nXBFlF9Wva+Z0iJ5IWus+OKroIFxKHv
x5UiHetbscFNvyz6GTZpfKX9LAC1EyLZTys7gQz2SwQugKpU+ZaXXYtTw8VaHEXU
k8qVITTCFc3OXwPh+W3wyE38fokb9L6fotGPTfA13egxr4Lb5kCMrsrhiSmsIAF7
XDAY9Q5QlfFpJruiJMtY1wzfA1gkWkSJiIRY8z9ttwijrWQM+pG5Dr8ByTYu7/PR
lJd76EVq4TNPuv1EkgKInX5Zac35yl/znT1jPWctbIxWtrQgQPHpdWmisIGF7tr6
VOz3DARtTL4I8Y75HWRP0bAU/WBDGKq+R3m+vn9KgAxguLw1ANqtciQNmr9w8Dss
GCJLt5/JntWjsMMhWZambu52eEayFt6hRNvQBPshOs4NRuyOWNcyco8yWIPtgpEn
qCSMOdEFmuc5qG2IddhkXamkRbbbBoRa1lqv0CI53kLvpUNRUkykg1pAVUAxAq5p
pUAToeZP3I/HJyOau3Z+BbDIGK18S2Ds8FWdrgGK4eWlH+XvOsZDyynosu+OM6wX
nFBSGPDzPMh2gKsDISaLjn7IYI8wmC1VAS8P6YJCCtDsT7OK7qnFoA4yhqi2OQoW
Ak7ysmLF5mBbce0gHlZcsln/k+scOr2LPtU5pTQmne/iAiwMO49Wq65NoX5dV0iy
0nxDp0GUIdk9Ugi196loMEx7DyYiI5w7e9H0hLxN2/oC1JVjF3O8at8dwXqNt+9C
VS2KTs7FSGQn8T9QuDiolP1RgZQX/SzapTezLxlalJhNp81OLsIEVW0PErkASYS6
1oUwTFM0pd05e6CNmdID/wK//ds0cZ2ZqL4ZxYyu9OvYSpyZF2kr/sQ7hRKwWccW
F8MApDMZNtdItwwZPM8XJ+xNtu4fFJfz4zemGSzYFnX5mqxaroRQSRY3McPsp1w/
LsH1TQZE2TQKa8aMi7ypoQZA8HoCtqRVDG3U/p/kcQljpBFHHvu0VMPtmhyNWu21
68LxFlJ1osJHzJBE2XYShRo0hLJWI6w1dhGOba4hXGfD/Gfh/mNbrD5cNko1vocL
cmqHM9EA4BX3Lie3AlQWqKCvvv10otPDuSWixknd+MhTtebDNRyjNT4Q1YvSkvUZ
lLwPCRD2QARZIoTKqAN7JhdqOhSuvw8rZKTEh3TmekukTdK3xg+FflYN4RHDB6r3
3c2M8u7CiZViVroI2WcoH0JAnwgp8jqSbLNqK2/JzH/Rg2LiZOpNlra+f6vmZDUW
DvHAWPeCQDCZ5ORM5FY4BYdmDIXW7xJyAEJwkP08+7xygZuqqMkhDLHFQTdZrEJE
RwlnqiRgJHJo8quHp+3JFAKvp2RFlMacclaz5BE84n18rPEN8cM6DjtbR9sdm3zK
ravncWsiddUBiueRPj+xDo9M50O4O5yuOX9yrdmNBdRxfTsmey9NTFrfAtIfjQHq
3la9k+U7KgbsmsjIfL5rpcTtqlcJzHRasHnYJRKwYeA3+ctGfstxeqwrbejaxdbA
sHKAkYwGF99LTlw9Jrq8z9PwzaWFXcbF1BIIJ2qs8Q/tLc4YrxWbSvujXZyoEL6/
OmEG/Wh1tNt8vgpuXQs1cVvn/tSDcnylMmsZLoaI+Jwqa53FefGRXJJpRwGWH9e+
W3mUE8of8xG62+jmvF1tDazhISBQABu5UU2NTmY7vC+Tbcz55g8baqBJE8cV0K+4
seuo8uFdKGSOPYZkDeFZofrZOy2gB7EEWIAbJGjYGxqeFU1lyK8sIGhjK99yUFam
SMcmPXtiNx0qCNQEomUZTb9ix99EOExqEcIY8Ibnez6Z1MmNJ9nj/+gXB5ilGFEt
hZGy3dvudIpGoUNoFruZws9SnLrNf0FtN2aW0odRS108Q1J/h9xO/bkG+QW1dfFz
wxWtJB+QhjiIB9diijLKREasf/USP2XFNHCTQOFSrlZ9ABUOWSQot6zC2IySWd+Q
dBqIDwQzlt23Warqkt4Ms0tjLvMXhkqBWabPwGHuhZ22V/WnfCAPfcC1z3MLZKbh
yJEd65zgZXGM6i8s6sjgIaSoXMct8WW9jm9XvdQa1NCASDd/eg2JmQLJFtPyLYM4
k+jNZjUFXBqhnlho5PcIxRpv+menBQQRId4kV+GBoTSBjZvGq/JVigkA2Tk1CiNG
a+90F0C2XbGIDxkfAiSEomTUC0abJtvAGP3HAuS6x+gFzUmUsjj8Js/qByyQ7hJT
Tg6IeOzvaycTvs1DxEAh/SDMBHgORxLLCrTuGShdzMOi3pxkqdmySK+J8n8DQ517
MdfhG2XYjR0yIWafNxz+Gy8UcpGVsqGYD9Z4Nf9IhXtgbtVDdUGIuSpNhroF+MmH
40aPBs+Vfm1JDNx8nti3HMN92XbDZ9OxgacpLlj4gvsrLkqlHiUcJnf5/vIH8BBs
qWlaMk1zjzHgq4LcWRvgyjkAGSPnZ8RfuX5qOWJOlc0RY0faQWuRUKFITKCaD3gh
ndCeF0k1+rq7Su/RAQLWKz1jQ24KdXVetHMpLM98npTHjqTS1kguNxX+IvU4lM/b
t1PdhqLQu7uliRwHA+P7GTDsRLXe+WHlslDYIu9LXAb9tyCAWqkdVD9AwAgsGpbi
Mlo4LWLR1EMSymxbwP2jIVfe/eJKCRYA98n40j6oI/wqCHZxoi0ao8Bc7VRFFDny
us36SrZh7tTl0ZwPiViOlN6YOD3kSbIMwWB/LVusmY3mjN/H02tXWIXwd0qm5XDP
n1N5aNjdwbUwCYpUavJQWPrgQAantu2/TOwLijCFrrCZIBxY4MJuJVXOxwg+tuKF
0Is+7Q/6Ngf16EKoJn1DllMh0VxU47Cl0NMcbL+AhSb+xuv5x9HkUc+qenbGJQO4
OHvFXaLFoIQ5PevmkO8A/uoFjuaex61mUO3+pPh+7tTGq6hShYqp3OTx6S/kVupU
8gShZMdWw3l6XdWBgMpfMtYH9JR0GKrvpCzB2JAYM2I+rQ2UQIDWpu7ggI3yc5Z1
SrwIOtJZxEU2izyKGNM2DCSBSclkvoAfVZIuVIVfB9Kx8Q5V9P6dKAdg+2SJIoGn
4k5+3SU+DOo1OllW/pZr4Ur6lNIZ4r6SDqq0eLuBLWZiRfRY/XyrrLJmY1aoRooG
as7Qhv57153IzL3aCCH4rvtpMCKqR+W7WJ3FRUV157GNHHT3SnxEBfkKXKmodiBd
foZlGyGwcIj0RDbP92VP9aF5Pd7oY+Sodu4nD2jk4U2PwE9itjnv0uB5IUNjUrri
LYzF0aGlFyYoex3lxfHUieucxDTbp2EFo1J7ki9DZ7Kypz1ju2TMc3oEEky0BkFF
b57GCw7xeJ6MROiSDR02kXPbHb7er+EIBahl80QdOCFK9kWnmGl8SGNNg7iC94Mr
9//kKRaH75tuPR6IpxQFqxfw0+3qyjFublMwEpEiP9v9/rM4EZndgPqdPZvffdOT
wnH0FLchTe4LUGABv/xDZmcEANDUhceueurcfOsLJ4QmLUwOm8TQ+mHuPMKq4eYB
05hBRM0GivcJeXG98csd9ZRbmAG9t5xsRrwHQhoOpYN+D5JwS1tsrC6j5SoyNgvV
2vZFdNYnzAjFZ7kgE6v7PPPBhIKUFtFwZEHEJ/eW3Yslt205LEXeY67CHb4FQZTZ
UDfXy3PNu61YfXLvwKmWZtUwkFgQIzcAo/FfIylMyrD4Jp5bFjVOX3GAtUWfNYkS
fGd43ckyuSBoSdX2QeK5cQn30m8Cq3a8R0Txw2IO5OV6+botjeEEiW96RpLB7xbJ
8b9B7C4X1OyuCv62O0BleWqh3YsfRsKDbbvMZsVbvyQpS2D7oRgV5T26jn38q2Rt
axmh18TDLhAsexI6/rOvp9r7A5pwJDAs/VmKx2+6d5PHAZcbJfkERybMWUXGdck3
XzDZ9FwyS25YoLull7rzpRwJ8gw7Z/i+aNg3Knolwcc0uoEmnG8dwsaQbIl4aSz6
er13q+747fCuqz+mZq7xz3/wXsMcj32liUUhE+B3zQPTPpz068NaXuC+ehdYeNPe
/ht/D3nZCsU/qgJtqkrQ5N4EPlqCyOVujYqoiFAt43vkyZMwGBaGO/LUFBpxZ9WI
13DOx3Vcyy5T2IFD5MqT1IxUbTKlIzFxX+r2X81mLi0XJfAKbg9Y5gP7Tvvg++Js
C9Kn7bTSXoUmhkYw0r3giqQfWoKqsafMo6eFev09ny8d5jT+sv0YhF+O+OtZaUGS
dU4nuWD8LPMALf4ITYZaYdXiv3e1Zeohw2+d5N2jmsM3z/dzqlaIEOQu8s6ivwiT
yaZRtmj36GF2u+0KfeQt4Vy1iqF7uHxyiwppGAv97crsz1aRLk83QWlDVkWNQzIo
z5+v7LcWvnTpAbK9WOx+1I4ao1J67LWD0hRARkON+ItbQdiUmR2KfFy3K1e00w0R
kH12W1dORJBhMA1Wyl2ZEaLLwo0tIbqrxRFBENJOwam61gY+KbJ3SfrdLVobfltu
cl/3C06ctnORPWhw+3ysC7bQcza9xJ6vPhoHLrjX7vvgomML+z6GkLtObdCBwG39
N/sz6WThUJzA9PaCmrIjuOsrMkjB386Iyg77vf9gKHlfV04pAFfjJF38lNGLBmDK
wicC8xgakKyjSZxOCZFl0GoBbDv53BL436xLi0q5DfUjDdX4R0tJdme9GB8FYvM5
2Qz+BucyprhS+T1d/nQkxnOGEuzu0E9f22eEwqsHNKFO0WmMgHSFWh79mB3tzBNE
Z3pM82XO72FYhntDpmkSDrI/hHSojgmKjqaLWKwTAT7IlLNtbQrd6f7hj2hgpoCh
Bi2fgDH+ofa90BJSBkjzlaPH0Tv6lMFZDb/IariAPWM/TtDaMTkc5tXj6d85a2Sp
gAyg7gB5A5n0M2h7m+8ZRJhvC1iSXGz8dYufF+/B8nRAu0wzVLt8764pCfiIE08k
C5j8PqvCBbSpsHb6EI41lwQtSQWG4p6tYdYHbaUlWCFXDzGLoaDP7C7Q2yLODV8j
EcABtzlxl52GVwaJc8Ch2wzQeCMS7nuKI72IbuxcXKwh3hqee3399YsDwTKFreE6
/YnK4mjb2pZseWqFIAsUfRqpQ/o6tGtncxaGCFIis5GYqVgHumPIdgPLjRlrmzqx
yfvkIZmkorOXp75Et0QsSzs1pZQ0tBKwTpTOKiw8lOl6BYB06swH22ouki5FNnZG
QJeiWcUfUWUtKTS27WF3hj839mcS9USVlbOJv++PaFUnHlU2OrD8UX3/Gtk62JZ4
`protect end_protected