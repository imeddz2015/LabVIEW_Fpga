`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 13200 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/9huKRhRMtvnNqb3Z+UU7TahEoHV+T8U3P3ufru7l1O
3DlgtZzb9QxCbOjthp9+wDkjygH0eUfDrEl1ovhZG63ucioC90uCGu546rUHpZD+
+iII7dDxywvpNSezQmjV1pe/qm9z8BbtW+AtKKJUMPVNMKd/dNvdjH9sbxngHpeQ
D1vV7eWwLtqxw8UWlmq8QVxzyVsn2FEIHPOZjUrSmLccWhPq693jba8Cg57sMAzf
s97Lb6CcysWnnBdq9iqiz346HgsnxmQeTQwlI2zUGoq6v8slBLYt/8jSDtkhpAly
gohaI9n/4D3HGAw2hfsF+8KhngqDBGog2mIlFa0JSrmTeLsVE9+3/ety3QheYf7Z
O3JT+MFP0Vy7w/7W7XEia66yX0NAJMWiAasFH+OHZkJfruwoCbgGgRccA4qP0lFG
8DMdirIRjfSNUvz1iXarjy+M1MKSfu+T4qW94yUxA4eI60I8fOh3Suw/ZZRFeAsP
inat3EeVuQI+C9qXI6jTzfLaPJI3myQ3xoAN+u1xI2jZDdwN2u2zHg6q7WQ0t6fM
ViqPmua+ORHnBV0oasMtOurJeLPOfmSi2XHgzDXEPxSsx3J2tyLeZlNcs3oBIbMT
IN3EcVtel+KVTCjRcWWbAk2vLudIKhz7gdpr7Tsa4BZnJjj4Wh48JIyNHu6d4O1L
ABft+SBmb1RhdMvWL/meiAVrlLTUKXQfLWGu6lN7+j4/5pK1cLD7iQu8ZMM2YaRf
RMoFgebAEWOXYIG7OjMSRkn1lRhxBQSZPvhmoc5ZfnYyuYjXYbrwi4ePdEe2zS0P
ZvNIOSNxClpH1k6gmNe7h8tXIODHXDE0tj/OijGq19slpi1pUaeezgYbOtRXWyVb
euh7LcA1rx5Q8EIu3wVVfq5Kb8vBzpB9g0xhOgpNwmlxeovjvmZ/ySAJxF3t8P9W
FUMPWOBxK5RBD/gRYjvtfL7ANwdJOOXgzt6cfypYZRVxSmZDjQsv5JS+sTFaBaVw
gFsFsh3o0VojQAWl8kc08Wv2jvDnWN9s2PAobQ4yOWMf0uc9qtqMUvbpYBUpFP3a
7EVLMxraPuyBhEkiCLJ4oRNJGMOhrPOG2Y0Pt9+Sd7KMK5iThEGzcPGXRClkngMq
QDc/3RSLbkRRI6P63pqogoXOdExcOto+qx/JNHo9vZq1+Wv3hqbWLP6JMSGZ2Iv5
gDWa2Qg1U1aGOUMeI0KhPR8lZ2huoC5BzCCWpCdVFxs4lCmp8qjGjFagiHzjSNbq
LXFy/ek3HjfBOn+xTySNjKrEW70Ufh4gj9NZeheJ7PWLmlNXBgrwib8OhsoHQSRp
83h+9ANHRBl80ZKp1YW6xHk1G9QHsvH8KUKi29cWapmeogJfyeVXvpSmn/bd/Sxm
+NaK1zrIDZvh1WUHc7pn/FjB+qi2X+xzEjN3R3++ZffFb4g8PGe9SiXczDujcTMQ
dalhUEj6ri7eOAvIadZqniu1o6CUbrguw160YXnwfRDyaC1EtmeF+3VmgPjctwMq
NEC5HPyNRn/fplZxsqjpVQ8t87YTUQ/kZdXk4x4d2LhcDT5mtIXj9Fp98KaypKBT
ZZz3L8z8ap1vc4nVOSVEqs0eVOws61Pu0jNuXCjQjby+mR0bpElGqMQ1j864EdNE
u1wKBWfeaxbqHtKTNE853FyiSBLtJVLZJbUAIdFCAKjT1E2kM865Fhe/iOjL9wxt
EjF3QvgzWYpHTGvAbPOfOXTD77Nk6DLgYBEOSGGWqmSCfsIFFt0yipbi2fOl0Qn9
iYGCUW75wSG2zJ0i/7o/+D7lfm9LsYhfpKWy1PTM1QqHAjNH3bxKdaeWNxmV9e22
3YKjeYxHvlfVNILwXk8ghKz+oEPvP7MvMtZRBeExewQnRm705pvU228gg20Pj+nh
ForCjxWuJKxLkFuFl3ixx+980OgA58cVMkq9UFsVCh6hAVN1c5DOqyIRM7bBRc5n
sezI7m3AP4lTXPFEBVrnMKPyVNe4nlGK2zpcBr8qSS89wXexNONUOp7bh5Df5ALR
KokOO04goR6X+4dVJCJPE186zXAaOysozr+j5/9jJWepcWlgZCyIjeY20YDSBgVT
BC7qC+/Yj9FN+FM7FWcbjHNXvGHTEMTtGxfBAjbkeEUXhF7uglfONPIpN7T5pXYt
POD35xFc8bimUN9XrpOAdA7t/loJ6TejRow5NHIsEnwtcKlyw34luA9bITN1IKVZ
OYHSB3C8HcolO89EC9eutQP+J1SlYuIxV+43LyvchxQhXrjYOQZzg/nuEKJMcQJX
ybHTrSRya8ciXm+FpKJ7U1tIVoLl9mUjG8E2pLGxd4fqjOrNAD9xawNf/wpBVs8+
t9DRreKeNqJU3yQLb6TeUMrZlbDYaxBwiAtiWV4fwuTcF9sQRSSB9xDVKH2wR3w/
y/mS5Cq4DzmbPop1joPxWooO6obqe00/qfszl3n/PZhLMcfbBHQxZvjyq6ekfZDs
9s7iP+R7rR3KbSWrMEe7XbwJTcACfkKqU1c2gaI1SG28puJGgAjrr1gs6C6JkYJv
0uMR3KDmqes0JquJCQ8Ah0iksBIRggqxd2GMygGVCHf2XK7D8o3Uu9wfPtUeURY7
e4KbJ0NxalasBKwqNy03DY8lbJldjWWvouWNk6mZJLER/vOL7T0emqnD9AUJFhnp
c5uX/vsk7aoE12scqqknkWtc/JTfe1xHlGE4Mvp2CmEHntrA4UwRSmCnVrnxaXUu
dGq/IRX1uDhkKlzTKOTP+m4SL0DX8Cfug1fMG0eWNwrDjk+bsIF+8JowH00xz6U+
2dkuSXd3Hv66LI4B+4wBWqVC2r9eusWvUp/bggPesTvsvfBialIYsdZH/6a/VWU3
1/ZakX8naN3P3sbkIuqE5Zuy0vxQ7wYohkeAyoEeCR5+K6q/7PsQ4BbwWkTVdVF9
48Igs0maG5MNuSYdL1in6tg6JEAWt0kfWvTEqCpasHZa8bQGHJS6iCcV7syBmHLs
ztv2IVk6GzleP+JhJUlU8VE4cgKf1wmMQCVCIVBpAnwkzi/m5E6+WpX8XmwsQ7ib
vIK8Fnxj/gfndzG04bRWs8G7e/QqNybm5wxPwIA7hRNkZoIIMZcfidGiRqDhw7I9
p2P+qQX8exXHF8aqS6YMjgyy4248jFUWk3YuHvyhd4oRkBEwoMIsCa90nqM7dm/P
sCxw2+5DLxgBnZmBTCjbjpB8aP+9Xh4D9TgkVT7gN4P5if9glEGK9Sg5qSAIdll5
4lunhdN+P3jGLpBgBFNkoE1LIHoFo1dIIkLHNTZH0qFSBEVAz5A7Lw6LFi5xLpnZ
sDkzCQLmV7DV1m+Lo7ke4/QNa0QUlzudYorGd/2EwlCq0RC615KxdPNlPKRwnyF7
nvvrgwV/yQgN8uKsLcVhczZkZfaO4KlLx2cMihXfS5jqzOVC7j1GBCW5CvARPUib
umArYQMn2RMgJB7i5pYXO0XXUyaGvK2iUqR0QZ+9++Cu5N680PmvIotVAD1Kf4eU
f9aOfsVsIp6nqaLp8P7j61S93VzYJKN84uQT6U+rMHYwBeI8lVQcK/E1svQ8qDg2
NYyokpC0RpgyejieJlGeYziTbfUgUMwvbHVDLOr8qFMQOE2yB4+mPjRQAUU6H/iW
k8K35Gej19Jp9KgoJABkFW1Y5zi6/ai9t0xe0HvyxWmzRluGV5JpAcxhq5boqPFu
yZF09DuZNiCFy2rTuqL716ZwWfRnT/NGYmCJTajAG0ox34CbvbtareF8r9Z1d3HG
9IpSziJixGMxDtbVzJ1NLHu+2sAR37pTvMmBXJ+YQeG0oQjXULdWPOO3LtFjFkoU
mtROvPj48JCykYX+3lYH8vOB3G9KdSGL75+wJADk6tS20P4uFZAPk9iqUamX+Csl
h2nj+BcxpBlD4n+8xkoeP5q+B/hV9Tt9LR/JexksbXeWhj5xajLEOGDdqNPhvDKg
3voDWeINnDZRrOXcfwRPngp4Ce2iCNj18NQcAYWtam4h0h9dtxic3kVeUsESpu8O
0YBEHqfOl39qbwU2nRnTRm3xaojgHS//t992Z90FEvC3i1EaxhkBu7Zn3qXca7pU
vc/fgp/2XWnRxS2CrEjXgSkF0Emuj1aWQ+8uoTm2/mYLRYrl3oVoTDfjRueC4i2o
M3f2eZSAE15GPRoN9ipa2oDm9R+xJ1ysDFlrh+AZiA/ZJOfR/PknLbb7wsmrvCZe
bGIbh/EOz4qA/Ac47HX4XisEuvJbJ5TeFL+H3zdgK1PQVv53Pi6+H6BBpYIStm8v
/oytHeiB7DNxDKqXxvQeqpueENiR7W2NEwgEKS/5cmW9m3BLiPOJuvPeN1x8AHul
0mm34WpvokM6VI95g4Pt3D+D43OU1p810ZGqnBjhQ9IYFNpUe7DUB5beUuUkgpmz
PAWq2fo6VkvDzKOFnum4sqnULXVQxUTr/63840i4GWotvg3FCmL4IKNJoChRWWH4
Mi/oqQE0e7zn83LN1iE4Mu1jnBzzjISI26h2XVHlDqmOVDcflM6Rpf5J5pqqbNTJ
2S1DUwQY7oQ81ml2ZQOgrKuQ2gecsSWk4Q5Kbs7vtRgGw3fOSsSK6AOOSMNT4lGP
24mWm6jVV3o/EC1Z7UCVb1mdKR85qAucZj1a6o0pJiFVAwYCskQZ9X07ReFI8VBE
dV1cQ2r3yOsYtSj7pZusqZwS2PXU7lXwUVrQyEdYAG6GTPZnfp142k7QfUdUrYJj
9R4x7JUngkg5vHQ6pZnvFNkM0QlMadMoR/wj2j8mmIM8Jh86XwDpCJKLCl7XqCQ8
8nRFT/BWxW5g0LwuvQEelvk2J3rLs9PstupPtz4VtPbAXnbaT15Nkyy/UOqG/cKu
RBV45qc+VzG6ogNInccV0qjmKoC47+vzKi9yEKX1K837on4eWawKoYo4hrxxhlsk
sG2UX9QHzLicWPTLLo0X2rZEOAIsyxIQWcG7tdULdxN4Hf9+PNdOPlGSxqXuoIxD
mi3APYzKVvHFKFWVNnl6c225TTHvqn8eHsgSyUCT3y36w+tIo9rpKfRLiTL6bHSg
yrPo+ouw7dtsXZ3ZYd2cl6WUmyNnGgGcd8gp0ZDZgfhHg0wDNijwexCb033eqdl2
+mEYOSxzEa4QfGa+6J1Cz+jfe581jkqDTu9WiV1eG4T7jJkkDvvhhk9kq6UQ8geZ
eD9atoYuywEmntW2WJrtRL6zKcDYkHpJnR8x7xh4MkYErQWtWZZPWsOXi/TQlq2p
EfMiMr9rNJKPUS+4Vtcvr6T0WvWWvY8V41fmD/rc1GEq6kRuX/DnCOKWvyMLlP/Z
nDVhMtgmXWny7xkj6UupSo2ysNP2//Zof1pYbwcNFllAwy03Iw7oFdd53szr0gkq
/AyorNT3RA/L1BJ/4PfAum9ucU5btwpLBd6GXhFEJHq/sPnjHd+QtC3a1VhYStJn
G7pK7dPkdLv83fsqLY22TM8T24aAFVYiX8oYt3fJS4LamODfk4gAWR7a/dM/PqEG
Yk/zcVZHQOkxEiWLQESy75btwR19fm3Lo3eXf0RsLpQRFzgwyZ44MlJXIVxvVLP+
+bkI5Gy2X7DBL6HWwhUyZchtu2QmBIJgT2n1S9ZX81+1GYEHX7HzUmhz7UJV9BWX
KqDUmbkwZOyE3C3HOVBxy+KV0/je76xMNbMlHZWuocJ/7PeGNSOJPUhCS00v+4CJ
7JahCLxkyTtIKrRJ0r8FEs4SGn54lgMIgT7FVXNaTc6uTi1S/y7JviOHLfh+Dre0
cWOXCWCMzeNLly4kHGFXtbfXEPoERqW4NnuIkp5M/FD6LwIEeocb/CS7YzJlbfwg
Je28Q7saVXUO89OEsJJkB+wlgJ2b5kSOIlyeO7dl5dSo/i9upGiHtHqAFFvJDmhW
NhBPLFvq6l9g6I8wdOVYcw8FqAfiGqQF2fstbjRx7XU50+kr3AXlcTRnw7Nx6OGN
zIpr1i5TboiAcgkt7fuOLOietc7UEpZhkf91yEI0y4ahs4pt2UtDA7/rJzieiL/8
n0m/O0PYHuYjvHMCyfSiWjtxflzY7rur4kdjPZvUbepH7RjHOx4E+26XPu4YRoXl
i0Q8/OWL1z9d0mDHA9bbm8tObAdG/1NBh8+nXQw4xn07c67vB77HOcbvU1oDCkKM
HiywN8rwJ3nnwkR+mFsKCQcGV5IPN09/43fxJS8MKs+EiEA5YSeLeNMKxYXqJ6/s
l14+1ifK9MJiA2lcFKfshg359EGkLg4TpiAqZ2LphfhFCFEV1kn+aEAD/GuzDbBD
57MnJ52iJCC8vnP2IfGhJOO1XDGg7wNg/hPhJV4xF6rAgxeQf+mjqEODD9UebK+L
C8Fu846RvXgTv1vuxJWOvnKrpYcYOU6UDeQCyD8DW4zrwPSB9qx7XgE13ZnpFGZr
4xrlg6NrQr3iXpe7+TEQrsEziAyiSJnN6E7wTFe/zXu5HtFQ1yfP9FpCP/zY68zj
nR66dUlrsGAVhBZg+xmPL3hKN+OeD3TCyRzZ+v2Hg/Sz/8ldcF34Zm9CfdZ3aK+7
hbvBCzxW4yDo4Skhsx0yqG+E29B8dDdjk1f5OW1mWnSYZxPAeBhrd5wXO7jCyE3F
DyKqXFvIF2GXJVmn2y54sgd9LXR45rpj8/Lx+yKl9NGKIpKlMwa1NVmm5rEdQX5s
iFRLb5uiZy9WBah8WSyicDjiV37TXjUSg+hakccOdXuuRYat6jZGOGhW6LH7a5Rt
pjAmgCkdrsMq7Rdv4u5MGSJYRFb9yAVhc+7ORPPyHHMQnzvsRUXQOYsBfS1d2sOI
EESedVgLt3wbRSVjvKrSFel1bIiGDSlgdxSwg3pXyz1alY7DT8nb6sbKKMclrpm2
MWWmR9SQ9QoOFgNN3Y1YgufrAGCAYNo3hFDuPaz0Y0eb5tdu9TZq1U9nxhYDBN2z
HREkUJKjZ3fK6SGqwzeMW7w1CCW/LhnroNWJwGAkT6L0X1g938Xd9mhj/twa5Hgv
xdNMWX99xUIajhKy+kaBrwJS52EdFnz7m34bkGXpEFmJyDwbLPLJC/5sSVXJv39D
ZUAcyWnei/fJ1oNz6b6mWGUml+Z1dDnZcNSb3TGEjgZhwn0InSI77ue0wLONXk9b
mmNF89lj2bdQ6a9HC30I1s745jJ9fbeQPn0NZZuibGQK+yqi///2ph6z5pngj94k
1NJBs0wBpZK2IkTTIKuve63NH7HkDrrJwrOmLCVLHFXTKXcSNS5hqjIoAIhOQxkP
kfx/hKr8hN3zQz92v82iyx4rsoiqvNdEN78Isa3+dXqOMPNX3PWPk/97KWDPIOdR
pwHErzBazvgYWwjd977rfy/r3f3tZElZ7IlUqy8aMwien7m6VelPEzRxtRBYim1z
1VI4LBti7AnOJ6/TNO2YWUrJ0bxH70KijawMsDXxyyzL7ev6vbLNp05h2eSazOra
ML9iMc8qbZ9yzjFkTYJ/0Z4Sq0NW6kJ0aG2/IUJ3lwpIPuH7iKCS+nAr2UhOpqCc
QU3cRwEOEANMKC4mqtlDgrLn94MqkBh7Lt80/n5ZT75ZqBQ9vg0sQhfZ2/H8MMrV
Y8Ht3fhPVsQ1Zvm/e54T0cg4bWtx8hbMSWI7FsPRY8R11Amodi7lPEYnnySAIWhT
hKr21bb734lH+XvfhPO65ICGkY/sYSjd30dgHsxxsyJEw5SJPfy5q9cjegulkB3q
3MJDiruwvQXD/sniCUvUfoc+umaeiPat2vB8oybtudlpN8zvC0JY+XHLWmKRDZFZ
CQ1hZ/GVJYmwOoS4fluRuHi+uWxIxG+XC2ywcJsTsSEZLKrNIbRYvJdZYd77GQEh
j7vTdenk4Y1rybxOAoLAQuOwbyodjtJszSDIzSLFWDLl+u5aBYPHUykvk9Jy8HnA
ncjEbY9jtevJcOhLbHttNBZWL39llZYg/IFn4AE5i/1nhG5lfPD0BT5RzTe8mv1S
jxJG8gp2SN8XsLhEM3Xz8pjXCAS9aYbcEVadnNlAYemVjFLJdVW/JiwfYcSmakkc
vpzdb7wFe6fDH7H9oWUSsgiGWWJGdinBe1PqtqQP7vigvfl3ZVT9hXMjpR3KcbQ1
OiG9QTJJM0IUVsohE+n3cuysP+UFUdL5KkwhATUzL4DC/FHt+ekhwDQbPyg8ExnR
kPlKvkx+OZ69PjqHt3S0HVr6J1OoGcTJtNE1Eh2sq9hbjeS0eHW8l6W/0f8hIHmq
NUGbSjmwpHLZmhgDBvLTpcyGtjm9Vg6XyZWprnObMtXCc3Hg68BZlVw2KyBntDb/
eXgC1GG9B3jVsKZXBIO5uqVBeUkZunIGHDgVQaoR8+b+gt/1S0Ia06fzzBDIw+5C
urVUa1RMRUIK6B7c/t1G/bGaGElJHwLgDmRDI1d48wmpRUA+gd/WDynKPAil3LTx
XGcDpi9IYkJD98K8M7KxgMUMRLFDW2cxQwMPzW9n57lstqMivC+mppSYrW+t7sx+
e3za8tLRPMO2uEdH18Jz7ZzqcsVB05yAsSbbKCFGIdKrZWtZqWdcwHbeC9xEpx+e
yNX2KzFF1Uui9xOXw2muYhPqdjjkLZGn9nN6wl9o0t/b49iBwJoNPDDHoNSFwmOu
meVFWbsUPAH5gjcFobDs/TnEdUsw14KGR/1/B9uM1MYNZ+bRhQ8B0czWJwDhg87S
sQMHb5mP4J+NhHbr/bzR+ikaIkkdAB7MdRB0LmoyDgQ6IlPuJBzy5SSSZllQgo6f
WSJ5/8qgqHbQ+L80+mMyJB3fW45+WucsVw6M7KaGFcS2qx4jsKhN22e1W6LYbMlN
35LRH7fQLwbJoOTca+aM9iUjh6ARyAUyne5UGvSXFbfFGUeEJqcz1blzLDQUm0CD
/fhEfUTRPz8fIg9I/D0HgPxj0Feh+uK7xiQidrHQ+FSJUVQ+kG7qe9oLEi6EXByf
LVKfA3DYjxAOGefgPhsImbUPmi6BczcDqacja45/y3c/zWPdcwIfl9KfUr/Jvfz8
eLdxB70ULPJ++MAJ1MSGMPYqqrsFllDCrph44N7ADTBQFyObNZrtvhLFoCYd4G/K
MakZnRmha9JtPW4Tds15cIWTgpc3BRLaxQtSpCyLwQbgiTG2N5yT9l9JupMxuhhX
fAoGIPxXCrt4AdLBi9X45j67sbRpa4UPjYLxPvaSWN1ou73FdcLHxmZ6T+xwFbF4
BL5OREqpAu9F/FZ3E3aP6nwXBe/Gcec6jtaOLZvDj7dEbB3imhckAFNbG2HoN9lX
pkfX2Mk453wiosgVjXUf6aD5vqKOKPtUll44oTzcXCVn0f/OAFpSRoSVEzWcGepO
Ikh7SYvJFBNU8t4auX7+7oXN6xnGiqGrzMJb8W9T1Fp0jV8b23ReZLM7cQfawhA7
TiLj6VLc267r3o3ZLDRNpGW5iEkzvbbTdWZ+XahW2cGkNcQ6FC8PZlxhKGen2VZ+
CCKPmHne8KcZlsU7zTkUEQ8xYoyho7CZhfk+M7OPg1juDNLle1+YXNx3XXBEJKE5
I3p1YoDbgm04iYQIbupOu4UgopbJgoK8AGiUX45BO+UyOLl3PsIGQY1bqfkkw0lY
763d0N+a0TyQj+5r6+qpxd31LnxXerzSvvvLqZgBGceDA5DsA0TiIb0x/Bxurgsd
ypn4iPC1brHehShI8NyD2MSnMht9JINYoOA2Hq9foYXSZex1EtM4XeTXaiXYijsY
XqCWOYBv/VqnBFTWiuynt7YvAzf1ew9/NWF4KOSVvq6VFJVU30eLPa6rC0mmsTZm
oVPteMDIe4srra9a1XOU/FTpONxp4+iHFMcdzUGXt8sHe5Rjl7DkE+ksgxwXrOE7
HTWISfN6UI8RlUilWhvDIk8+CjKlrhuj3zBj2lqZu6jKhmtJsiO0qIxzjt5ht6aC
H5eqYbrzpZZDviHSovDUYXH9vC+vllJlq0SWGBAvzvTZple0YrPqC9hdNMAKDoJo
yeq3Ig6NE0uhc49NpnoU5EKxHqgLQLsz4CqPJb8o3rLUhdW+Jmz75GAoSw2ZMw+G
DyF/n59ySlhhnfiqNBEk4sdnq74FrF04h/228OQ9y/qDSOnOldNlGB6oRnZ/EEV/
kkQc4Y1RqTR7UwCu1/0retb0yOzW6Wwcyjh9mv4nNL2UbPVJpBjaqfkzssFjH+Su
3dkVxKfHUunKi+ZzGWXM1wjBMHtZIy9mJw0b2kXGPVwl/CF/Cl/lEnciF/iAo86q
L6nZXOqIbLv6QHOzUg60W90QBvuXTm5d3gPiHUWT5yo6LNJi+h5fj3ZRkqWXZwNi
UQtxcBid5Fat0FwKqnE+SLgpSjnIRxFaKPmDeMucXzT+B8lQiI3hjv5dSokasmwB
noM4+xijbQZkSCag4Zu9o9Gf0NiiASNIwxxZeKTq7mQWEyTiigbjY3pyjoYgmEOA
Eak2iGlk3bGJIUlNDmueWAUyXr8s0CdU20Ehw7M88pfTfTsQ/bNtfAaEnd0gj4C8
PofGQDVADcpfLXcqS73Vma9mV6abQ8EC7DwCrVxHFmZhUv74heVdZZE1BpQJVlUs
RPlSeSSjzXrG0UmQPO77/dt4qw0sDgzcXJZBZRFXzeMeX1y2F7WcXcvKWkU3u52G
qYGdNfmZq+tcW7AFMQjomPso5cyIhIPgCIRDokqci7Z98egzVD28fyiKZJ4mJSkT
E4ymcz0sy4GxHqIKvsYLcwIICW1osaxhTgaHSC+qME4bNfHzBVVEh/pcfkxCVMa3
BVGbcPmgw2ZAnR1aYTmTugn0eSSYX1XjhWIiuGWRf0DwinQB05PUzTJ7HC6czhiU
p0EoQ1Z0RaKEBmJaBBNPDdQxW/upv6wAwAeUcXrUoBwJTrPw/viIIZ5+sS8pkAJk
OUCzwc0kd0tPiYitI3KZZUgkmmZWhMQS4s6pEVutGMlOYOYrgqAYAYFlCrqaSzpl
OCZ+AV7CADaZ9Ozao+Ve69y1557j084YaTh9/EseNpmE6dnhqK4x6SmOuoHCWejk
CQAwGJD0esqyiMFTr2H9aQELj7KTZyui0WlJCokmctSY5fMYISsH25qoijiHrkb9
xft0MHVw3oz2olTj09AzqsAuHFSDf5O9vniNbk6qdKBFhlB2g69SgpoXKiw/dJ6v
0fC5Isji0MVST2vmQdToh7E0j/LFtFPI8rjK6wopUeM/Tv5LEzwRMrkV+mYar44l
S11H718jk7NUdUI1rsquzXeesQWCZQlRs6a611AHS5XiDmwAdNQn7lGk4iBLA2r9
qbG0QI5SsAaljhXav4FW9lgKgtseJegNZYrq+ncFO5pg3MpPEw1V74iASAaRd+e8
2Nyu1NgYAs8MafvM7SLh2g2vF4mWawVitcTl/xD3mdp4XiDNab3dhnuigrTbaxOs
brma6MnWYNkBLvMlj/VCVZSt2oix2JLoqLqiYgDkcb+PMHfes4pBeIiSoaN/HD3C
sf9kaaPy/C8RgGnbup8mylnq/xtO++lbVYkx9ckHwZ0Vb2Qx/FhD9AzLLNUaKQTi
8Pnl7Dj7bvnzGjBkemeboOVTa1r+saxItvo8kApliq1foR2wKep5J6yBA//CJNJ2
cvK10QbpYNPe3cFm6tK9E7moc4TFz8xplfbYPI6Sgxiw+BpcEqqvgkifq1LGrfLS
i/ce3LnhJMscyEuCnF0v+i9e1ihrrMLDOXWJ5UoZgE3bHAK/N5SstXMcNnTRadKA
ZuSBT7btbsP3aj6/aHxgWOdRS9HkCRO47xLOUYnGUX2eYHygNlQmUoXBqjS4j3Kv
fD1spD67Ap5SHw6Z4UGhjMPZZf0YMA9Q4R4M3k0neq3ulgpq/k1KKdrx8G+Y1xQ2
KFCcD7O/vTlOIgJb/8jJcWJBBTYf7YGPESHeh7i5gYwTW404BFJ6xVAUI1rFctk7
W2nWLOseSfZV+f2bQT1UE27JcPQwCGNrTiD+eDSPc/jMcL8Tl3OOPFVOABZkUBhw
BVor20GA+0+fUL5lHZf2KuLdVo5UVHmY8ap7M2vRpEwcQz/140F3E6XT2f/yLk4j
7umIawPJ7hWWb/plY31+3fuCbe8g88kybEEZmIOuxtUXRwKpXFtuFeKlMMNFyz8S
kY3fOwjz2dXmqzwxRvvyoCFn52AMbSO3rd24ZGEXOzi1a7IjSY8O1ejElZxhrERe
yJEJqKxd9NditMUieIcB9sz36/6nV8BB66knTLsZAdlHdF0SNlZS+j2m7WvU6Pxg
GpS659uCVNRT7iM4lXsAZq2+aDAHknNfny+8BoMc9PLH6DUUVVP/scO5L1bG2kRU
NZZ0ETlc7JWOYQfOc40Fzv8ZcElyqIa9Y8dPpwZOd9i2D2JA8kQCmvCK4BLwJ0P4
D/wiujIGItWWH/YifnE0N3RQwNSj5fuR9ewzlq/MjjKpBtMzQRZqsTVaamkVhg3g
V6bg0vTjJS/RTOdHflr+qz1nx4dpSAJb0qxfbH+6Lvi3P7/uUDuBcOuOy9/QhNKz
DsLmHyclTUQ8LIhrqmo717SfQ7/ib7UUu7qi5dOXitzPIv3m5xJzWwRwVXEPsUf2
1qfdEQWL11LaHxR8Ac9Wudq56G2fTMZ5aJxmDDCOgEw/JkkI+eurD44tzsxoDOK3
owv+sAdPi6OP6EWvrzzPAQgzayD90nJi45N1Umac60e6jwUwCPtRdEMCHuDifKAj
bE4jWaLO9GuY8j7sx5uyPZb7q6iL/846aXts1Ex3IUB8sSeubC4voLMOd9MeuMaW
CDuV/vUck1rkAQwlryWKrIRqgmOrwBqi8v2Qbw22itWvOvSkhWRQgv799hRFE9Wi
defbEoPa8cycibONoNBHiVm+ajhfX45MjS0nUFtfnV5hdO02TeXJrQjdMF5RndU0
a4F+atFRRXLIUI4uNKT6NN1eXrCkhaRdwq2NnkTiTKbTd+rf1t2kOHmpJbvQUh5L
RDxt6OpxycRNTNdooUfVx90D7gUr64ygkUtVHgrS7/J41emC0SETwzD9qtZ4qWsV
nyFdAnT1o2aTY1Bp7GEDJAdjJGGB1wApqf0qYP335xE4Ae7LlZId2iH6tRHQVd9U
Y+HmRB4r8kDtREqz1Zz4FcBbDoCWgyn1deYR79PHXbM5BOoRwEewLf5msNMFHuiM
QnnR/bwLzFBXMcRL3oHuSclQExt8LWy2G+uE/vGJnZ2yljbtOS01J47WojBSbjhY
NHkDsZq6OqrQKH7G+SaKICjq3n5Lb9IeVn5nmdMj7LlVDvhoAxxxLFhng2H68RBr
V0AUW6yYyPawg+plFiRLZV5pWNvSlO0kPpdndwcB8n3CY0dYd3yDMHslUBPjS2J9
LzomPGYrDdLM2RarHDT+4AKRo+7fImw5Z+4PXtsiJHGn4WfHLvpmgdgDs+X2mxQd
qUdnie45qjTl+9Js+MHKP5EmDzMPHQs0J0qRflEIqS40rnR+UGPc00m7IPsH/jBR
Tg7M0mwOWO0AXslcZH4PLyu1p3xWl2zCBiOZbyrQN8VWxFlwulgdZpRllaF86F9d
vfz6nuIzlTn0SRHsVjaISn4+h0/tAAoy+bmc+BkMiObetKK/S8HL555qmDFHXmNy
Z0bouY65JAiSlV/aoHk+5cTnzfEOPlsqTnc7RpDTmsjIQ603U8gk3D251BsSZvxb
fbqoYPm57uGTt5rpSqqzyNvJS7izei3x3/63r2B3/YHKif7N7DwhETChRKx5LRIg
X46+9g99T9q6ufCEFVM64iOF6aj9Lq8/dj14T+Ub4C23Xl846AVlSLewrjyuWXH+
YV+CgVTgADQIpD67A2W7XjrQNf1AFwx1loSOs5LiCau/EFrQj8u/Uc8p+icka3KK
fHR7JftNH6sgz2yPYayaY8rFK8jbBFu9C3raIrFdtRqhqElTNEfCC+qEncpSfPjl
DjzrQO8rVSFbTeqzNy9O/atpeBWU62/ItOLsq9G9VzdkrkR4d8Lg054vLzE+Hk5+
lj65bWIDlSrf/iJ4diIvSS+lP8VLK/S4AnnDMYrbQc+2JymahdSswVjyqAosfHHh
2jk65WexH94BG6nolbs0vbiuuHDv/xLCVlWDN3UwFn0j1I1T+PYQjtA9Q2ALobEF
7QpvRuoIfWnZDrjUVrREzY+YmtffUEdTOt21llJbE6daashuNSS35ZG+N41bLLb7
e5MptwETt9Pp1GQk3T/+oTc0AeqD19sUvDpFap7b6Glezm16KKxhWAqkxV4JTdYa
ie7mCunkYtXT6jy2ekue+Es+SKZztGpqeWJ/bjuqBafQPibQoqOqjGJKR6s3Dgp1
iGKue5SlAvtAvTh8oCSRWhpT62dF8MjCu2Ag0Q6F3O4Z/Q1mrl58turLGHgCnAJ3
DehIfr7eCQwlKRBEXhNfzkXwgk6vk4MoTXWGgGjzVqct1xkVi4tgp0ff4DUs8Gdy
zs5UJgPkgyVcFy3hjiwnMdNRu2YBuYIbFCoTD/AGg3gM/Cgm13+LA2tlnWXGq6TF
zomWGmh7HovVob2ED9sb1WDmjO5P6guzONz8oTS5C2VHu0qV0IhLx3G0uxnGUPx9
se9YIqzyDVJVRQkHStwCH0dveXHPlVzb7WpturExLlXrhq7/31oCwMgE/3c1xnAs
gC/A0LmOUEwlR6CpONxoCvjwTqWDUqFfl5PnFEzEWxGtr6oPeVNHf3I+oGzwjka4
2gs18UYurszjhkRZJYNTbBiOW7gSJbkq6qZ3zBqRAOsYmCfNPJlyJSZsTXNZ7j4y
3El8DzMK6ltONPJCP07pmtbUpKFpTHvwQH4XQxyR7VC+ErvgU/mN3v86tiejuPC6
utpOdCHUB7TP7Qrq4nF/fWqumkc9Ju+AbvWuC0GNZhXT4J/Kh8+gKEdgj0bX0yj4
vGQHpnq352acTjrL0rhgrqNzcEv5+WHGNjcIywo0HrwawCzmfr/vMncvD/KDTPOb
JqmggWduQA3nwsPhjzpoLe8jUOvqEqrUBxKaP0VXZnpkrJxwaTBqWpnd/aPA1sUw
PmZi4DLbhZH4zn9h55LPeht9n+SJKBw+oQ6FNCRaNJgU5OnD3gAkyEg0OaOayL7k
cCt7gsd7iTANEoucQ+rmmaxZi/9THCdoKenKG7t1RkEJHAeccZq6lTIq1Vnv6Swi
Ifjpy6xfSO7R4RzFPb1cgmzwZwolTuak6JHClBx/mseUovSYUwgQGFMkz3tuOLq8
MQcuhw54GeWyvA/nvv4NCCyASc6wHlr6qylyECEgIMZHZj3ia3FMm9D8MFP+Wt23
dAPOTnLKiqCD39yAAIfr/5N00Fqf4c+Cx8XkA/dCSnLmYl8z6sWicn30GB0NmCf6
EJbIMZWi8Bv0jwMpHM3OUZ+JRUDA/f2zYaHTTn9zmLrKgC7vb+aFaYorREEqKk5D
bQ0McbC8efeF1kKBfTnermhRw50ZRnkqp1xDymz4lGgOGRtR3BBoA11/zgbzulnR
Qx7MAyEMQXb3XdBCw1t3ibR65/MZuxENWd1d4ASqsbDFjGKUn2ACjUysnDkj+lF/
GR8D7X4sJ3lNZQqTJ/cshLKf9lQyA/M5CcNJ74xjob0ImIAig/mJkvNA2aCgRgP7
qXJqwkqIJk7Z5uZYUhFgjAJ9j9OkQPogPTw/SfborFkDRexuw5M/XcMuo6blFP/y
BDuHi4Hjy+3qZODhgy+oibU50wdr+HLn9bwubn3dBa24CKoK12ly5siabAqfrNFp
0Gqd5+pLBofGFmIsxPtdW/TZssLtXdUTGAmzjcBdo+93M5jkGOheaw9fp7AUPw/9
X60Fu5+h9BNgEZn6J+xzkfHvXMHonEOI2mZx/O9tGbmBCRJEh1AadzNdonpV2AJJ
DK0mArPSEpxoMecLTbK3kq5xpix8BF7bdUNB8Li7qNOWAF6c11bejQxx6KDCrff3
BjvXnVxXjkEpa/4uMhzwvtsvKiLj5OP1+oYTU3rwGuc60PaYrrCE9v+rCLm+CElL
4ZsQbb5eTMEba548YT6Ygg77FtM6N24JnEZVm2d9xAzyWvSNqRRvmT4EemmceESZ
mBg5EABlo1Nn6/YolcdtXzNai7ghkjIa94Ttz30pWLtztAT7UO6InWNAJTa/IeH6
3s5gtfOgVCrvsATzfL04eWsp+zxnDtdCQoDVT3B+bAE72Sy2vr7QADKbuyn3u6Gf
tlAiLEIFKVVk0N6RVmZbgzQ+s6V4TIYAnWvZ2kWmJ4MIk73k8F6gVJ9YXGfgNwUD
bxaAuigA+NorBMYCxhVXY+3rdeeNIAvEu/8nfyKI/lfQOITG35AJY39X1XrIUEOo
4o/r1/SvSXoxrv+eaYS/oNKQgdXT9pCHmu2ExHwj8BGXYberjrbymEqz4xUoliN2
aJjwSwp9KCY3eNFXIs3LrgBavzWlTwf75iF3+F/dyvUXoH2wauPMMsGTpsXayU0N
09XY9LcdyIg509Lu95laOVqwP4TLmq3JfQmd3kAEQ7f+CRBRrmcbPfTDY/OgUcY1
tnjpdG1AnbdqjdmIFcxh46fUa1c0hnKoniJuhev6ukHvGwzf5OaXnFYB8uShddBK
tSqytdDNCmCogVjgn7y+6HAhQ++ED1vw9uM8f81f53P/G4Agge5bETYZvPcBstdj
xTc79FQHCWw9YsSRo7nWjqe7DVGrXiH5dS3HsFACJYERl24Y/wdyipdPMwQjmMTJ
7no/tcX0UGClDWzsCGgngzHjOdGu/YjbifDUmRx9QfhFB9HhFySfNQbFCyrgUtxE
H2zn+tOOQ+dkA885LPIUNDAgj6Slcxgfeo9ludGVczCTjUFwPBEeF05renIfwdfE
1qLlFUnm63alhdX6RXRt4GvSPcQ+cyBU1GT7TeKg2BC3WlmbxLCgz+BrCqRDcD5U
FPbLgDx2FZC6eS/18zeQKVxJQpUwZhtp3xPmn+kMUbyppWJzBBEx4VYxrrVK8Tru
zken/ejL2SV73HdmTt20fszCGCEiLjtXXMItI5suMgiq85DWKg60wHEDSA+JYEf6
XlaCEx4fXEKCycN7jP4yra484uSe4CSrPFTo5cNanmMe21EdJ4uvLPudCO4BTVgy
0gcMpYyTr1DxyKBAT56vsvdBDOq1yFjenC/1oTel5nOS7zX6ZFGou0KDPjj8aReK
zyauy1AbRVP6ZKUKFolKpuk1Z0yg2pzXerEhjyOWk1ngUeMB6Fz7JFzGU2RVfuCI
9fgbjufpSbe//e4e2161Ase9kjfbF5BYM/kmQYV6UWhKMNhAzhfCemtaQbfvWz0K
2w8AGqENEfEmuHvIsZP1w1NMlBY6f/TPdLs5A2x9kZ1+UVwi1yQv26Jge8tDM9gC
/OPR87r2lmODBLeRtqzna3WJhjnoW/0kEkLfCLfb2ZZSL/zD7MyEzVN9th0StTMv
hURR209yP66EheiZDv2TWNfLHxcWeObk4rFGk8o9n1AETXAkwITt5HNaigUqEBs3
J6znnn8F/A+gdQtWZjNygOUqHSg2/mozy+2QMgAB+InrhtbZzxQm/ZLWJe+XGFjp
Rok0crGHcw6GE20blwj9bjm0GhVjCLQLjxLasLZYkN+DA+PQoGMA1JGTPra3cNO9
n0ChRklF7tZgqTuFAuc5tHDwsgl1+i43y+w/UfaKDv+ACZ5RTtx7F7HERWIOD+vs
sQwfjDim4VO1mwfiJoDsmyZpEDSYGSQKbyu7IZDFt0bPzKAd5OJv4bEgStToLOcS
`protect end_protected