`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 20736 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/9huKRhRMtvnNqb3Z+UU7TahEoHV+T8U3P3ufru7l1O
3DlgtZzb9QxCbOjthp9+wDkjygH0eUfDrEl1ovhZG604iyX7QkdCLcstvE5bcWed
hilYqnz0e2rjvK3W0ej8d+uyyYqNI96xPtuSglDnO4g9uyw2XmPZhSNWPlOLCihW
3mzmr6eK0RhuLGlocSpHPNkTjBFwLa+H8VGuW83P3rlBI28PooL3HCskAsrxFrLu
WX1fDPMxV4g4+74A1Hf0mR9YKb5zanrZcvS1c03x4VnakJ0AHpXBzebCS2gSbSAA
fY2OibeNvriT7GSCWJZw+2cRr0sicoweIGo08jeaw0J2MKmCHmeqbDQrTe8N5yjU
sb73+NAFuR5U1Bx6OHyf3aeTkBxfn5KlUmWi8GSCnlNm2cd7cf/+s7rDgKKZPdSA
nw7XAg19Vg0hMx+ky2pa2MWeg4rbe5yhX1B6DgpQ9JTAht60RrdgSKkxVQMGtUNc
S+l/MVThUwY1EWkY9+x3cOYyjwug2Tg6smkpsd9HvXTmHs+WO+hJsJ3ZcJEapOe3
KKwix4e9wL2zQWx1eXc517ZBor+Y6Ue9fjsv8QlhYa1xd+AuYPfg2NzxbkXj12yn
s0K+Hnr035v6Fsay13zaktZEIlUz5E16dfPrdw5OxRoWPjeYvUlnPITke+IzkCNe
bjr68VwALCnoAvDL8nK6QkehCpFAGHXREVRP0q85Pp5497iA6uR+eDeWIjOvCn8r
vMxUv3NYble9i2zoEgVFdacNdxrucuv27tbJi4FEWFuHAB2xbCumi2gePEQ37HIQ
CUhZLo/vL/XNxmVfWcJlP+fpflHaB2uoDLXgxAnMj2iX3RknxTzAFPKHKhRFnHBS
UFWlWOcaxs2e9TWiN2szD6YOip98glIcezQv6ViGdrLol0ZTfrgVvo4UWjCEDE/6
BfY+uyWzbgC7I3nOGPde+hFQWq45A5nVeYNAuJG4p3ifIzv+sN/ni4aCPJVsIkyS
ZbRlIcJYMDG6Rs1xZBEux/WkLvRH1k9pZx3V6sY0GKW1xXXcgTHtFINzNhyCCyMD
kZLzML2BFbVlZ4DIq+LoTsAQimM5b+znZa3trhXRMPwYnSZn+u7HAQO9Jnp2CbHy
SQo8NibIj9AfG0BUhq6niOjT0ih3E46j5kB61mR8iSoMX7zT/AUshfHziC6MYBAI
7F2a3qvbz/bnW+MSIJkk4nMsGpyHHVAxyPhp2zqa7nW0LorrwLAMiS4ld1g1SfGW
H7PlotXHH+sVJe72AK9bwdLVYkiI9y3nvDlGo+xth4ik/VV41hKFVDPKh+rUDr9V
s0gbm55yHWkOjp0oaqp9UGEi5HaUfUcv7Od1rHrr60BLeS7NPRopmwg3foMsmU9t
W7vNxsZ48z76+QQ0zugGtFgfkFZ2MUQ+2nslDKwQD47zxe4tJxtjAuhnyXx/MlW4
h91ucwCf2y7S9Q8p+rDr6KEGhO9Ker9UXaHgdTZ078DRs9CMDlnPieDBiQzX6Eka
2eb0ruCqPK/JT7msXxeKT9P5QE7RkhH133SwYx+tJsCMHN9Bar640ou7dS00Qfi7
7PatzEukIGbx/WY6n6OhIyy+gwdoguG8Spv2bJoZzkLGaTiqc93Z22AS1bT3sBPm
J/EhmCoZgUa7MPOYEHmgIEcw7mA/acE47EqCS35BkjzDHHeWSGpFU1WY7ob675LS
Gg/8HFpqfludkcM5Zdd3vxQRyzJNemly/NJnlDWgUYUkg0BqJCuVGdvd4QVsu7bw
CN/CYozO5CFcE7U6Ldw61q6Zwg3r70AhUiSASftAtPX1sR5omKW12mo4O0+agBIT
d3q1dY2HI2SOckKIsTA5fMeLbYBpSWHKxL+LrYr+iqI8S8err3MW3rrgjzYkIVSE
gF3BpdOz4z1tXY3tpNP2+fHE45k7/F7FRQWk0//QmUrO4WjUvxGOiYlDg0vq2UJ8
Zq0H7Q7+nO7O4RGDxpsS4lAQogRVtrZQ/7ibJDvUTomfnPM83ckXNsIFOJN1CZ4V
jxss9GRmc4IQP8bqGTW9KGQcrq/JrHWGxk1b1UGQXfsEyUQFttioRpHvxFDfderk
0TJWwRUD5u+/JRFt4LInZVoaSmN2cxS7dNyxeqim9MEGty2S4zNDi4Wl9gTTiDmu
ZBbl39D3yjsbIgn2d1WI8U0lqvHMrYKFwpwfQYHig4B0/kwvV5deoo6oUf1CgGm0
6rxRCPR+4RIypzvWK5rtWZnBX8Ecudry3mdSBVyRBAZhSuImK51Mfj9Tjkxbzj3k
wtGL4pFQjumDUDLSKW4zv38yVhOHBe8kKg6YRY06xNf+tXJE3fLNnNk5tfKlMuia
g0qNJ4ANT/+3IoGfAW8BvMkv9zA11no4K+JJfMwiUvERwb4Y2ryDE0CDhXptKRor
SCurUZMFaoMnZqaQjsg0H3q9qUI/8JM8H3L76zVd+5tKa5p/LFQMfVIqFL7oGWIb
bUFwZLDwb6l7DSpEh4HDQLnoQ1PRftzhS+3pyRbSLFnPCrK7MLmvSusS+G2GAABy
x5LRp+0923Fx/meAxEbWYhhfPCOBOobhbDp+ZyZWnLDj6twW8/3/gT9Jazs+AFR4
tExAoiH/Uw7G+TJlVZYBgJyaKV00gbZhaeuXI6kxj/tljkI9lrEaWAFKGtHx2hlj
UIG9cNWUgnDIUoVJvKxlCE+kUyn0770a9Rk7zDnv7MgW793aWE4AG6LBB7N3Sdqr
RaQpINQAGTiPaProLtq/ZJhuX2mE5NlQu0M0rWMO5qNH1iqyuDTGToi/N6CkU73Q
60VJuayc/2WK0uGOLkmJl5sSKGA6C3n0I0AcB2rbXjKooB/DJ47DMu3cDpwqWTq3
A1eppfKg6B0VgfyG+GouXXnAZpNC4T1EpvFjyh2F/jp6qJGXJRvmbD/FHt3XoSPf
XDhPhXP2KdXvMA0e3idG5a3plBKyfH869cBGgszcoEcd0i31MBd7uZofUKGOoQCK
4u8P/QekmmDr431QmJBKNmDAXiGn5kkVi8L0Rl0WrG28E67EXtZ3iwDO35O0hZAD
Gp/4PLlk+nu8bZ9tbYITX0nyPap5FWKqME/VKuYA4FjfOZZoEuv/lz8aN8twZjiU
JRsRkDuaVCjfleu2GlOmL+2T4ey9KsiaBh6VeToyM2jdcnJp4Mc/dLLXrrQqnkZK
Hlw0MzH2p/3AnFDpPtPOu/ElOH2Rtg94HOqXM8QE/65yx0/ha68Vds2rKvsJFsO4
s4XT6470Xxd+xpStuJO2DPre+QtZPSc9+Gk83Ra6xVlYfE208d1XSh5IsKZ6Si1p
TjyU6LY65cC35hYS0bSRVA7aC24iNdQ+7sB9a9+OfDYfB/b6JMtIColbazjd16Qn
OyYhllMLV3SZD7xMGY3LY/lKb1nB959WjV9Gw/LF724aq+alhXTcWJiYN1Frs0OE
wAxrcgYF0VdbIaMLUWZVgx3W0fLa8N9dKfyuHzSPCY/HtjVbvfnVe108dp/h+AFZ
fXz9I4K5aA5ckEPQXXe6gBjMinUI/Qjl8+8wZZuiDOCHHUJqBfZJ/Wq6cs45sQJ/
hazd/s2YLRQITpd4AKx1sb+Npg9vF8J6dLk3Bjjp7HRcgqPvn8SVb0p+KO8ZRYvN
R+eVeXbftwQJ/mtUub47mBSq6Gw4gW/p0g0e+WJWY06X/x859nItF55baQeb7GPo
Mm6mYiCEGAMcKbcBhkjf+2DhIAT5VPs6BjPw4yM7FvuuE1/F83pgCy5UlpwS/ATZ
+tZkeXNRJ+DSVa5EMK5y7lLNKQjS+JQ5ToswFtMZ5uWJSGyV7IwfqJwZK3zWqdJL
yhb3M0RQJBEPfSKL92vuiWoUWRjYws1j/jxHoGWba3B3eWj638jWGJHCouhPocSD
w55OYlkKNHprR/qzl06SzjQIIouwBWfbn51CwyJ0toYodo/tSXwhXc1q9Bhk1t5R
hZOuXGfahDfoU+iDHkb3fRdIKEys8r+K5I4r54K40Dg2EdqCiecZfXSIG7dHwbLx
bmSVtdo+oBKPLu3p+kyeQcsXFPaGTA+gsC0ZghWVw80nuNfzd25rQumb+wus8HAN
8eokRkTCCzwIC0NDvguo2LnAJRHv2tUuIE5tFF/MVxV9EBEKqZONlW5MebD6eRz1
KbBA7Eyd2lGawJfVtjssKiGtpByj/fiv5s2gRu45Jioel8HUEFulFFLUzwgF4oxG
y4i4+7Q603ZldDQPCO7L/I08gb/cHxJS0AcfJzh0rfk9rH9l4ade4TdRo2hTbE7r
lr69xYAnVfCCqqXCPIPRgo3Ip0s7h7b9J41wcpEQ2oquhytWnQwD8x7I9evIGB8l
DC7j2RJvKe4klcu9wr09p/VnjGMFpGDW4drqQar31rmVOSX27opp8d6S0USZoeYT
4wzu54KSVbhUUnXrPL+HB5JTJBoTLx5bDxb6E6Z2N9L/eVWhdoV1rRVHI90zv4Se
7li76+WWbApukvq/d1OEoo5BxwSInFwxzx1fGpnx2l7SGwJiBnBKAFBxhJ29eiYm
LJG/I+0oZCSFWC3funf9Vmh50CqV98jCQsFeeJCD24JJQDpGQT+2jDBhX0skG3d9
jSSflWGzY3fEx3VA3ENT0XjCfmAArYsDY0xPdtBRnnp6OgKPi7dA33HyNXRv72FE
On+ddurK7l7TogLZaBVKOKX2nYSoENfar76iMHLrSIYFL+4H6aBFgkSxVC0d7LxQ
in31i6/moZDfPjWQoUf9hXGA6m8++CoqIXMq6BIOqlEqgbVIK85PZLw2EuziHy+W
++QCXtnriQIOMKLYfctmkkzz42sm+7f9FXw9GipgGN14pVaktZCPj4J6YMV58q4w
Jb3ZKZxCxli0IQvpWhGj7PuAoRnQujK+ur5wgnqpNqKs74HeXjGI2oviiJE+/C/B
VPC0Ual6BBfSMyuxaaWkiA4TB8ty9iiP9sefYGIY+0+eQTmyEqjmKfqDtIe+91Ib
DXy/eQsyy34W+AT462AdTswU8GdddDyd30bHDbLxXXBC9c36aWx6rCsZcXhtBcCO
J9Qk3SgAzek1BVtf+nlQwugcQvkQkPgy1e+ibpghykLWIMvfvlRJRft04ofPE4Uv
R1fhcojUaiQupu2pm7waramYIAuzOkRqGn1ALCXarXyEosbIRaPNvtBq8LebHSRE
GNiwaWDdoPPFu/JtKGRq+UIjhwdh6kHo5pcFsHYxA4u43QPpF5yTU72ZgcROQk+4
ZeGhepRFxZzRcUiR+RfA2iOMPzdPPMTlh5CMF2S6aVH/0Hk1ENRXeKL0eLezz1No
ktpo2CNHd+PEcJU6S8rGNOQ9VNvZ1vUmDGfulcMXQJt6fmPM+kaxygiNSfn+HAP7
Dnc+1oK95hrpspxUP8jDe4qe7L1cV+SID05ilD+IDh+46V75I6zUNS2Mg8KltLjG
UAZrPEfQSdXBAf0LooXUwJ36trFpyPqgmW5Vq3oPke7jV3WJn/U66eRydexHzOTr
kaPgTO+3+loAu7fMIRGWsczEAWVpWi6f0vYEkz5m1r9tDszCnE0au62aK+pa4x+M
b/VpTRg1B/41nFr1VIEoOfMzmBhqzSG0OIKDvllsvLHyxGUfDGPCOj8pk62fx/Iv
q6i3Bc3+ZPn9CiUD1NDG55/IOVmu6Yau0DNsbz+Hpf6B+WXR/fjwMQufLESLgngm
dQsZXsHEA8Tqn3Ocnuum+dQMtN59Uz3Ls7Sz+V9m1iw36FWbXwqqIPvES6hV2aMF
8CxP8R6QkS2bcv1cwVd/DS7P0bfYnuhc1whLQCWfYvvcdHikct3JGkDHuCrl/0TN
eZ70lGeAbSib7HgF0pIP/tvF+vwfV2s18XLsaWhpa1RRcJYp+tUd0xr84jyKbg2P
jp0cYaSNa0Kxe3HjyC/SdSG/WEairiEPfWpfx5ddRi/1SYwGKuv55tcOcNZXvhEe
4qvAPfdw4uEV2heoE12hoL7mXM3g9zzkhyn71Ys6T4Kv8+G/jhjq1WegM2Vd3p8d
RoXZxGHoks96TLKHbOFo/4X/i/D3qfEa1rdiCqrJYpB9E9GBd2Er17CmDVOrLlfP
dMOxm63pitjwSoduAeMfP0bNcAhAgaPwUUV3xqOJmLIg9Y1KxxuPoJj/7iRM7PNO
UDhg5x4jDtmLuOd/SW/n9dr4XevXpcLa7A2OqXh9jSpJ0Nw3AQi3GYWJOLrDM0bs
utcEEL+aNNmD0LlPw+nWPxrni4LfRKqIbgPwg6R4ISIkOB1z5XvjRrKwsZKEiS4+
zSazPw5gYZqjISgoqbwYaKJ42HyMFQ/nOABH8k0IHIWx5IP6h79B0TgJcL/odFmW
5CH+x094s7b+qOOpvrZIotsvkAZLEew09MkGhE5kaBsBkU09p9E+yCDAZfGLGPNb
dPWaXVt4ucTuSapfJO8xfBHE3deqNq4ZWfc6vIEg0bOqKRkBLaOFQEv4OJGax2zt
aMoXsW9b5HffWd4OL8Aa4QlFgqIStZJKpmEgnMpL5ARza3/TMqq2ThjKDPiIZGWe
GIG20tEsct6ex9STuBJHyK39QEQRz33e7p/cuyR+jCL4ahMQCpC4+1L7YVpPvEJQ
TSikcnMl8THfWY+8FrN57XXSaccqU0eTjscBpD+5XowlugZNU1Z+eSPWdeGFiC47
JJjrwPFN2Ffd5EWqu584NqntIgINcMxiHuGFX1pJiXJFGp4kwDsbkMHtOtH+ouLM
0EGp6ordztig/iISOz66Osle3rntWOsOcwbxNs1IhLFB4CRAXVDA43Yvh3G9zwkf
tLJ/965XryhJJc2SO1XA31DDgT73MIsL4tfzrlMuwwV3DJj/GxsbXDA/VqVcmeTr
1KI0f86BxPJm2ME0E0cv2jA3wCbxRimN22HLleV9mqkg463si/1x/7aOtY+Ot7jW
aINQOBYi0C1RQSj+bGAOkdWd4hCXxFLseZnkWB9n78hEqH6lmER1Zqxio+uodAkW
9GLeqxer72f7MqWRUZUrBIHSJIb5pl5cDiO0NLzuP7mJgB6zalm4gAS1I3zg8kmY
1D77hEMWA8fTz6ux35Mws+VU8Z2EFdQngkazOQdODWyHCd66P/Ur2ZWFHp45d6kr
Y7ACUQvJrPVQUDlmv6vsB3PEc7/MTRxhumR0ZYtJUfJRoRVkqfLmLVRbzzM+UhCK
CuB0fEvZk/LGB8H2Ym37I8HtMPZyuqm19Gv3d7Y2bXHXKIF25U7jjb5fEhOpEXE1
x6KXaGHYDJeWZGj21wA6JprkpQkGAv/IVYuaMzZUukBxUUA8wt4LIDrvFobYWxX9
n9UqA+XtFUmwxWHw7j0JRUs7bL5TZ+p4v4qtZ3esMjTRXVYO3oZhg1NGVSjSL/v5
USaT0hiDXRiYpPOUJb7JjS9s5GBJ2Yt+KuvRoKOEkKFQb10OR87CYqh6QOTQ3QSa
170k44gVJ7jYz1dp3Nsmb0qWidAb9WBshoODZQQlZ6tEAzL2L8STQtICn7piJyo7
GMqwJkqkskYrG6JT+adDBsVRY8XZPuVctjzzUuhgeRxQgXaQ+/ZngpXZwFFCBHSx
r99s0Z3CGwTqvk9B5gt4enHR6q7HTeqefmr/hvjQwhWsNM7BylFiUS+GmQD9fkE5
NX6Fy1R2QqofcjqA6FRvjVgW23kEmhU7RDk3qgdWStXKHzUj2LrQvm1loyS6z+0M
rjI2q5X6Iu99DWWH7jPUcfUUYVobkcz0z626A4JFLXR44ch5Pp8K+oDUlZs1QqT+
62h2q5Q+HKPKoR6VrT+ZnExNQSUlSfuG/WXMt8GP+ix4tfXXzO0rP5ae0wUemBvC
gODdm8s8HT27ZyHFvHt05Q5zocL1Wg5eiorIj7wyywKGcC1axh485icFBJBoAE4E
TOmfP++sY5gJJs/k9Q8cdhfsZ5go2xKC7/hy37cxRjhtWSp1ADvP+R/95Au8v5K0
mdcgzrsYjXotwAc/fQMINS+yuloKmMCyL1ZPnf9VdyoKuNpkTdKZI71jN6MntbP9
s0zq9BiCbUw2Or5tQcVG7Uej/D5244OAVxy2HETxoLnLtvEOYu4TjIwi3SM/dhmG
wA8ksNufu+HIbB6FIUnyri9XCh+IVilHtwsbRtJaA7/YXDfC5UxsLZDZuTzMD5uw
7RneIRYxdYwSuHUgosANp+1zZnesElyGq0xIJiEEmLhpd8htVJk+NO5nFoSD29Ij
hzDf5xxRMtNqleyg+rE7INY72vSlKF2VvRQsy6+xv0HpqgcRBYzwq3Dwy8m8H5JO
EG2mrQwj4aKZQ19UB9pxlotq0fP6A7TixB9Q/uH96NkGRm7VQZ0yLb0IL6SfcvVS
G6ndxt8KGtemO23YLQ83xmRdQL1fru+juqyDM2gZjfDqD/KEGBLcY9aQfBvYr7/O
z9882EeHXT3v8ECfgs2BTIE8NXVmke0iDLUiknfwjtvwebsEp2+1ZwVOFHYB1+C3
LXzYnS3tuDonqDjrQurpTP60MfspgMR6vtlC3lHaGCtGOiEBlyjc4rhH9IyMUXMl
QTw0rK5pagDfCxBaPUehSqkmGweA4MG3VonErx1j/Gr2yZcHRQSgjei4+uhmroq5
9UP9IjfU/aWxpOjD3EE9DopgrpHqTjk2amne+ipOt0XVryy7d0tdyf9wAIGqpFQO
Ez3ALFby2uJgRNRlo53KfnstLx7D2Ue7FidpHgPpaRaDKerFRmXuNU6P66Z00SIf
bBO9jkVEqX/XbnuiEFyL8E3XTA0v1tmr2bTKD9azzKQ0JKZkef0fSaD5jy9Vrui4
+lPHAxqFCvAAEblqYQnUQmnL3ojxq0LFPpJ+D9HAF7kPa7oK++s2QP8Np7z7Wpvt
XbcHNMnJxxagVd9+gcnT7XpNfqSR9dWh56YGi+kspgmIL3jgrFyzEp7n3pjot82I
RwjBNSrtFuavK1qLERCgUQvroKf8Ms80X6V1w7kBZguC0cyLyQwmMJd1+YEq/Yhy
EOJnWSP6CbYOFVF14lhutsKnFDPvmG1cS8POWwOMYBcKxoODxMSjt9h+PCbFatFZ
XAu93FBEB1BtAda4tKuESGnxl2kYZgUkQXtngvpajtwBKwk+VxoveiYxFvxkbJMo
v8xlMGXjpg1wr5Kgk0KcV4u0C8nhaNns925wt8NoyGBUoelXe2e/e/I/5tORuACL
yl8UnjsWt8IFNMeN4AwETa25F0fPTlR44bu04jcXz48XwomHN5uZoWBSSiGrv11k
No8ZAGyIvl924q0G8C5EG1ywBqJHVnbhvOjEZjHAuuLZKfUT7kGUjf4/qYuhtSoL
XL4ZNlW9PzR/xqDbX+E0c9iCYgrioKpe1COiipG9RAFhWTbBSWiq24kHWieFlKho
+Ry/YLIEH+2XshyKn+q2SYt43KQy0sUnU7jYvr+rZMzZ8g10G/zrLUzpZynZEcch
/o4X9BYgb98ECc56KVLSEvTjB3skXQ048txAGZHFWxckCJJqCd16FQ1QZQnkullT
xbXRpN+0PYXvDAV8hLjB2VAWysCiwpGVE5ufLNie6Y+WhFHgq6WJgD6u3zGT5h+2
Y2KdE95VU4L1LACfuJ34VYCh6s5rX4R5j7P6yYjfTbXH0Xk8hXei6AIwYPwqijtu
coOL64iPNKzHD3uLoxwFdAUEFX4hgp8caJE3PkPnrYgQy3PXyyvEvJ4tbpvzYGan
Q4OuPcf6/696yuESLUJTm0r1lJ7qzU0o2csijwXiSMakxnK051JbXJaM/lgeEGdf
MZXkDFABR/w4OV/ys+uHhItacaGSMpyu9KnFLHKDfE04nVF577nJbhvyr5qVWSE3
IPhJTuJRKt6PowlpPHiVYjD72KsVylG3n6HuK5WMHNRF6H25AsIwHTmknFiszJrY
DvtB74K5qvJPLRtXMlrpT4lFgiCkUPsI4AOy8NziVYIZgAsk6NTAoBKnsxdwV6ld
H9oeIu05moWPZ1IsjTRnawWngxcGWXXDf0b5CaFstvvt539vEzmAAbDgYrEogAwy
CKSp4R3jOn8/pbNnFOMSDlweIl6Q3ObsaLyGmn4dSNtGVk7zA/+rsVzyUYARUaLM
CrFlAIIsDt+/ezV2tNaOXe+yEsqca+wMLl2p6SqUjGulL2V0X4iaewwV7cMRor7S
hwqRHVlPEqpOyPTiyFCh/Rn4Ng7zRpQ94+x55gCX+HbzWkpfJAlI9doto8kkAV+N
qhwYFvhUDJ7Gg04rfJMuJy6XEcs8qyKe4sEDZFWLYD4FjgVrDJ8efwrdw2IEvA/c
c342w50kYjLTc6aBCgizNYCHcerBe0VLtJxBvSjDZNXJbi1w6IZo88QwD9fnPFFt
pePCHA80uppiv0lLm1vJMVJgTlMHhusHQfw5bm9z3r3/s76ZgsPJajfLxoPQGchL
z425Xv3eRjnl/e5pzUJJwgcxehCgvpA4bNTJ70IjrZ8trxEuZhc79MgQFcJ0hZ9R
vUi+NHuHZ3bhlRPQjzfRDtzAnfjBasMSrs0ZmV/YVCUxYKVY7oP/T552FQJih37U
9f544b+zvAcoWXNy2OmyefYDUc2I8ryFD9ZmDOJHcUrN4IXamfojkK481M3XICpu
NaN/FPPM325r7QDm4rsaDi3FtjGrSv2p8liEl9rP+axYLRL6SLtWdEYD5NJYH0+1
XR3sf1bB4VIdBFyubadGHz5ojbEklr5tOQ5d8PIKUfhTh6gDeB7yQwNgrh5CBUs2
ulkCtv7F5/RG0NCzE4FWdHou06uS8ulYS98PqJr7I7WHYTk6020EKLlMteUnuneb
ithClP00Gjbz7rzPs2h2kZ0J5TRXt15hf06++KRN4JzSXWAm6rg0ufK0/Wv+mL3o
OXU4cMt0TAvgxeYfwWqxdAcySNE0Zenydv4+NIle2XEtEPNHBwh+Rvp7iOD5k6xy
3L0H3DelLBA3nvuwP33fo8QMN3WxL5HM8aEJJtRiR8M7Ac94ezQtuXpq7MeIe9kK
SyurdpveodikhFzQLUHigkPGfIVMEnmh015uDm0+Xkjz7st2UFCN2LS3StLZqZv2
UaPLql4tr+bgwMiWzXfwxLw+aI1WQfjt45sbKuoz7FiuxqIcy65YQHF6IJetkRnT
17suwweyfEixAVYhv09Wyi7E2Vf7VhI/0wQplUECEsdS9ZD7HdRCJ2ewVyJMzmuk
syVKqlhB8puWLKPCJOWBvWwkBY+mnYICFyrm8cCEQIqo1/4Fnfx9qwZvF6BRu+kd
4f946REXcixpzXDZYQX93uYHdpVKpb29lEAPhczuUwkjyuEvOqI7rzf46Vw0tPaH
qJvCzSziSDw8k3W1nTN+0Q64FeEivAi4/e8wlf7OAfhkYnDrX6HsGOl42lsU8PxW
+NQWXs6G17dsHykKy8NVefHzJYT3OzLLpVjr9sdTXEVm77w2Dia10IRdWOu22MxS
XADrHSROa6ncw7akMIQ42icepDDNG24hUhx1jdxGB7sETe4RHVvmqOuh81gLR3xv
veC5TxM7qHVoBkRntIvgm05QvGu+TvQ2MpDFET3ipDcsUicN2hKRQUncQ3Xro0Zq
SzjTx5Ds+xFVD41OKXSuDDc/rTQKrLDVOaqYmkvzsgSDbyxXhsiNdkVU8bVfGxM1
eikLBVlR/SgF003susPICffGQLoQrKWz4VS/gA7sSFv8VbzwI0SFesLmpOHgaeax
QyVDMJxhjhr7a3Leg+fuFEvvnS4xhG7nC/B24XI7DXaDM+EfAoOwtpEdNP8ChkZ/
TiX0drkpix3tXJTnrlGNSnZ5D7HGYvEUcMHLUzAbtxJpYN3tLsziOwrg6k7yGEFt
8QvURxuCIk5NfEufEUdEPgg3IY76+C5bSIH9LU0ql1eyMbBnr04I4jvq/9C35zpn
fm5F8pFGSuH26psSOT/Ae6n7OW1mNZb2VB5khqix/WY7Es3eOgT+9FnASx+m4eP9
7TikQ+Z46oRxArCJeXmeCYWHbBn2BZo0D6Ngdljbs+zAcnBNpdSy/bNj5Lbej6ZD
XR4Pyic67i5pGcO9QzLfXbqEIiZHXcsLEtHcNlSeoiPlwXD+LzvTN+mpoZ16SxmT
ECSTOkWJ8IZEe9yGcgcS/JFGmcH3UZ8vaYr2tqWY1/vwBcVo1FchBcETP5hSIzv0
jrljyxo6mW8QjBAp5xCKhA1V+5k8Jc7Rk8ZR6WYKTKDiECBzwToxc5+nk2X+AQW9
HBaS+YyVhc+wbRhQ2vlr2uWeETO+aeKB4DsxouB/tjuRYCAC2yrkO2eAezPfn5kz
jQb85XANzH7nBxYSCjLKqepTylxBW/6haZ8O9I+0VbuiK4wfGrg13wh1lu6nWCjh
2B3cEwrcfdXOPKMYGLuY4VPGoGmAvYH5K7YerTuf7r6vGcATnXcb3I1oudMdZw+T
IFKME1/Fcc7CITnu2QkCx/JQcNirl19qiI976bAZ+sl8oc8QDu4KHKpBCNlLItRy
WacaW8soZYxzeSk+oqJZBcsIYEv27JoHw8sg51/+Oc6Lc2PLkUu/sObnMMd99Wef
pHR/krzttirDA9N1JFg/Kv0LGfJVIMIMllV0/YHIm4zQvkRS9Q1/TmpaWUwlWgFd
kVnk4i5Vy59GTJYjRX62KbDSi/xJ41h1dzyn9Q4+J15OZ5dgCG1MwOcEFX+sjBeI
ADXZGi/A23kD5Gn5J9HgvqyvKrvaqVcGlbk21FLHnefdXYngGJcR6Cn4cH331ti6
CgEgbG62P0IqaSFQkxpCSw/v7wmk5NwFlTO6TjFy1kFp+uw6aMbPe1KBPtZIdPmv
aK7B1hAuGctlyKxUlGW3xCUjYDEb5puwkxJap+bOATZnJPhNykuRc9T4jnkXJPo5
Y8ENvgjOeyFS3XEuSRWh6gEENvcwcycE9bFCVhPKQdVy2TfSd4TUaX0d2SA7O+lE
YXuPZqryvcZhd8fqY4K9pNgLnaU2kfOwXQn/ccnM20coxitRrssB6t2l/QcXTIO6
sizstawFNbn2g308a/1UpwUTpGIe6VTG95kfbafFF2vBq1UIF3jGMmBQpbEfmSLy
O4DpLrK3WA195/CHiVRz+MYDETvvJfaio+nbTXYmEPLAaLbtar/wyFNJ29SmYsyI
jvu4IOc1GCjHU74hKghWKA3/6OnnCn+weZwAwMfaMxY84wBD+TvNsMylMihihwMP
T+PSZqSGqkOQ6OyGgla18RjzqRhsn42yo/qNMLvAjGfd8UfY9XrTQeKVargjJadt
UhroS58K55P3QoKluUhmYngrqdrOVdoT84yOdrtmme7wYtoCvqpgl91buROdrBTv
BFMVJ2Id8aaIaCpSfVDBSvqzjkJGm2SUrJGAapYQtBQ53FA3Wp0rqY3OYl/5xLWg
/3+A/NRtXdrY3PFp4m6yzhFk9kwb4V+iaY58FeFDM8uP2M5XzbtjtD9p/Mw87zZ8
BN7BD+BGUm30Ft4buyWSST8v9uHg5Lf36TPGJs/sO3LfBr2XjmiRI4aI7sYEJvnS
lfLv7nw8h4Aaa3bVjJGhvh89uZn2GRZw9QqXTNNcMbVoFxyhLwotrFiRz9wMnmCG
cMT33zN3jgmJFJ+Ri5jf0MF5SMfplz8NqkuXkxZPzjuxrtK2z7ByvRfvfXqko8dn
w3pijz2MiN8fdMn0h2Dpif+elf9powyZqjinFP4GgcfXITma/PNBMZeS3Jdb44m8
p00fKartxlya2btJi47VyDLQgpvHz7bFJNi5rSTXX1bV0bg5W8AMmQh7jMP0mQNL
oPCFOTZ4gW7lwu9za9G7zw8B3Xl+xE/5Kmgor3qdCAZYV79ZzLuSHHDX0Ay8RfUB
QKc4wSjh1tin/Uz9miL2xXp05jAwLBUpDQ1t99iZQy6Z5UBXN4CuRXLm318OAk7w
/xkOYoZWqA8rxz49VcZRGL+LTHXRHOr00K5KHtUi0xPtwchVlFACAX9MXWw780I7
5jf4S/M/fVLf81NtQV9MGFxco4qD6vPJYvA7tekY+ZXOS5PxSZf2PGsKAv9n1Wdq
jPtVfPtBNidg/n7n9q9boKLkagq6r9UAr3gWqlMsktMdxJbgzoECsDVnBtLEGuGA
RRWQC2kP8SJ/e562UUPKcpPQLuxJuZSVgqneImjV0ZSiwtnizvosVRz3SvEP8dYq
VXxGXrYLdbiyvGx6k+jsrAiVtAJHcOzOSqgwIgbApwB3ifDuIUFbuWYIPIMCqhaH
EnzhGYZLByb1wshO6I8ICYEqC8GBqjc11xFky5R1SJcNyEAyt/Zkf1ZIgFloGHUd
ZY9ymkFab4tD6Tr9Z9vFMIITaOPc/AeIMzWuXXfDl5FQeDSYHDDpMTXJxwYlzJMt
LuRtvmBuQQr3gmIvq3M+lNJaQXgftUIlmTwWDFxtu3n9/vcW8QRrSo3YrBWGPSAV
ixjHPKvCDmf9ktYbsBfCwNElXS/K8A1kG5pqtL0s2q7DHuR9s11VClf+LlEyJPBV
xHDv/zIBAHx5CgqnbQMHYHevO/PbflNl+f1yyTcTtbT9FDdHKdM9cFEk3A2XslNk
HlfDxfiIYJSlGfF0pT4hZcbzwEhreb3gxbPl2tJGvXSZZUKkFtnKKnlZWGA/dWfY
YJrMn3TwACC1vZ62h7Q9Cs7pF5lNo3dZbgvRU1acaptX340oMek6VviNnJ+jXYBa
4UolfSVdKYH5x0DEI92+AQ/vaTLV0j7VCFhDdjQTLCZ8cmoy5jHRyp8YkHzilclE
Wp1Kv9xx4AF4N9ighdbklU3qteyo3nlaukZPvx0x/rZfp2Po1Cr7SJ6tqMHIPC7U
9o/OhffB4lyCWkEYap2yTB0TP9JfChtwOt6rLfKNdvoPQnvC02qRPjkpCUE9Kf4E
RxarPKzyRfFx++EYcsPKtpPAIZkypkJB2EQhgPD1Qwp+OOA5RiiUIf3hbiuqsSL/
PeHXTWP29BbkudaLdx4ojEL6QagCCdw4pF35hSfQio6mMMKjJtfrYUIhp0v7xe2/
MsV0zOHuL7gPdBVBS/NyHn+cK44YprZBhXByLd1fDpLb8ichEa7UUEK6s83mk3sG
OIJmhrt3bowoWiKGC0EdHxH2GOVnIr0/IbfTxguUh+b/tr1EzYegPDhozpuhXFDG
qB6M/5NgKF8wjGfAYoZ2a9DdeAOIBrCWKawbrmb+69rtkqMP0JFVTWUcz35SimA8
HQb89LlzVaG5zU5BcrXRdaqqVdqHDRFL16hymWVZ4n7LJTxSZ2I9xJDKsja6Nslz
0Uu+ED7YRzEkYT3NpRJMmlCm7oY44azWqiCsNErr9owHBZ25Oypy7NGvgmot2I8K
i4bhAvLPVj2kNfVE7k9IgXYr8l3dTOi4UdXhcoeq1ikOYg7o5VDY+olb3hNad6/L
Z28iYYXZa0o0eEqCKfJDYoYtxIwdG21idy6KKLkiLjpLRrMeNQPIQPLCkYKtq76+
SVdHMgt6d69wdua3AzF+HBbKJSPLGcjjL2VUr2IJFAqAgADtLRaKVN4l5rJnybFR
EONnsbxZLl+cp5BkILDkDOoXEoxZTA38hF2rJcNKr4GDpEPGV+KO5/UhsWFQe+0O
xAYLEFzH6oLzIF3hgbchq8+gOUV5Z3evikZ8067i6J3kvv4sxy4Ayms1qzD79MEb
69Eu8wWZa5Si+gUWtHCgHEN6bWldCMfzBOuOHDHSMN5u5IjLgz39Cg4bSwEToxoW
YcOzHwgZ4ycyJnd4ThC78nqvdYdKOPXCMknB2NEDm3MyKrfaeNPqnERdZ7ZbcT0z
sxBBl7fmI3XU55AN1pk9Q6HArO7e8JMXAlKlAxLgkvCOdhzYvEM14D0V5iPguPyu
5qexy+JFQGiqooW4+BCqhdRb6rvJrVKk7hpn2dquNPeTm7Ym74zthD6oVCAOtkN5
EhfUGEIZzLIF72ko4L4aTnCleKUFe06jO1GmmJ2Pwfi2mXIpCCM9vpNlROea/FFl
YmjZ/65nZ673GipqTSwLoqvWbEhtP+I+pT/Ya0UPGfOD0ezWoW5pj6N6iOxc4hZ4
v9rwy1bSBq4DjcxRB3gPiMBjPSHtyTX24oTOBbaNnHwEbCKHnhLXI+oF7OVwsotR
navLuDYzUegTiSKCXtMSoyH0AftYSXL5MlJCPrIVxP/Q9/ndGImByWH0Zttr2DtJ
x0ugPS2Vk43CvOV5RBClEmN9+Ct083a2aLBzWAI420un66FF0EgMpke7huQkkZ/I
zKVYbcdqgMXxiiwHUttCjJ76jP/qCh5z/EL2Wh1M+YbpzAD5lKoxB3mrNhuliZLl
wtNlCTC3XfYb1GlIgJ9fsVFbH9n/8NIUpPpv7kRoBZ0lzoZH73/NABXfizonhUHU
xXw0ElTL6ksU3feE8odg0X1zLaFp2WUt8DWnmXNu6JjmkrnlblaFfygx0Dfs0Utl
LQ9wJTVp1a0C/2qQWly3VqCopSyCI+0Aqgw4wPpN+DjMidM/rgvojQe5OefKVu6F
8Q7HCNPgwM8RUeCWFzvNUPezS6U7iJ1MPJCX0gfaQ83kDdJX3+aRT9BohP7RDxYC
ZWDWHja6847OArlgm9851ylZvyig205OM8ca0QSTBXJc7ujKgiFF6nylaSrb8iei
7985y9E+3dBoWyknE2kunwV+k22KWkxE/v97YrTrM1knWVnfVp7NG+Slfc57ID91
IUhTbLY9m3ZgCID/83eJZdXF4gO4r+/pd6Masw+Eyi+4yVh+tMJuO21PZ2odt9CJ
ZOFULiBT2bsAbmGsKwyigPHJD7WDlqpc+Hq0KOdVvvept8R/b+qN14ZE/ujgCtjr
LJ5LXw8CIl9XYGHxpgJUq/sHc6Y82NsvMGlY2n+X6T3Su8nIIWZTwRp9TmNyxLdx
XPTbmIPilSi2Q/TZuZFG8b5VsqkWSs2aU4IaCK6HH+SBnTT+3YieMS5crG62S4wf
mi2dzp0qkp0ojyUxImvKrcTjkCbdBcMhkF3iB3OV9AYH7AFocV3VzsSebtqWRpxE
qx5r3+5HL2hNYvLjsxHb5ZB6bGxukhcZbHd7OquU/eO/8yFPZeEU5gXjLt6CEly1
QxGzwYoT3aWJHOSgvABV/L1LzonQpLRReAOy2Cjvs++/6A/rLH+AEg2aEYBmyxKI
fi8aJZ2zd374rkTwyKvnKV5pKA7YExNP37ucnXO0QgXQhaOm0Vuc6MQo08nRwc7Z
hfQejTNzZ2ix1qeyf2phTlNA/1k2AknHWtkZK6KoUYGda8jr5IHX/c2yw3qMgv6a
OkqX5byE87VV/BvLPgz3sdE2PghXO3VeL5vK54ksmlO1KqQU6el9c3E3Be9823A8
c3FQDTBOT0dMHSZiUldtYwT9fmRY7W2+vHODX7cEMTa8L8KXLt1pTwOIZK04T5I8
mOs16o8ToVSlUZSzUdwTDem4Q5dHPVOA73FA8yoUg27WvgvpgOY76bBJ41G8ylnQ
w7+n2Fe9iLed/denu9LFpX+X90u05dOV0CBuzTmFTN4tC7jIkpEjyYLZWJFOK3+6
8IwtW/FB8Ca2erZgRi7ybZ6DI/wTYSTLVjDkSRM57Sd7QZFAFaKhNfn1sd7vorl4
6HfoSl6MQjhCJb3pUVygJmOYoR11UQMyOQrq6f2bQTgFYJE689F62jAssWOOCgTw
kcSSpZoOf7hEs7iavXXQpUm4f3GIGPKp0ioGjKK4jhLcKPkK/bxRAH2tg8MGCZiv
a83jx7rpVTA90J/52KYBSPas5rjjjJN8Gp0j980iJbQyFNRPNvcP63hLxBieWNNn
+eGRBnbVsqsZs4UTRVw5V3m04qTzuHfGYMJttiuBD7mUJZR4gNJ3cbwy6cHvH8JF
5o0wyVNik7RIqUoz7L7//Cdn79hk1dLXBDi/iK5gksYSH21ntleTmN9hVp+uVzJT
TcSUV9krGSbOdDeeuOYd+Itk2g798SWjbHL9K08itr54uvS6EhmlMuhhFv47/fcQ
+Q/tTH8wciwsiw3xItNxj0Qimz5vNyEC510lPSwUCC5V0jwp8yZlV3fbJQO24xqE
KFNuIXlE8YwjuHk9C/LifWX5KH+p/aM9FlYWPDM88Qcf5zayP+93gaXud5Hp9PUq
uIHEAVUHfR2UPwqimd2rDag57un5eVu/WiEp28N0beL81ZGC0Q589fAglA81Ir4E
P980GaZYCpR++zmsCyxBw9Ma/DnvtGbBg6qIkuXno/52cmhvn3FTh2B1NhGQtuJM
UN6/XQJGjW7dSUlL5KtigjvRB0rrptqgkH0vJGPjEsno0kex2dRxB4ipQaTcXbQy
4YObBXJj1FOzw15mIX45rSAbp3EAhBrt9tFDULmjvLMhTH4EQ8MS4hfupsxh8AKZ
9MUJu5agonwQUktwxi1yE1tn0eF2WiRckGjsRAljm8b8ADx67A/Ws4iUh8nyOSm7
jBeW0s2G/+TrqIgucPka5UrrmJF/ljUEaR9KxhA7aJB+ukAnBgkkiwUZp5Ke0izN
vgvLg7BlA/tzmJN9eie3/sAXx3hvQ1YKS4jN5T2Rx5tIocBjoO9KSYF6DexRR3Eu
Mhxw5dSMopKX+jQmO9GNZhhfnjJaUKxiUF6V6D3AmpyjiNkY8WVdH7YA9NsyeOYo
J43lfSeQD5+WUxFD0aZCxFeUfe7sqTlA6J/YCr9fpnZ+8zm7dngEfqCpVytC8Qp1
Ob213xFP9dRu5WdEFFv+8nh9rUqrrQ6tLig4twmNreHsgJpAxBuVZKlOAkmAb4C0
bvhyqDQel+sDhS+vO09Ix8J61gp8Bsa+o4TRF6lgcDjkR5dLMumg1BxD4U5XFS92
CuiXYjSld+rDGfynSZnZvc8KhqoQcu6g+Ye11otd/D92metIX1oa1ZqGiGDJQaSj
K+uYtCb8TlpdR9P2wyDpKkOnqdbAE7hYL3k0z7URIH601wTwDfWC38mY/22KbpLG
Ks5VbFRdDi2C1QWKFutaMrflHEORWjmDXCx0W1sEZTfs5jb3fZd0l3Q0gGiyM/7A
xDXUxPhrFX31cw/s1PjgL5FIeUuSDMnjkH6A80Q8x63X+tOqJuZgJGANt7zIsxkV
lF0i8hlnhGudJB6wFIWsvtYfEu19P7/DRswrY14FgY1nJgtDrKhFMVq2GatiiwXm
Ba6MtzjSCoYDZ7Fj1T/5GVLqnPBv7QhA+CmL7x+EuPTvHi6WWIdqdIrnqoUXoTIC
+KafkXu1HZPqEAzLzptvJDvsSQOdEJJdPHxPrNau4SznSw67BQ/Xg1VTwMZY/E1m
aYHGkp8ajAI47V3HXXXkVzRSMlh9eGeaDm1HjY8SwqdsEWwYOf8A3bUGonRukY00
xLAp/rIOb+REOfvPNa5GU3q3AYFgAeZApxdwAL1demNRnjsCQ+7GitrJV1N8YIu4
mUtm77HNQWHC9bo7EwG9Lpn8BpfZnCYFPpcSczriqDrqvKxszVriyYU0ocudTB4G
QaTTPalv7Ieod1HX0uyZ4wl+LzRMvjyPGVAVYl1rOFonl38cvhBiuWyEtHy5yozs
/LvlbPgLneyh6EvDa1WAW8FdqElkaltfoOprfizWB9/SIaJptojpqDfknVjUEwYc
gYguJro423QVDBkcFLc8NyBAhRFwMDIwaAL0nytEtXyq8lsYB7rq+W1PwpVee6FN
As4FMLo9CV0gEyZ1m4TgySVxY9SD6MsWDywW0wLqaLzveSFjzx0rd63LpTT53MPp
DuBYXMcs1BxtuAkURRUnf0zdeEwoVZLZ37cU3n8JIOt6Hx7uEzhrb06xmx+fS3az
PJZQ+oB1DmTDKBFiudm28fI0eU136b4JCMmCQrGA29Ou1SCCKVWRNTBhBO9DWZFb
9sGA/jKrS5wmOmBRc913AAtVTPKCOVusyLNwRdELs4tLHBeVeSvT9HK0fPgW7DzP
s+usrGqAWBXa0X45lmTQufqatq0XyYwWMtGZgXTZccmYe15igmvRG9r2SEJxAsHg
Imh4TScIAb/HmCn5I65fNED4jWfKgrG6bj/E0F3J1+KrdHcVLxNz/6zKJdhtKwRq
joD6OUHtaD5D1H5/goTKPgOq5eur6zR8FJ4PnI78RUKWOOOjHBfoJx95uHm+i8Wc
HENqK3iUXeCgSmRAAdBhQKIlk/0lrKK+nKTKyVeqGu6q3+HQqDUKecTF8C9/neVX
b2xw+mhv0cJEfkkVCXsxd8yHugk71mb01DhWhAR2CA3VVckikwkZZqfqVfZHa4el
TWfllm2HYzYsmOOY6AvBHOJkJVBfjJhUuMesk5pQ7Trq9LtMbkcWpbv/g1VTP4uR
XLrB8zjx1IoKp/dF96eyEPoiElN6x9HEt3DUh37ExnCHILdovG0eJC8lHXa/1OoS
f9eBACqvkX1Iwh2HCO1BNa8tm8BnzQeF1Kj9u+DgscpYZCoQwIsi7Y9Hm6EHQrYA
/N/cptQSyxmyg+eQuGpdKy2yyt2UuJ6TxKsDQ/B82LyKP6TPZi2sEB2u1dwHRmhz
C6oiTATzTxB9p4uFGpHBvYsy44IC3YTdOGHSK/F9Cds/WON1ol+DioTpCIFmcg7H
omEdPDPzpiwoYePzUssx5NnVSUsLcxOXnnaqMmyhAR2efOLDTW5baQ1uRwsK3ABG
evkxasuseLMiMe1Ja6cXlg9SdDd7BS8XRmlxJdM64pwrOT5zBudBGOZtXX2tPUor
5N9QYXvpuw+z97X2RX6IlJRPsJDbWZH97G+6BEVXG1h/7zbAfmjbRDzI1NdlsN4Y
63GlxmW+FWh8B44FMSGMeO2kZvuhSjc/AYu4BjEBk0dZ9fGJjCzvB2t6DZ6ZOzRX
vkMFr81VbhgRXGGeQk8K5U4Oz5eFug/Sy8Mc/dPVeufh6oU26DaktkuB/ZywDxmb
XEc++2QRfB1SBPc7oetV9VQ8b5UTU4ToP7dt8aicfdp0VUlr6KAZi+fQFBKV2oLD
dL3tSvQo1s7Dvano7Ofv/YUJ20Wb5LiDmDK2ieP8TpER8E5s4GWUAF/hUxeG/5m4
J84M9OvwUBwuHijRRO4m0b1F4V3V8JNd7kTXbxpPqhbJuekw7evUP/BnqG+5zNxZ
7dFQqce9zVg6y6hbwBd+HnTHShCEtAxjPNvkHSdzzzTK34mNmBOE3mA2iVKhUVpK
m8cslcDXHYESaIMaYPriy6wifT3yNphuDFdKHVKJkcRApW/VUjqz8Hovtj30dGNp
017YbHCNgsPsrediznTVl5SmaeHrdt2ao70wBzeR6No6Q4DFvOfJCAe1NpABRkKw
u3ECKYIhkNxbQg3h57zWnYpXBp8hX+/L8ibYdwJLXN8TKdP93UdtrCDN0UB9OnC2
jvQjE0l0VhShXLmU+2U2BvzeDrgfc7QjB6CHvynHnNvucOVhL/ZEAGf6GzLYa1zu
aUHBgFgZYb/D0CUKGttJmAyLDNtQT4+GejiaDrOWkOgMwdu+xYJV9Wyhxjzp8iFa
fmgQCykCrI4Joq7ihPulQ00TFENXOxdHQLnO65OKxQ90mGRcygauVAjdW2P/KSX/
DCoUPeiSSOZWMur+/9LLUVAi+I5IOJJSWlpBZJ4odwjCPtTXJJWyoJXj2LsDxbFS
axc6kR5DBk8+fuRNF//C5pk4tOzXmL4j5ACj0zMhqJrrWqr25QeWuGKHuDYEHpAk
kz+FSV+6MNNQB9Wpj27dkjAbRj6e8g/M2pSQhrHkaaSqAo2whHRHm3Si3upnbjlF
PH7klIvE1dDr72uP8wE0U4lFY5oLRoxf9uiiT75obTRpyF4oeWo3Qt+8SgSWWJu4
MfANROOAS1K9KsxcrnvGX044u0duZDX6uCpPd7AD6qEOtqEn3MPH+SGXNC2enmlq
06MkZPkFU6ip38T7H3UNJNW4GU+pIm+o3rPCTTTynmjaGq3wiYJfrW7eNCcVPzCD
pw69mWtzc8aDff5o9B1cZxkGBtNlx3284UvHRYlMBS6S4KW//uzHMSx41E5WOKcU
P6dqBEQuORteBmmeh76XmqHhGVD5sTtp13nOcmJp6wOVvw8YYmZ8ph7BC3L8ZLo0
yx15kTpOjfQDcWOzReEIhdzM5kIQzUSmortvpExv8WsMiWfboDefKM7pddCZoo9w
4zeloJ61A7Gye8qzmOKbcnItTBUUrbSJDGM6bFDAlDl3wv46OXGF1Ogv0tS+H5p/
Z2Mf/+Dqn2N3HloCDP5YS35aKqf+tRac8z/ET6dePZBFpoh+vz4YDDhYEPzUFDNq
i+Oq4ypsoYLCnm7mdyAYz6hFsgSkTLAnuo79c08f+7y+mJZrFU030TZmxek36U4D
SRf1wE2iH+xsa6w9zgjydeQS1G9ZzVJQTOSFukH/r9Ey5/WDsMMJOwXXRpdN6WP9
31VP5SOXTM/N+519LycyV4nX6Hjgqeb+y0iQ4dwTJhLIaLAuE79eR64t5HtEYW6m
cMj3dfvQOxNrdrSNd86Zu8OuWt1fouBhfR1TCW0HAlJ7N31Q5YuVeVB4G/EnjuEu
m3rhGu4KLcYrd2Ji+DZTLBnC4VrIoH40AopSFah/keRXU3PIEPk62hmhjeOAQKg4
49ET4Dtct5aqOXddZLMGUpK2Cd/V7vWg31mEaFGjat6WoQq0guR2Q9RR9hXkWUHE
EMzHHz+0dwewlYKWlf5GmCh8ol06/eE8i1dv0XvLWH3p58ANFRRG9WL60tXjpxb5
JlV7NwMPZ1jg8tiDeFaEAAsZPDBj75DyIHtFc/fgVa7cJgv2QQk5WRD2i004tSmG
Td1rZFrOyKEgLqDRQZmsQBgJE99WsKt1eNja2QvA+jFbIYiJLdOq/E7gmESrVUT2
lzqMr6jgQuA/nqrdZWI6yN+pgot1DQ4NmqC4mj7KHeJUvPoHwMRiqMbxKC8b1cUU
VDTttQapGiLhATK7LseVoEN6jZ1QXrMVVQNspwaJL54T8IZhaEnrT8/OkS+SfuG8
U5PwI5yJrILpAqBomPeXE+vfS9ZNdgUNN2Rj3fTPKLvQs2o9LR//jatJiCmOhYAR
y5x23Oby+6aEZjsGVQQzXuD/Uoh8QOrek8idMp+HJ86H3/FsnSp4nCp5CN+M1HCF
pNtrNBYqwU5yEGgA5qAI6thY3f0PgyJgtpThmMwVefYJtAIlUAuL3AUeA0+U7qMa
CFGh6Z10bgNu05l2vWUDwcpBcwqYHOvn1Ct0j7i0rIxa+/v9yNMANahxU8DqTkjx
wnJ1UkPUj9vjKGz1mcRCTlSelyeY2ND7mt+L0dDzFRAJmpWmZTshXKUnfXZS8qtp
crDdeZaQIe2DlTuv3OFEr23xC6SH07R3dwsKvCkU4qS94IurjbaIDlgb5g+aK0kw
z/Xdgkr6FiO/LcmaE/VdRTF7v5ZUuPb81BDUBTg9zqgeyQWZNXAvBHzdur5q4gFh
lcWUmp3l0ekvHWft+VBBG5fYVH4gpco6RH73upND5zJzXCv3O+Z4jvzOFET4BBLL
lsP2zc+ySVsuADIzkHH8SBpRgkpCps3fc9xwpy0vS6DzL0RN1GTa7nMSM5Eetlxh
0gSn/EmE8KxyFCtU2/clw+62xP1XvAOfOqVUI71Z17j3yzCVczIsPxuOQ+GOWP/r
Se9SyqzoZGKaBEdQE3Q80IJojvFSvmS1MXCRya1gmliV5GepLb0ETDEjun4cu3cW
vo4PuWpbPhmF0HFdSiJM41Vn5pITf1qFTImNXqX2iKLtQFGPw/xZsQblC8E0jRX4
OYQb/Ij68OQ6CSh07rztOAwR10J6xugQPFe80K4Q8FH/QC4LiKsUw74QV8upEtCo
aLH8tM2T2cLaC3PGWwGljebxCO2wsrkUo/x9l83dDOOnC192KO93tekOahE+IVlt
240FHo+8hQI0TIEVAceRY0onBU0lHIV4m/EVx/nSqQRvTTEIxOgjR9BBTj5kUVE2
KvB7lbenngvgaP2VcS5KUO/c7Rt085PbbJCsXqxiT5YHaH40oopV/3OyD9pdf+GD
Za5JH+uHIAiqmINYXmf51q1Jb3y/hNNjTBcDMakoCzxPwJUM2Ip+fBvwBvchacop
x53XA9zY82W7z3WvMjBrkFf0pZHR8VHkS1PO9tAuoKJeGSWI0HmCqU9IJgoLo5Zm
Bi4Ut8HDchGkgSHz3vcLU59v2JR0VZfZk6l02QGOr1SWOV1b31sb1ugAqLxk6kIp
CAuPOsNFYklhX8712nQsqwr5+lnpLlXqC1fxswzZUpkOZxa/YVHipEfm4+rZyDNE
Sifo7GtbsNnj0h0v+ANyCOqxcj4mhnY1uQ4WP6/J2X9NKERXRUhLzVsdZ//XBL7C
1Wo74Klm9EVk1/dyO9bYOc10nBw+QBtLkWQViVM0XuNitmZQ0Sp1EQuLhJuFc+z6
074owsKPN8d+9n95vwHB6MmW+2Fe8Q9wtwiJiMJMX2OfRHFwgvmld+MWRzATNc3K
h/w/Bzrn+7VaOrqJ4JKH/Sw5noT51aoL3OGG5pL6EoT8ShHiUtW2BWznRH+ePZk2
w9UQcQBeefUuZhMIQWxbxoNdVn1dATceW+ZhcHJL15jCAyyQnjElwQgHzWz7j80m
6wsMcxbUyocG32Mdn9jt940mNVqpB5tlsZ+YNBhz9koVM854asGZjaXsE88sM8oe
d0JJbygU+M8m7DjMZS+YLZG6w7C8kcp9WYBG+LPdEvwI5a8Yfii9RLUZfS4ZJHfq
+6vb54/sFqW5h/gP7A7OhNadrJw3HoZxgmRgMXd6BynW6dDmcwNjWLGs8VasVdIh
vM3CZQkUpeTQ5XfPtSiudwrB/9+kyJc8/+tlRXWq4m2dytHDv7x5YLyJKDUFSFJG
3ilO+cA5LFPTkQzoDc8D6FrT0HUm7dokOra2WcIFpipCYcdERZ0PtM0A3NDS8occ
hsfum5avJEoxaoImYjCRijAeFHBAISL+1mOPJ2QshCIuKo8XlbNlJrPT+Nhc6WOQ
jUnz9SjI2hOkaA+Vhi7VW+S147cd2yWqcBuPFnUs3TsoFk6wjdMwozydVRKBPeXT
KuwRvwi2EnUDZabGPnEPdCP558ZJkAQlFr5q+m/JBTnXDpv6C/n9cPhM4khOM336
oyPEpdwFNu50oWZdEDk725mXVz91FfX4H0aWOsVD0W2vz2Mxf4M2htCq/oFL19l2
303EOgGZVLaDeLKzV0Jk1n5YHxQnthg+3VlMDSigJ+17W1s8vBARkavIGn5tjxTi
20MhOgP5Q8sbV5M/dXUiks5fJb+Y7Ch2sjcbUwCrrQFYQqlbrY/RHYMeWrB1M5j/
S0zDFFe3JmiXbKLbB1GSO2kLvw02VwjcUrOFIed3DpOLjHwXKcILcQKdI4bY3Ya8
d/VzebiLhv3NyN1afpjFSc0wOxJbAOeND7xK4upKXNb+fgMHhaTm6lvVShmvzFay
ha535f+XvjKOqi0XgNwuPYchRiaAoLLsTWl+ajXYVLEimMVZ1WodzqmXGVRoG38X
4BsQ6rdRLPdmUG3dFWY7eCYzCUf34GHLJV6wKi1+UnqCMqJEe+arK6X/2PdAusaC
u0VSgHhhh7VRERLN1ghuQ1ggNttP1KuQ20kvNz/nOGSmBWxiJV2GOCoMJF8XP9nA
JxKB/9mXnjI9t8Up117jW/ombPfKcAvRJkdl1Vfych1V6IR+3llaKY55yy+daQCN
5UtQ95UPQCNsTUAsv9BBmtOr8KAtNbM11WRvclWIL2TA/7qtjP1KK3DGmdjUJS5P
k9/FKzVCRYVe7pU1gUZ6akXbzhR4iEVc1dwApMH2mbO9ofDT4XEPWC+dCXymIlqo
R3NkNleZ8VGGVWPh5B+rU/CGFfP4ItFK9gOYRn7p6xkfKdD6oUDdYb/nKUHG+KdW
C/kerccXH7SakXSVXQkipv/9EnI5LC1DdRsckU+B/9uyp3bwFN0au8wMNeiHEf64
VDWbANvC2cfTMmbjKZ5qV5dw+stfzmDJjt9loTzre/HSNlhbEof3SMbmNGuAtdVr
4cSZnlWOnMuqXN1a5TcmwMVO+hEcb4M6HQRrKzjpD+vtMk0OABvQLOz9crWdU6go
Bcb4H39Am6KADa8ILfnGeSUaf4LNmrevl8jph4b/cZfNkcsNm31c+Un5okV5SWME
jnPkyXgXkEdPvm60i3vJquRGoO/rRvX85z2/WAHEoweQNMiLpoPI4lGR5L1p3ZDk
+po/x713/opfi2a4ONmxOlCCxRoL4KKePB6WOAfDjbkGgpmvyoT3cG7gPyGnEpbx
mDY4ihlylfJUBNRrc16qwXuhoL0wouUn6gpUdcZaXBvBmXOjmeWCfWTex58wigvP
wzEN2zWnIKyUY5T4BlguPWjBXNsYWTjw4JJHJ20dguMQnOqFX+79LrWiM3hoprct
L9iPdA4us2yRgl9QNHdW33lsFzxVYfkXR/goK6m+vK/ns+4zukw9Hxkk1v4xi9tD
RJFH+y0dK4TBcQH4otCGk2DP/7UVPThett6Uvlb14UHb6ck3rH9xTp6zptTbgYA7
2MctHSrMhfzu1KFfdGgFgxn62qe6hjzVcJr2St60ZOdlnilW2wmZhV/feDa80pv9
CDzZ7HBde891Os1cAEiOkSdn6MAqeCUZqt4rdZMIfi0UfWOqFUmxiO16/DRhHJZX
aNIvPHantFyMV6ZchsS/Wm5msRZaexujrLOpPCq0GsVevPOpiza+MJdbKnkc4wPJ
6mNtH/mzIMTfmYJoNvO6mllHCLT/UopoNj5VFM7la7ddh4kO/tMzEFtj7AuooylJ
+yY8oclff59pt968qsDdt9z1WE0ZbF/uu4inBWANhRZWyBsP1DJwWTVf4wfsMMwV
+rT3Tod8O2B8DVjxU97VNpmnHUspvXDiooq6kZ5pqvNAJF0jE/oHPxPZ4HZHpg2a
CYDW7KGluzfOqrukGtds979RB+nxyPiNRw8BLvXQhVqnzDyebe3oWTGyW2ioCDVN
plccpuvBAKpTqTwkQbpps6hqiCjZQYUUCHTfb6wVloSBFS5zbHQWLj1ePfGDPHFF
LyNYr7UqK5UPR8347MLFTiGAUC1bgxUABj4C7+L0uSCIR4RB1sdojxzHYXo4Hdm9
dVWVKKQBafmAjIFML9/mMr4G8GsFDIhcdlQReUjmC9u3qayXgjnFi91Viqs0umrX
4C9YAJzrlDc/4czm9Q738oBgF9xV9ZIn9OQjNs97TLxMPgDYQWjzeL4XAkw2mNaX
L5EfHNtTmjhdLHb61p+l2rIhMalPdenHlfDx+hi5exVu+h6HVgDZCaHkjQwSNzVe
EhRC/flo2tA1k+QBQLbs2soA2/UT34fGMuc7h4MPv8xbmgdC62fjJXT8WtkGhqX2
CcPH4XKQqk3YH+9IrWmrXpDxY0ps7cMI28KKrmPp1JKRWktnwPFStNtfqFNtzHJA
2g/GUnWOllRk0tX2QHmShod9WJAmzo2v6qjYW5zepF+4MoFEKFJOc0SlhPGNiHjY
p3VBWT7Ka1Qrz1NaOt3sHNnflX6bDZq05keTEa6ZXgMqnFqKKjYUgrbCfKBBPSQ0
88MLCjWS/MOWJ31CubrJJbetCPxM5ugyWzMv/5A1B3l1XGRTWqXoROZwOMtNQ41Q
DY1d+6Qbvmf++EWsSb0hmFUWOrIUwRc3Qx8MFJTEEDq6BqRuI50nh6Bu/096uULg
Cy+JEiaJTWFz3RyeIKxDYqez/h7cxm9ZVzI/gYqJI+ZGQFnaWswcLCHnfmpaMNEl
NqEBm4wBUDPTFJxXYsdF3NISgdg8eycRcJqu1XxiTqRfthbHQgoypK+BOfjoPfww
BgeSD2QtqMMDOtnu6gAAeYhpaHVZOjEZ4qrgFd9NoW7rFfY+OLW7Ya96LtJTbafc
`protect end_protected