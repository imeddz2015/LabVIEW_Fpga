`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 16496 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/9huKRhRMtvnNqb3Z+UU7TahEoHV+T8U3P3ufru7l1O
3DlgtZzb9QxCbOjthp9+wDkjygH0eUfDrEl1ovhZG63mjCW43EJWrzaQmBQiXBFy
Oa38u3TethZEtWn0ljgaRhRSw0FvcNDFAZdP1I9nzL5DRHt1y3IvCqqTHYLiMd3z
DG+IcQOXqjaKrtMRwwDyE88H5hugKDnQvoHQ5qXKQAylXgYM9TebkpXDfDlBt11X
Go6SEdUVJmE1SUHxS9rskGWUi+LfuXLReyLOoRGwB3rJKUuijKqseqEn4jD2oBi6
KDOgZxv+BuYr3zkyX7giw8ZC2oFbu8LNPiv8CQqYGSWydJvgBFhSJB1TvcvR81O8
pH9sCcMRprwXm1cbv+Ukv5xCh6Ot4tWrECLPMSyXg5itoPnA1AwYfbiA8uKlDI+n
gN6ea3wNj77NY41rpyMHVWF+BaRPdYTyaKnqrosjsjyTy1onL8A21Jx8D/PLCCIV
M0YnSACHKEfUMOh6UF3EyZSjCjx+TRdYam1JJlkmTd1F6BvLHI7VNIadlDBEfkhT
eqFh8JwMTv4DFe5TXdkSOUoWj+sLQrglufunHpBHPwC7f1PcJdnQ0DhezWgfr7cF
6JztzKfYdoBUYcYLQ2amE1/VrZ8VLGWlfJ9Ro6w4nesh/DO8NbjEqSlai4ZX81Xv
iCjzqpD1qWqIZF+OS4xyy5CA3gZltPlk9eFJ03m78Q5SOBU2yC3v6u/fQM9S81aX
GFsM58JDkTPzw0yFH+U/LjeYi0glGeoR7wrPegp14sg0DnR4SSs8eitPzLu4TL7J
1XGVdCsDRwjupz66qiH5eML4HNRZv+8kO1pO9DaK1gIYh5QKvdVhnN+JUb5FcUg3
zuDcde8wFtSbP9ro9ZBtvYwzO3mSVLVHhsUI7jzmYYJQenMG60p4cgLEns5RJDgO
wTs809X10jQTisRe1NfGIBJAv3jy4lueH2InV8yWOIEukrYCE0sOubfs4bBpEOij
StGaX81dIJdci9gt+Ud0l0JTA6Knn6YYBG8ADJGzfWKPm0rJ/WD0V1pEB+xlYcdD
ncTqkpTsfmNxCwesdjo8a2nHuP1HX59q+2qu00P79IlYfudj7xPWRvgQd/GOAo7s
CKvUMnNrk695jnjAUr9rmADith/zkipOk5bnrnxBbBrde47iIkazeiF626Z0as8W
lrKTYp0NXicQPxN9hiDAosyP6DAeEB9HGIFB1hhfMtbTaa8quFomKZnbBiu4w0j4
qjvZELonrM9d9VNdNUI64JJnTsJun6Za4YdLaV2y23JRl6WaBkZbzQZyVHCUFjYJ
MIVtpVMOtD3GcM3E5Nrsalfrv2dM6TG1O1KPhGRtxiPjYGyleC570xyf2uTf55mh
mVFZ6dn++hqwadIJIV+e6Xo8zkNmh7bZ4IlcOBNwJCyQ2z3F27M866FSzJ8pKGNe
7v45lnSVxcbSbJI05jcbNoyjS+JgOBKveaOZ96GFg/3e8mRWQANE1f+VQ/NLRFqs
rECbFQlaMj3+K6Zc/ZKLVH4PyIfq5hzB6vMlNhiPL9Pq6ny4zaDBC4dLjB5R4uhi
9yDleA80vrKVe+OdDO8eGDsCX1Z8kkACA3sSzmrXX1l3akngXxHoBd7TwF0Ss+yl
vpc3A5wADmeZ6nvn4+ZSP6L39Z0V+F6X5zpvFjddbjFjKjavDa2xGiTm2lbWokuA
/Ug/yizieBBTLgMQuXD5gE4LhEZFnYm0dPCEcaEepeAURvspqHDa09G37UXeUX9z
9+VnZafXnQKPF2J4VEVIz6dZFS5TwfH8ufqoKK0aKGmvPboU1YAGvsWzct1edykx
74ukmqe5p1UVHHtpC6697DeQZGihrQuO5PoLjysmSbh9HovrdYh7W/aYG2mmwhMp
zdD66YaQAX/0OMWSW7cdNvTRLZja6WLo7QcamaFhYtSDyblncr/jA8NilQI+/nIG
3khHUZTfXwLLyiQtQ/hW10XI3fGg7EFjSUwRUli67VvFPXkR86PX+RubnOLKNrY8
hzNCMDOmNssBR1UmRdWxUwuGRqasKvfWS2NAOZzH03FCxo/Zm8GRIf4Vl48Oxhff
HW+R7m1kpsUDJQp5lg0s/2FrSg6zNQ7rspqc4RlpELVa6Vzn8WJRtnWADywn1y4H
rtvjiRwV6U/crfh5CbZ0kcaPnfmWYyqFkZMB733Pb7Kr9k4hfeFZCM84amRzG0su
0b6LyhhSzld3yo2qNqNW0Zq7iH3IQaYUf3LHE4hMBX5vFb5VEyvykyiMeQ0D2sTQ
ejtTToabxx4pQS6vPZEpk03NL31w4Cyum3lLhclRExD7XNV1h0kTi+UjIidDNiOl
IlYOK98sjcPV67sch5q6FAkafSDm4fUkTZrPY0R7y0cXeykzVPNAR9gNHQBqgzQ9
4AtrwAO7MZEDLsJTwcmwVg/kR1KjInSQbIvTG9ubzgIOB1/+doWDyDfvHRLqY+gv
uLsGJuwp90jWc0rzHo5/nvx+9ZrEbhrpnSLmU3Sg9Ynba1Oxb3YPRs/1xRNk197O
vF2CwQUIu50QjQzdiiDLdCCBkHGR2N1Ym7sG0dUps89A9IRLH/z6D9iRZ/Sdn2sY
Vfd3Yemy9xHmu8ivGY0Sf9D8DqiuEF3vCoHv5OP8Fyms11XtKsfuBkNOf+lNhulb
9pm8e6W22xy0XzCdFOk1C1k4x1S4vjRWYYe8J+dB9wgHofV8spPjOXkH3AZnmoe9
V3bqPBA3OMWkPAa2e+6KFLnjKtqJ44VSZQ47Cq5nqR9NSysxVhXnqSRIZUcPWZvx
+IjvLP5A9DBIEe0FjH8Wlo3wPieeslkHUzhYg7YfmYG5DJGLv5ZSYr0x/25m6WKp
qlHPlv5sspTrlVDmETHyPqIuzNtXskXdfrUc/MFvz5loR7Ikr+fK1ksD0CnT3tB8
iiJoP5WFEloL/gngBJ8UuGHf3PdkY8oQWd39/JKbF2MNFp0wjMwI7Yeb0z+kgmDX
qxY+L9WSWJKHquYAz5Ge0cmQ0ECxd+FSt9cVxEGsfPvUPmOG4/uFScrirFmCxhbN
MjMiOldxFHttpXdZodiw/tHWasPQ7W/M1qV8Y0P30S7q99dPkvsWmRd7IM/CupcP
LXDuBY8VOBxUybCgxqU6LZ1mgXB2GFs8EEuIRgcfh5FaeDepaudv/+wog/TMnj4F
B+jeyO14rdmhchsd7iJhJVYHYwLIpVFcfJfIlZ3UUSBttTldkZ4Khnm5AaljFVZk
Hc827uq6y2/NUwQQBqsRUpQdAqSckC5ULuyiN4B6ZjiEhz9+fB1lfCm/57gN8C+i
qxSP3JK6mGr6tKAM2WraClgPzsqSKFn/rx4Voth5fSCbNtMcZ1MNfdS82BChkCiG
jmX9Rmk+bsptiFnxWpEykDeqJFg3M3vO/6CJ9ag3Kl0vVrMnL2+ros8aUfkuspY5
RUe+jny971aKOMvg4OrVDJFaw+srbxTHTmBUO4+ZKbvXKf35TwaPMcwlBu3xE/Xe
SVr0kfK+UWx59L3KiPKXKTt/J0avEgwAQ52EDhtSs06c3/ef+KF6s9ntmGFLCo2k
V+oP4GH4IstTRoDLhkyNMXRfxU2eJIRLCbJYz8UNk+43xjSk3ZW3sskjaK1VpP2/
EyvvfwRan4Vi0/yGPsExAgwCLHWomy3tYN/wACjx221kltK96bgnRV7csg5nkgAp
00ZEMFg1bg4fn8XjM6mL7bi1wOiqr+99gOWmMOVocru4beVYkzmk5N27CHUt4hGr
HAL9I24SGBzjMhAQRcHgfcJwtK9aEg9sUxajoVc+lisHdybzG6I60N9yzu2w8h5I
tCWgmRAOAcKzS/42I63FfrmyUmAEio3PqSld3+A0PnUkbcbvs75/SQOU51JBSCG7
oYYrNejHEYaaqCQatg1Ms1P3+zNYMSQfapsvpxLGnP5SJJdsPeu+tqhvIy3z/QVl
HWYm942lZRn239VD8hf4gRm9F/O+Qvn8InxivkTUf41SXMykpZ29LxmPS0o452di
mYWFf/mFDOWa1aUchT7imEZtqTwxGxCLyhUu8a6GFkzuCw9QWlf89trdp1rj8nKD
FVUYV3sYmcPBVGbQgWL/cASuj2uWyegQ+8Q3iz9Uakh7FEdr6jLK6wimT8yA0Kzj
4/EQHDCmqGTJw+epSGq9JS5EOWKnH6bNT1PaT4Flizq2WKngGzC4G8kyUHUu3RfK
nDKhp/UQiwpyOEkmnzovDwjxPX1idZbr3xnqFrISNdNFmKykz0ZIopMrvlJMXwib
L2SRD4dWxzYLupuroOQoIGD+k0tGKaWbCWrEPvuTTS01NZ4dafCTFd+miCgq3PqP
56Wui86gy+YLBTtgLdrezSl7lO3rFkkrg/xyMktqKTuHji2KPy4hxD5CW7Bz7CWh
JOpb7hNOxDqm0uty8RaiZOHycdfpd1Tp31m2faSJCc82cWuNBM5oNP/2PRasStoW
a3XUCURZfRbye/KGrTGxwhUWzfTQM3IjrPbkndvKhKgRq86vk3UlSqFdwBxU4aOZ
JDRkANLQ10Na5AakWUA1rpFl8VUTZkWo3UGNujVe0NsbIcIZBXY95be9LowZRrpm
31M+hs0WnRZWen8+lzrrQ7w1QBuHwPyVPf75e1D2aCEUprCET6a5qZiVRJ05mH61
pZT77b828Sp4E+LupqklZFAWsn1eEOEhRxXpH5Bhkc7dGYt6zYCev2TfxjF6Q0Rn
xWvN1km+l/P+9I2HMlFv77UsGFu9JVqavz+XdId2otE0klhGurl4RVnleIJLA9C0
6SrfYEPYhcl75o5wYpOSyca3FUUlr+z8JxxaMLjK01+v7mBCn6zk/qmjfELM92js
PRpOhDf2HQMMzxDr5Cv3AgAuu8aVpHhq1JazmGwOWIKfc6V1ZDABNtpA1Q02r33v
UrflN+IgN4KGtkG4xohd+JYP8PqDzINenwBOLAUDYefimROOvAjYlYTyx06R1Fjo
xML4tW9zVJm0KqxjxDxA+2sqyNN1wljoq6yOgtlwgGdOB3q2DEihcLXc7r2oN1WA
rNuDgnHx2cEcHdczg4Bh2f6g5PbuDJqFsNx/jG5b//Q8skvdhjawZNraQndKXTFX
OPqrH5hLFh8Wl5QdOkibXuDtFwm7U3tPlHc2YdBr6LI/T+P+Q//c1arTiWzMHtlJ
LsaNJ46CAZcD6BEVdr9xZtXoxT+uk8zjNUW5UiEYm51OpJmKeMg3hV949MgC95Ng
78awbbRsP0GQGeGeZ24e3++ckH3rz03sfmCUK1ZCnqC30fG3VANKO6FWOH9p2UWp
8BOGHh7o4kgF5YDevJHoOmox9Z2hP3qmDEB6BSFKTNJk4/6Sssla1CU51Yjl7NRj
T3HV2G2vydTsCS3ecksaZbjba7NFKc0xsYblF0BZFh35Y+zKJFRfdGXgdq8mwH9N
8zUxHtyJ6GjkDyjVkhRV+wYe+9XOXk6AZtt6S7a+gmbav4LWLom7X3tkJOzkdyMG
uQ7hisA0uaZ9CdFTVM71oMhqyqNbZLKnNykC52nS5PJosUnes+yMtBU0wM5/UKY7
KIF77ExPC5q6FH1CS8bqMNxAjFAODvl/FR++VeQ80GI5cYbStVdDxEpnMPXVck9F
4P062f/7cAGOnoe9KoPn4TIV8EoAcp33JWZAlHrtvZCrjdXF8+Q5jSoWd9u2hFTo
F9+rceAY9b4HNP03NpTgVqTumLaU3+aa+2H2+WbbjCOQVsDxLxI35vL2YZHP9/tN
F7o+8+8XKokqFUWFMoN0SJNMdJqvt+XDVeCimTQlOyni6GXskfw48AuHb9oy8yO0
DeZc6jE347xF9C1XHyoCaUg5rQ3tr2Q5QFTn7EwZrFH33cRHZmi9qs6Dz5vZ22Hr
uQxwylBlpNW3/jmI+rT/9E1JPJe5+x6sSt/NjheTVy9Jwu5pvJql/SXogLxpXqXc
wWxEOtngxtYNpEctJdfs/+lzlla2iz+JjYKqHTl8RV6YYFwYOMyJc+3pNLMstB3r
+hnrZ4gkbfXZYhY8t10UmH6T0YcqEFVIdyRL/a239Fvl8eGQFAxOY0z3g9jGyKkM
UUFb4Z8M6LrTaJiHk02JZB2TfUqIJb52pSu9Iv4/fqEGI/jn9zLL591+g1YzSm5e
OeEmVc5OZ7Y0eRECCBdmjA1FtsB8me7MK3fnaq5MdPsu+RS3NXadWVU+jGZ/dfOk
6hgJnAXa1pllR5s2PSrkzqdlG4NsEgJsfcPCgbYYuhf3iMmID6WTZlsFUAaT9U0D
HfCZeWZ0jNBqJ7OGnHIcCmB47mI9i6chyIT7/uPbTkU+moW/upxaru/W0faRWwb4
HzYuEPX5x69UfCB9TkMUKtfbG3gFQ4d+4D2DaJIxNY+besoNuUMODtrv8hoR9M8q
mO4FzE9fVki9OpL+zrVZ4pC00Z72Q/fIskS0SWp/Bu5iwJF9mXR6/QZI2RFs6U++
EepxYr22Y5KPMgFNfi3dplyAXchR6oHZjQA1pYFQ+hW3pr33LD8j0nAdR1g9aVkN
2galO1qzbI10nGxfeNpaYH0yzh593YdGQwvepkbPRoEHXUCgcRmFVhBXcWap1MFV
0bqWSbUwvHLOH/NGJLv0c91bkLdvjHIKcTv/jfTCvAp5Hx+3shUOO67oChKhIdS/
ZVY3/+luKl2vEEZtZZ0D0x5mUUdMmgaynzSHoIuD4s+pY6G5SjB/qhz5wBA0as2f
OAz2Jmfq0AMLb0wPfOnuxwCeHzLf4hXOqkrT3Fp+5b/levJLuxBrTYRN9lnWOrTA
iMS7oorbjc0XLLjbX9aGyWqbUxJ52GzdT0JqTrPGM+v9lxFzEK5mJbNpOZk053Ud
nLATPSeg19EQbN3VP5ClTRxpri8WemJMaZ2O08iqF8EdAvKL07cc+P1mZZJ+0pV0
sCbLWDwgrWcWU28+XQ4M/+hqdcm8BAS0eZOPbLQiBuBeRsQUgM1vLH/lBi/v3Lm+
3C218QdA9VY+4XZ7FQDYoWZerhiuO4VoR6uEx38mdoi4VY96eZlQ2c3kpmZRO0Rx
cYs1V5a+b9NMCdcIqGAZP9rhK4yfFFRzT5E4wiTIvxkOUs7LzQmLgkZJxNq0+fW/
kRV99Tuc3ibiqvFRogQh406jBqpU7FG0TPHCjwLfyN5TVx/ithPFeLJtmGeIRAvm
RhSlevUTVvhVH5mh1NYPbFmKp88AaX6TmSLVUiZJU++PY68/rffX7/iGQ3Q2p6bG
rm1iWwlNVKG4xGwPARc1WWivrHofT4C0fkY6EyBBdAn1Hd9z4goG+kaRty/Ywy0q
U17TrB45lYifzyHz2vRDtym1eazUdwwWd8A+GLsKCXjSFQHFKI0hfO+T4rBt/n6x
T+Bn0ttwA0Bpadul091BBGKTDIhQ/Y9anHZXnOiW9Av0YNaa3V4b+tOQqz3D1HSJ
ygoe35cwUc2ebxlLK3jUj8b+dMl/1tfKFj5l89gYdWE1/PTjgyuXZqkDYBtlTThL
OEvvfmzM9Esc5snCjLdVd2VT/Vz2xlWem3RQEiP1s8wqtRAwjKU4YZyoNuiP5g7u
2fqiy2O49AX28W60/M5YPa3r2gnx0Q6JKMG7uYcAOnM7REe0p7MN9uSFMaY0ddOU
z+1YwLadXhH7esvClUbCZEKI5Kkt/U6NzdJ694caoqkk0Lx13lWKFASOqFKWo0nI
jVBFdYidNZxVHyEB25kp8HuSugjGz5rrfY3x3qicsFlmZYmIus9jC59MrDLdc4PJ
cYVb1pvwyIKa5v/Dw1sqC8q0RSjKevI6qBoC0JrxrWflonGbgUQ+pRFt33tA4UnR
vF1djS/uZZfCzq3tVCJ3t8g9ABxLFzzzwrE64mxDsu3uYrB0b+ctuZ7siCtd0O2w
oLRFeq7Ml3/sXagTtom5NUykcukfNduGTvs6To9/lMqw1shv3tC9gZszSGeiFh7H
s8MGL/uxiDSzc/aN1+87vSUZu0Egq/+S5cDrrActhVkh0wZNjHxGaS5VRMHzmsq+
+MwAGXpxwThb/b/TR/481SkkGgGXvvyt4HKVeEV/cGK3oibp3qxud8VxoGWdONOy
HeIqtk3JJ/foA7/ngBEmi5TY1C7eJwqD5sHbqz3+5RRHxRDeEQHC7Iw0YE+0Zw9l
tf2i7YgUovl5wPqpobXWLzowlHvykKu2s+01RbLwit7qng14yBgXbmzLycVIypCa
B9QtgYK2dJxM5wTMr3DGclB4W9ahanJESK7AthSvmpVfYkvKymqhCqIqZnely4Qe
jMPCPaV24YZinZYLNncaskqgiCsKfGMSFv7pIdBgHC5Za4Foylb2iOkGk05Ug3fB
3xu8b/pos7TPFnwQ/K5m7j5z8lFxpfgOfJN6cF5oQlYoMAoHlbPnnEry7u1Gj8X9
LJDXrno7Tj6G39cLRsRpz38T9LCMwymznRTuqTT+TMtFdTLfVaabQtY3hp2+ZPq3
2BlcQ3w8VGLPuX2UzwMb3LyZ4G6HF8Aol5AO5d4E16YqzHOOhyQ8yLngR3ujvmoz
0kPjjDTRkv89qhwsITdimuuCHhOInBv9peB5aF1b2VqgQ9J/6wO3flKe0ToXY8Ut
PzoJ2dYDZPOnBl/L7FHsbQL3gGIQ2bK+bpF0tmNB3KL3DDS6WcwlosTEKVltMDq6
JZUWETwMEX01DeFXxfwHMckvD6AZOqGwkzgRe6ogYjCOsZaKoMPlr88wHn7TpOMm
pj4CMrCgt3LTmfTH1HW4R0XJX6XLN++GMv/jZffn68JyJ5sR2xZ/i6K37lF0/nzd
e4QnKRnZ1QCXl5V8hL99gzDYjvRispRbx46omPP4qB9rb+HuDoN7JHX4+1qxqqK/
Ws3BYTcByhRR0Ap3LVM8SWkxf4/+VUq/O/1pDjN3Xpm3Yoq/bgGj9A8bisF3Mygk
lDHhSZUp8emknwVO2eQMwueTlrWus3nzxjXG9BJkyYNqqCZwcoKhDWJ6OKOGUtxs
ZrdPJZYd74qDN6yQ3ufr8Eak1jYGhIVpaydo7D1dStEpaUgpgCHCABy2kc/wN8Ts
MB5OsOxj3pRJU8S217P9qIqn9gxg8yKG4pX92yT1+OlggBlbL+8CUtDJrPqbX0FY
VSUiz7IOQ1Txdz+BMJfl/biRoFezx61kD5iS0Z+bt+YxjTgzG7/kHMhXpgIwppGj
kLP9zZVzXeVtvCREpci2/7YmfHY44BEESNqDzXMHD4q25AMbxIxBX97rI3qkdfJ4
12kvGF5T4JrCHvFG3xHtAyPkR8xyF/oCqweigxRuA+4G4Jv3TGS4KZJql+tCkYHl
DoQhZvP4Xk94Ty4uWCPY4kkfwQiuwcEYUj0JNZs2tVouPd4nTKsTPLX7t8e8TXop
rTirelg+F1dIymbK3nrhplpZxJh0rB4eiB5IIalkNeyxB86oIvFwqxDADmCqmrRA
jIafTPXIv3LVgzrW4Ceo4x7/qlsHK9Ocp4t++M8wEzhytFa/c3i+DP0yu9pjSApr
x6hbSu1FRO+eswmIqtDRmqD9UocdpmnCfmfcnP1gk9D+KIOyXROUGWdSpnJnO2Dk
hIL/KagHOpcvPetfB8Av//eP7apbE8NWByVuZ/7NNF7g+9rYhm3dFi4mv5CbGi8N
aOWr2fBkbjNyiXB/4sCz5CQGTVmYE6EeAu4rU86hBY5iFnnTFwZucc7414w1+b21
XysBgFlyQaiuhg+/GnTmwPdYmg2VIUkFFodpsynjsjJV7EtAKRFDmrpsCq1A0rNn
2yhy9UPWfs/SQF76czIvoh++pxw3Te944PpgNh2t2QYZu7SCKK5EUYS5jXfSbkWu
yA/Wl2S8HLWYiisjZUYBwhmiGvtyZVPFhpaaQ9iiMcY6AUAmRMigSJSWbh0uVDWp
DHM+FEiDIar6/WGu32eSou9xriKRvhEJwu7EHBFmV9mGoGlyoH9t7oBNUyBdMUST
lJJV6uWUu8QFgMGG8OHC4zOB9wNeSxg/GmBenz3b1SajPWPcIiOv5bJyudYd2WEI
lyFueFtmXR5BxsgJBiR8Z3UwmIGuwT27U/BREU9GxuywpP/0g5nHkmgEK98JgYN/
cg0Lf/d56PQFj6JLPXDqEUxBtzyFRoBFU/6DKwfROLDF98BctTxi6Tf5xgDxRMzF
1LDegXY+c0G5pCBAfWGxAja7Pz/yUVoCvxOiM84pJ5EUs/EMbJy8j5yWP1HhT0UI
rwYMSP+1EgDdYufQt2UOUQHfY+Il6DcYVXvRjFskSOEN/2+uTEHdIzdgtFiiuJl9
fgdPmZVXjOK/Yay9nzoMu5NgK4Ig9j+ibwjR44nJl/txIU37OJtZTSNamzCNNlSi
WkPzyaaLjuHpXEUgvZcXSmhwLAc/LlJ4I3AF+q4F0Y0bOlzSci2xPNoyvm3LIP8L
MW+lWmLTohgSvFVcdvEislz5jC9962vKs3mZi/Ek/8JfD8RnifywbABh75D/IoqJ
829wkyzLDOTNz/XEWRObPtO2IM+tWt4977B//BqmkHYYo5kPgy0P9q6JaouBaP8m
Yn9W93DdDpNbR/4N+aPe1AdkewSi0GoJPesZzd/RmoJuQ4xZrlRCMNty+SIUlkm4
h6q61LLj1JVwtyNCacMZoai07l1pYSd3BuJhTmXBL1bm2A9WpCC/cuJ0JkWiYGOU
f+UGE0VrYd2SBWSg+2JADGRXotse6Bz1T7CM97y9BOvwCOG2DniRV2pzg12hqFii
9l9rJXM26dxraLbH7M1J8R4LYT/0+SrS+IozD0h747cc4pZTC8IZkp1FYAW2HvYx
hdm+kXlDLo1CWjzOFodZOrKO2WvR8XRXqXz2pb7K2Y5znSx8rv45Hd33xpZ1GPbj
fmS9l0IzjWR+QkmDukAsuqokHqbZljEGLgJaLnV2EmQEYHqUvsJJDILHKgidKg8Q
7tMcuMIExMqTWU7BCYNMBVHXtL/JJZqPTfvSd/wQprR7nEux/381pGlMqKxjGa9H
9e7/K43IVt3j3lgsrcptYQF5Dgv16GpfpE7GkvRdQA+MSyHThrFrqXUOBsXhdB9w
GddJn07iVymKCfNWEII8F/WG6bBUH1mJXeyByVQlruz1Gqyb0xXFq4uZxbWwTtHs
YBFJH4AaIBi0z9dbLl1+gSYMdZRGtpCbfBPlq/FqH98qXTwkQ23u2I9oSxE9AAj9
c1daFabzAXbvnZNagaqf2MczRZn+zA4gZDbfH3gF1GBDkg7mdFby5PWBHLucAJIL
mMlhHD7GmKfVdGyqjtmI8gsGU8HLuAPUGSVLHqir0Luwc5uGXUwfOd02WqqcToJv
1163DLI9KUQcNyC5cHZJLvNNqVucvVky6jDKoEYZmHZJ8DJUgyisPRRFm/OlAmE3
Bodav8hVWS2015m5wWWQ5/83yt8Do6075CAMmKyts7XeyCHg/X9mHoDuDI8YeLqD
8g+xiqieMjK45XTRJBXWxJJUgAXFCb9hOcrJBNazQ3/CdIsPHID+YmdxyqFcVcsR
S0m43/gnACPIYOORKBtwK5JYnD2BT3uuNctk+ugXaCYwhjan6RQc92WBubmU5NzK
uq9TIVrmz9SNaUoh8EQfnUKPGvUujzHYaQ4bPu6XGfUiI7DYukPLx2imY9jGwY05
2Zeg25oYC6fC0jP6ys2XjAegWchoRJAFpS4ZyUnQRI3VXhkAGKpmA85emEgmtNn8
D+7X8oAXRsvnMd3L/X/RYXEeTl1KdB/dbcHYMeOlpOHZHQlraHL/5ZBE4WqouCPN
Ql0SIofxlkbGctPy5C6ic4vfATZJVMyCDPy9SNHF6IkebnFdMQ1EGceiOtCiDhP1
UIoDImlIcLbcFdZ4s4FbghrVwAq42LEEFpYy+sDPQBLJEhtVCorUTDH2QkX1nIGW
i4xkmzZeaBYvbD4Si784jQDLWeY+5Wdjz2NO9g/lXa/i0LFAeXRbJoapz4a98o1M
rQwRtJFiakFKkQYDCmsDWjME16kHN50JjOeo3xRJxopp4TC4J4uI32khFWv4J3oP
WHOMlfPEUuGNKxNNTXUhbxNv+5Fk6pk2KS/GWwlpylbOSF9axmLw7e9OSZb5+5OZ
tIjeXEnZq7dSyw13ykKLDlWdVUNc9KPPNfxWpINL233pZvO/M5AAEdZBFp74tdUX
ktlP2bR2ObgKPfbveQ8k8Jm6uqQ6jLqZGldlACKvsNsLNDkqBqSU6ejCQORjnE/X
LqwK5FUtc0FPaMS1AARrqYP/nrf2I40Um6d2dkdSNEAfg5aybPac+HVIyuHduxKK
ynuqKnChzS2lC4kION5Wj7zgmlRAZBT8RJcLkrJSgdB01CJLxRp+vXzcNSadEMF1
4Dxd7B7Z98+BAFNC1se9C3hmQweS4GF+nQiXGOq2Hk0BqBQT5VVXb6j1tlAdUGPx
ihHMlB2ke3n+QKQagXolUx//rtOkzmFGAf/e0za7OUlZwsQCx5Bi5iKkva6CBDvY
H5G9ZgQmVRZdcFKcgAi9Cjt+ZaSwXkPVp6zYvHkZbsyP88b8TlokTN4HhbUprHsa
nc/UjMS4G7KiQ9uf9plAV5kd61erHsiJHE4Rbgso8JMBN87pTEN8fkwuHQwQRoeA
9L6za1E2T6jFZxILcl+NmWdjh5d1u+pq9EYXN5K+FIiOtaVaaWwgFncRsKdGdClp
c6FdlUfcWXcdACQPSez71Ms/BsUKYRz7rQ2La52rzFzm+pixIDsh7MKHGevIOvLB
LJ5Nr/U0Npqxevhrm9BviwNsbUtY87IIk3TWOEBXzaqNyMXq3ll5BJu2uL/F46pH
TrpO/IGDdJqZcRvihiCUkF2werXPexrBJOFAHYIuqqg30/yg7n7BAblH/mfsYW3o
GV2KWlJOYNxdZ+exwDkmWHL2Q1DUFqhLM6Z1NYmuzieW5byM9Z8rI5OD5dNF4eTo
LpgtInhqIoLWSnXFoiqlyMhN9oV7PC4x0XE21eHUGwgF1rRpOSHDuzk+q5K/Jf4x
xY1XzKPxGcsT1hxK7+N2qCDi8pPl2um1qPYLQqvIdA04q+hEioHs0Rz7UiV6frPV
TWgYCg8K9MuqeoRqbpPRYVuuKSvH+dlzF0Lq007lD8XB4c1negGy9I/nFEh4nnYQ
M3pvZL0gdbDSRoH7+gpHanVRppQKB9jBZnrmteRZIhYOpWp+JQdzTZ/4EetuZJdS
ydQgj1xDBHtFqTBEftx4OldOlPPm/ONaT3x0sgs2iubGnsJyD862jPv1tVbH2pgB
Zc7Z32OoyyhKe3NOU3kPB2wk97IZ3uCcKCdxMPiTqFA+T2YEjsSDEgLfqpnx69XH
f1KxoFpB8MGbfxt4bxsuiV+npyLyhIsxBukuDb6tVSnwimFtT4zqZevfojzQ9Riu
TG/c3rlrwHrUoQFCJLBh1sbCQJBG2hzH4nOoTqHRGbMKVCENLBih5YAn7k9cwav+
zltgZxn7bWaSOaZ63l3uYFKb9GEeWyWN9wMu4FkvJKj9g4mZ/tnFniIzVZZhyL37
4VF5k8StMB46wkzhu4bQTms1OJgUFZGHRkh4dYI7KO/JKaF6xVfFwIReFoDhuBWi
QGbPXYD+Hj7Isug0bxgtA1OaD0wFaTw+Tl9As4OFkcDvuLFshFVfgSu8mAaWVdMB
4uWrqo2ijfp1oolMajkV0LSYDOfzcdKCtDNGdkPL8FcAd/1bCgjh8x2sZ/f8Cxi/
oi+xPSXW8686UA8Z3EVIcQDe3fglZLSGi67Pv/91QhM+td/EFObvtvw/7J4QlFNR
NQbw51Pc/mCdW4n37YglKv2exXhD5pct6lo3NJkbFhd/EyeWlAPNPOgioj/BhYlK
TcBAqkc4nzCKyFqha2Ca2eamOLd6U22+ARqD8XucJklsGNruiisAUuuORP02RDel
hj0zot57O+mtcR7HrVJwSB0h+7JNv3dsolrARtlhMEOJowqof9RMBNnvrXtYndxM
L1WglaqGFESa0iFfppUJwQGqoL/qDfgkUJn4TWy0x8WqbLxgqCheQlV1MfReoFp1
rSH8Ins9kIhOVLNpmvFVS+vCJhU4nee427ze6BPH+TAJHdl5tTkDLUEuE3dVJq5o
CGRl7v7rYM4t0FpUjn4K6mZgW2DfYL7HRe+9EEtp0+g+h4acxuwMT0qLMPUfp9jB
cKgJ0ytFcFvb4enkzWC/OMXOTOYNifv8tqoAlpunASAsIVgxlZ+8c31KqJ8wFeBU
ZevA2xxNb5HTlG4F7uwGeV/NqOTOKJ5uQiGT2Y6t9KYcZ7rr1pFni2cUiRnw3Rcs
Wno0VgNRIWANbFl+TMTJytTQ4ofkK0TBuCe2adUW57Oo+TcMgcO4aW0eHHMkQZfc
c8/5+PJwdnaUG+4jCmoa1MY1uM0LsMVF/c2fs+AUYL9tvxnUnIgIrSQBIJmsPfM3
xKj+XpmTfI0yOeYm0z9BEvjR+ZDYar3Jq6ISVUSHy8z8M0TlDiRkNtHH2iAT3w8b
hXaKgvBmxVTaBPwuJRTPYY4d2q5HNlSvRYGJ/HdTRKwMo1ABAGkqo7eI7Nil4wxh
qkJLVnrJAK/Rh+Bm6bxwd0Lfc8tEvYcR03EVxC6LfdKEm6WXiditSX4mWV5A7zv8
xgWU+2ubFZ6AgINObBaUr3w+Osn6bnsiQMPst11gaBCw+pa4TXOZBV0K56l85EAl
jZD+BoxLTkqkQGYPJrye7MzOtHDHK2ZchDsR6eiHRPNu45NHCwYUpHtgj8ZIBOui
hUEih3QD6kVxCSOAU82kEKztz8RvtpPNnSjv01qlR1BYg0oCsv0/DJVywCrXpFh2
2KYVYYdMAOzJTiNiTwu2kgiPFwlaw/TomFxbOWCxXUJaYfzH7Vk2dHs7Jb1m/QVw
IZ9DA5KXqFXvtPCEjLnWfNaJwrDNiPMgWjrKJI+YQ08TTurztGGjL3DV5lf4DPCR
+uXjqMguf1p0MHt1ZHBkvuh/oz90+DJi2seJViTgrWj05KafRBOfT/GqHp0yjCsj
cEDB4W1uz8STy17o6OkK20IqcZFgKBxxENNdVHccN5jgFC87OdZU1xkhrxSHN6fH
SNNNN9VMaHGi7SMZF/zm9AaB5w503gVNo12UWGDJJM34OxyXEEvmVVWn47ZZl20H
PcLUCuxEWZLI3Rey9uWTSTbMzryydxcMY6hV5BKSv+a8BuPS579HANHAqB0/ayCI
OHxfzOKkfNJhbgdBLD8AGsOZphnCcRTPtGvBuzl8iArTzCcKvyzQdCdVOSACPDX1
XSeq4SknU9ahzIhQP9/Qu/Zf6nvbkRYYL0X/mBntnaICts2qUZo/cVP21EUQ+vf/
jaXZzOjWhSjMkPatfS9nHD58ph1h42YIeOjTaUBt2dIUCr/V61WCnk7Q65KFC9ny
bGhuPSa4WgCx5AI8VQg8LPfZPCj215M0e4dCkreNB3XB+xwHlvnRXfHeLmaGy52x
hlaL+sEjHBUsMGtNqZLH7iy67EiDbvrUvv/CLzR/b5J33TOyOiH2HdkAcJP7DNMu
hl3/2dYvFWJ9tqyHjnA71RAt0iiMcadgJ3llOykc6yUP6y8Ymgpnh5GnnT4lpHbr
mI73R6ts5lOdbrjpW9axoQLbEWN3Po7jnih0MsPiQoPNqs6dmKEu9KnEM071ZVro
1Ta4SRzaF91cK35RhcD6+CM5G0O3+x90Mx0ZOC1gAhevJeaAN5X84y7VcYPqqZ5W
sWhVCZm+gqu0w2vLFJjyzF8RL/arf9NJaQdHhtz85QlUv3eSurGl04vcNqaUPeaa
8M3bI4l77QoHgaNERrPqYFDEoUdkFGERZITj6dmgttC93gwpO+AJcmA1uZYaqqmC
AcQ6OtDiDA1EbxoCg4V5wefYZjxabgSdjjSGXKHdW1WAZzOD2MLVq+B6ftI9EO36
vfsBgdooqii6s5kr1E4hm3cR8y2WWTjVKy4sQP5N14TI9oAX8mnEyJWwGmEdYGhO
iliUKcqkuMMnu6a51sBRxgPZo3XVGn2YgE4yr0eNk4qa1U02UmNV8SvTpsW96k2g
7vsmJ78dH91QXu7iM3ak75/viYKacX07ohgnie+DR/g1jGzkQwYgtQpR3QslFP0L
oHJAuTjZ8s98qPxB9Gv4FfgCtSqNg2ZmnGqstPFtdgDWdVQ+/0gI7RJoLUefmb3K
cqR755XElYVepXXTT1q2EX9+y7nADNJYf+nROfrb/MUE+KB0XuabUS4qYcpXc7JE
1XFjfvC/jCedLPDXFtmEy4vLUTgy40VJ8e9mO2Eh+XcRqcheyuJHcv2z8RkTDQPj
bzUVMQoqbcxqRgNG0hAGIevjlYH/7IICI89tTbHh0phdAq3dYufwf1LOYVcuqO0J
kAzTP1yKhRF40iyh5gOXbY5CNObBLGbTlSNH+xQoeRo8k0LA94U6l7QOhVhTIxtT
JBFKiufHuH+f3LJujKbmN737o9d1F3s3GFugsrnD8JXGJDW4Plkd5Ifp3R7r0J7y
hg4gof4l0Z84D7UFfwyUI7oWuwALsD2pxu3ySWu9AhWAKNBXduDqxVgYGPzLwE+j
DiYfj2XuyjxlfPWs4wYESKj0oz/2ViaFk2Vvm87TSLCLC+JH6WiQcMKDZB10z3n7
NRuNB9LDogJpPJxBfibAbsbvv7HOuEoP7OZZpco2EmruV8sX7HeMAfCBvSV7yKOb
TIvEIYxqAwAR5l0APHRm50Mv5RoTlB7AcaxM4XQWO7tOOAeepZ2dxRN9pGBzXqG9
xQCbkipih9TnY/2xUWkWmjw0r6uxPjsma2nyJT0WplZsaEHaEX9L9ksGv2jZ0bhx
1z2cwjlOoovW/UfGdddIn3Iys5AwBVachzhSD7PGV1iL3UdncwyrcKRTLC901Pbi
d2k7zGhM0PkQwViM2dkrYcjVjF4S5DgysYnMRc7GbRJLFxTF/K2e9CR7GxWp1C/v
z7fm/FJqyvAgFOYfFe/tfPJ/Oc4uSH0r4s6lz2ukOCr6sgjm/lOPwdjoO3g1olSG
dzIq3nGbyeT4INsVGRJYQ8SAUxByMa1MkX5yuiFhJAn3O7i8jGHeKGxVniBGO9y/
zjYB1ql+FcknUZMJ+6pM156wol7GV44YaUXB6CS9DmAd8/PvB25rcgoW4+NEm7vC
/pW5AN94VOabFjBkyzCkGnyblYC6MRbh4q9Su5YMMS2007zYMrhwTWPz2b+5M9ZD
Vso+Yeo9G/aE5gyzAgF1ESVoRMz3MEYI3I7T81Jey7Eo/Cuk55CwIASwDO+goUwM
J/PWAlwuUOLEjPfwaPd7aW3cHa2jeAQPhVDaZuWoGF5+NGxGs3uV1IIrvMYcu7fl
Y3yu/p5zU3gzJ2NDawKg4YSgBV+gpoS5uG9Sb0PzmOSfx/iXoSctI8qK8dZiP4vT
VKkzrMfpDNdz9vqA2LPWiKauwYAviaInedFaRPcxVRlQ0KK7lBmnDVq+jMfYEIAb
4gkrHW+0qFqoJ6mbSurW5KEykyWm7mnp4VlmtG9PfEOZ9DZUiTkWy7INaUlSFiAH
xIhxAVjZj1V5vraxJpxOaWsNS/iq0CIT3dJV4egXmGHRw8Z3gv1ielF5daCH2CpP
oA4KQeC0MGXN3rZM31kYhdFxb+eKAmqyzmEHYc9BOdU5B3+L4ypUHKA2fd7Bv+Gf
8XBGsdpFCbqZuRgO/vtYOFbRCNjClZfGp4TyEfnfbVZQIzBswwVgDtT5DHjkjlPf
t/Mji+10yobZu0IFw+WusXvs1H6QXyntBFHkGu/5byVy08nv5eBUzK/PZ0mg7nB8
uGwvxfa2m3qV1vk0jrR9pRvRYIdlo7nOSJAwZgTnVAX0LOkdSfxGkD1u/vEUevWU
/zQwQupn6IGD2zjSt6g3G3Z4VZXLOoTHwH/1RdGvTxNQhz9A2lNuBbDXc95+5qAP
MIP7hFkvIlta3/SpYXYuYh+aWO/pw29xntoom18cX16Adq8GLBL8Vy6IjbcMnJQm
f7rdK9KIkSpirbiy1z/2+L9VYjjSLIJt/BqdS8rbjGOlljPLf20zd8ZC/RoTKKXU
s3SU+dJ3knl8q1kqm2VAjM4O0qaGTMkgT1lV0b0EHNpbvfGL9hNpuWBNZW3cf2zX
R0dTK5y/HWj4Pitrx2wVWprTRAi2ebVi4JP/lKcFebfI0VWpQM39rwOFnIpa+Plk
j2RU66njAhl9u3tl1CGhN05UxaReRILGb/uMKqynUUtI0btCDz7kEk+vhH8djr/K
rXoh+CjVa9Pf/xRl8fF5irKkUgdEbRQrV2PR+7dhEtW75MtUyhu7BvwFQnZCNES0
NwAzNFPyNKok50tUFPQGG2LTwsog+Gj2RUMzVKBmulPvrkqKrKTGwnM8qw0eaA+p
BLAk0FOm9XsnGrz5nrCK++4iRhB4st1iN9P3auY1Reggrgm1aEbjE1yBzPzo9gbj
k4+BmbOUiaKzUVRFbOk21L9te+tPaZeZX+m4erSCTM+i5pXUkOkOx6Vdgxlu2M3C
Ng4yQpTBln+YuJTtSd4bh0jTiZ+4eJUcSScHKPjxcodQTJyiMBhWJyNwv9A3MtUQ
aICOMoC7stMxMjFUNRbusTlSeuS7x4hnoor2HAayZC9+/VGiXS631sgXLHP5GJks
w25ao0HapKybe9dBKJXlqnRkFw07HKh30XP5/9Z8rmfi0Q4zu42ZR6DJBTohIuUl
iDNdJU11czTbP/lApM+x9kLtlRf+qTygN3SXtj9DSJwWpD5X2R3Ggnai8DSknBIE
/XJaQ5E7uxTNeo/HOTHNdmjKKfEjfVboNgzN9qLfpbqi7LZxPPqjvJiw2OmfrcDb
b0rHKqFAza5BIgzjI1CaphyuZUo6asGRUFrBQSPmeuM4hMBqQgwCQbsIs9KsIdlj
Tg9/7nUwzSqx/cErRsxOk0lQhesqiDayQVe8tdxb11eWBWfbZcx0IQr1xShF4zxB
xj+V152dtlEezg8susEsGN/e+EIrvPHBr0H5Dfp8+cQNtTKxTA2apkDq5uPWzRSN
pJ5Ji8ZE/n4J89vpAjQgDqoPUMByuZft7CVe2OmiAoxh135zCvWRQh7DQspbymV9
iWkdlSxkh3T9BoV/+orTGypRz0B9aZbc3IVNQLRCMo4YXD3E0EnS3doEo8bWW2B9
VCO0huzxqYDswuJ/HzWEug47OWf6GVS8IbS7C+OzAHIvK0UF/kOcPRw8zEbF91bm
sQx5H1eitdnCsaWyToNKAm37BnD6FgEehXDMdmq+WuQ+lY3bFBPjNQCDplmYMFhf
RU4UYVZilcnV1GU3lu5yr8w7ir8G9/ViQgTUfnF1rRf2UuMn2YrwMQxNvJIQUmpR
k5pvMsGZChIOWdZ5bL4zsnGLMGKU2kc1LRR7F4ABo5zOd2Xr9AwevAysOJxz/MQB
/g8AXHcA8CNNZNGXqErL5yCHFiEojC61RZvbm20R5Ql3p+UNsBhbKZEersrU4v09
RiY7ID7VefR2WG+XPi0MVH6c9kox0+Du9HCaeRptWyyRcSh59Hh0D7mCUdqjLW0b
GQ4G58vXASXbckeWmqvhBhqcJPDYm8qjytzj6ZSUj5hdJrD3dhS2Ill+33Xl8Cu4
ro9pe0AOoh6pE5/L0NVuPGnbRU1SEw0I+kn0Hx9GmKWDIgtX3dMBR7ILih/RQ2AX
HJNn0nz0Q+gUgqKg45FWWRf/nY+1tIfUktX7tXsLzZ9xyAIyoOEVFAOR2i4Oygu1
8rEzatBs2mCqp2O136WTYNyIfANN5dcyIicWUaSrJThtvOwFc6rIrrOdVAHh4t+B
RDMlj4ngoPVoO7hI4vT+sADJ8EIwflVFNSr/j1j4LXPS574sgb1dsS34YeaJTcxc
/JgGiA+i4w7AQOUM8uHzZHF7k5ocEDb8LmcbsusdtY7nsXM9wz9ytX5hlnflatTv
3OSZMpDAvE2FIPaHNuZHlkrzq0ZLAmzjWkJ+WBHNgPTJviTcFv6dlLJ6pculOwUY
EpNHOcwkBOamJUlylNtJ4Y3XSXFuB3Uh7MLWm5ZlW5egx2avt1hlpNQTm3/PqNxi
sR2m3jxjZR4EYthw/h9uC8vN4VBAOb8cjpKMepncQWJadfxMFdL1Pv1ouxhurgVF
h3xB0w/kfvnf8rosoEhSVTNUUugXYZqKHBvYNr7Merx6IJtkuvvT5cja/7+izFVD
gUMGKGpmohafsOEC786FCMFJuiC9eXDJ3Ba8pNe9lG+qtv1BnIQgzn3ptFPIQhzZ
gRq2HzUoUTHpSOKlg3/XqtMDfxYlHn/KJ7KJ+NJ6tKromn+6E3mlaqsRTHpefKeV
cGvrWOYOK0wbZ2+NdMohcueQL6HWyCLDhrOOudgPAIFaDzxgbVi2R7+gTK3WT6VA
J4qOnt8zvndQ0he6P5SNBgN9l/oExEBQSKGe3C6lfmagZ0iYQKV3H2gZZkmlbTKV
DXTKbFBucXNc/NIuk3qT+xGkDH2p9QaJArbpoxT4ZDImznAEIQ/9M4bRyiu9FxHh
F6+aWZSDCI6sVoScxGHphLYrW0mlmmgb+uC9X6A1up3rtdhljBdQcXMygwY6QwqE
jVjRpS2WjVh2EhfyekytzcnLMygRPZfUUTt6RYK5jFL4n9zdPCzbxky6HcP96y7r
K+ZD3V0p32kqL2tEv7Mn9eb9BSOUFloLXXQd0V3NYjwrk5tNHmtSj/wvCAfpUV+p
Eog7SIpXY9rKg6jQOBH2B/uH6Wfx8qCSiJg+1bcKokF2M5ruNowNFIc7l4AYz/+h
baYg69U8K9o5PUFJNWjrJFRjes+Z+jJQv8248nl/KzvHn4R93NzGEGGGEDoXRMjt
ONnwA2JaHBOa73WtA9ShnVCort88LNLxXvogRgmUNMIv3pcn+OEJD1vO++rIs2O3
nrAog0bL2gJGxQ/C4eXitN5YxJb2D3LLRFhe331Fv3Yyhk0lTbbKzlvlSYpwTtn4
ij9tbu+oMg2qSftX47By54N66lXVfetaRZMU0JVX5CqX+LsD+K003oulLsZqWiEg
Ar2KHSrHFTylVf2ddLjXltQJbGdf4B+ot+45fEfguzpvgeH3sfyqznuPd6DUDc8f
i8ou2+REdaj5WhPCH/d6VQlA0wk/oJ58iNEN5isaK1GokMcUL5qKCjZwbXx7dRQk
rM/xJ/5Ia+6N1eIpen2o3uvi7wzB+Q/v+CdNlIdabFUNWU6T39EYKV3tSkTONXSe
2RbwX+uhLu6kwvFm1wEmv3lnm6zIBFyI6XFb07Ygd7R+YVh8mtQ9DVX7NCvttlqL
/MNQ5lAewqO1e115utDp5bNeKLj+eJPNwAmqKMWiykmZdBYvlYZBRvM8rJxLQBuj
OtovaVx50W5kjHIsK1z/E2koBmKUzqCK+rfGovqHm4G1vw1pS5di/DZdDIUbbknY
os8QLyYInQs6UssuhGXIcZvwBZlZpvs89reMSpnnas391ClJxbNXck9n4jkhsNUM
+H6dLfCz5yq4WOZffNhqRzKHnKt+HOCaHF3lz0zHQenkYln0+GjzGfMsJ+bnQyCY
oQSr3hI6EUgPZQ+xORAK3WUtyX09T0RAJ43lTzGt8ldWn/PecdWNr9tr/EvOerfd
bP8w1RPzLzvFQr4gYis3pHj5U02iZ61whspOmyO+itnTs2qvaQMdVdRIBEg7MtSF
bSzPuH50+MRTpRVAoXtOMEKids5S094XxfOV97JUhahD+TjVuDnpeK+cLrftX0KE
ef4nknuSdjMWeN3bhN3rjPW4iVOFF3fEqmLY156Cwqt9hHK1feMNvosCgmfRHRBm
M6mEYeyZc80v778gztwI8Ccdgjn2WiWgjNPA4KV3IdPuM/YeMddsYF90hbzYk0Vs
wlRYJuG5Q1fOHxKDZSzmZPlD/N0zCOvVT/X84qO+GudhQFqtRtQOWFtCouMnp+Fl
OtH95dztTP59cC4Je/iIw22R1xzFTu9lDTNvXn3gnonTC10iyZhhSmpEH0yptVx1
GADEFFRYZT0Di0URn1EgA2D+9QYrJXdNvRjRM8olsYnME2yRRDG4lhK9BDOL3uUh
x2zvTgNcwaLSg3BhuZLOe9KoHGlQuEhlQfuVrm5ttqYQrZqHn3ENha6/R6Ye2WL0
ZhBeCERX0iIqJ/XeMqyyLqjmfFZhtrY9kNx6esyPhIw=
`protect end_protected