`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 28592 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/9huKRhRMtvnNqb3Z+UU7TahEoHV+T8U3P3ufru7l1O
3DlgtZzb9QxCbOjthp9+wDkjygH0eUfDrEl1ovhZG63P7N8sJIK0F5bdHJ5BtJEh
jWj5SaP6UrQda1dJ4NSOn6wDWThwZfYTAY3qagobob8h1jeBAoQmywPR7dAfRV43
L8IIEmTOpbsmm8aqTtaOvwUcFTPQDHQd9QixnWsj59Y1INh9VolMpQU9Ai3FLeI0
Dhi/PXMWrzpCHZ906D9Qgorn7R37EdDK/ga15EG3HQHF780yAuriAQOQGaz5+TEE
H0AeBHnc/9jTTdVb4+UzfmEmiOvCw20ksh5mBs6qeRkWV3gRWYa8KUU6BojjDcNq
4xsRPNPtoiKWbD/ImWypTQ3uMu1QMszlfWG1qWebxgMiYyFNld2SaLm2TQSXu6zz
wuBCj+NSYmBeZZuiP1ygcwVcW4ywWpU8zCK9PB974ujVUMwU4wQTqpLegOZx/LXs
oNgG0QdbXKGyioyRWybR/iXWG69HesF5x3XaQAihVbkzigqe4QcAaRrC1a9gGN0d
y4kZv3IFCWQ5jw72xlLZUXRkKo+ZoZQ9tl+TJ2XwgtaDK8LxJo4kxyvJBQO6Vcbe
u+CG2D414pksBd+y1Ls87o10rk4GkyDTII8yZwTGkDZxFIHdeG0WKqd9kDHqM/hK
DjJ1bGRpvFfVzcD+lGCsUNWEoRSDvaXF7pKspeejIbh2PAIr1CLmKoWZdG94JlzR
L2oktJDalAG9OAbVuVIUb1Z3gFn1hZ40XCWPzfouMJ5JZfrHB/KdQU0wTBtdnB6t
v/Ob9aCVTCq/cLOeGqQqTDP7kUIpiUSfLrKdOSx/eatyEZD72VHzGjo5AM7vu57r
5jN4cnl0W8EiFsjl2wgDm+CQCyX45whj0TfxE9ol0z5cJephRU0bnp6zYme0qK0K
9UcTzxbUSGJrI8oY5tRfX+2uwBLvblC87EaXrkZhVWnVDImvGBuMr8WmyN5SbGny
6K4YoaxA4Vc2yQCdlryQjBN3zus0mabf2ZfoKtIyt8UDciiQHnMTgO9+vVU+JEH8
oKyKd5yMcO96oAGragh2ZdME87PWGJisJ78gj5hbYMyDdAJWxjwiQrtl4+x6m+UB
3c1lg2cLuo+1OGk8Kw5MkzgL5mfJAq24zXkbe9FuHY9YhkkFQkRywhJcAxWTy05S
hgKl+dfWSqgMpz86Wfx2sN1ygnjh5japQJP+Rf4peYzAQd0zdGsegWHujq63bU5w
LwdNxuEwVklVlHGZKRRC014p3VnJkqf3ScYlcIBvKWgGn6d9GAnRFugj6jnrGWsT
hdSmSVMCf96pYGR4tEHrW4RBLg1+FlHJ94rnVlg2rYElgW8EVb5xJC+axTdnvzHX
T8OtaqCwLILaTFzI66aSJAKKJfXQeSHUTFc8hNfwKtT0Rd+5AlwZ/NWLPW0mc2nY
lozBXmqHD0pCQuqQU00QBx+Nf6YGKr/l0hRmmhvuTG8K+peiVFsTiBz133acK+FG
fYxN7rj1o0M9yc+5I7bgL8//KDTiDsYw6IC5lcr6/WravUjspIJOOlRHGc28I/pI
ApdH4p0vrnFq7JbwoygO8rdl2qGQCcvfcb2ZHKmdiWXixCxjlZD9kuRxoFQoz3eN
KbiX7qXDyz+HS78HFfPdxTYZhTPFxbfe21AunnWvtORuf6rQFgBKMoiinRx7xEQq
aO4RGHnvO8P2/07SSXgRmLZzAqLpMeCWiSYQdYebvePFq6JlCn0H2AF9HPTyLvjp
boFVRaREWDw9S3l0DasN/8O1aXXUTzgZfALD2gZY0o8M+fLbRXq5nsPNZd+tK8xy
GCxlOXssAq4DvVjMdDI6ImUn7i8AKPzyGI6ATqZlbfMLF4uF1YKJBq3hgjlzYqkv
L4CxtDb8XZ591zuIA8iH5or3k8Y7BpEUHMJxYzZwQj3lcf76lhlhSQEB148H+Q5M
fmIUJM6L+yZD4h8i/4gH+TnEisIh0JLs701xd381RYFVGjXxaFcEPXgWDOqL0+Bq
2fk/WB7rgmsFdziFsVUJzcZP94tqy/DU2Ir38GbX8ndUanfq5+2DmYva3q05fa3m
0jKCzQsl7sT9/vftycglt3r1p5dEoQjQWDspGwma87zpa7wXOAdZtgexz2BmtS/6
DPBL+3J077xIgGBqt3idzb4ID6Ood9V9qs8OrpTmMDAcgSGK6gLxYAKULWq/qUQ9
n8XTq76EMW//SxovpPCaQinJU/YTigus1a/ObtqIrnHs7ZG6g7bt8OsqDmIhv4ZY
m0HBes3KpZ/aSQU6V30W5bqSeZ0/bkDvaHJhjKoAhQYNumAvUVGGSdwLkazR2MfF
GEGpgP/LhOKUT5pGdW/M3K4ZZK/42oMqYJ7OrF5rmjzvVzrJDktum246PHuqtthe
C8DRZP6LbFhpYJflH8GmfWsAaNbjqwFFA8R0EMvaCoLVnDFPAc7fwovabkHsDasv
akHpTBzqKuVVFTMqQQ7gtu+CA86rSlHQ+vePf8Zxgkc0WBUdefoHSr+B/rmk+0rV
DHgTrzGpBgheMeYHduJxnbAwKyX7T3YtYk1DiBwHLBS/8sx9QV5gqUCSq0vBU9yn
w7xj/jN/2lipS0+4KsjUN9sai6JfICyt/PTjxU69TOrArVpSfUWGEsOGhSQNuwsG
BLkkXfeWcvvR1vh89VoV57R7jxr8sMAJ6iIA5X8DnCaRCwuxxTl2s3ogSaHZT9TV
fxrHzS5ExpgXhSNxRxMffVx0fF25D8wYw/e8iGhOQLZgwXP62DDKm9xMNF3D/T2G
DSn7aRB6eFbsucXtceqndZ22QrailRenHDuWajA7QwBFr4ajR3ReXm6ic5LTsBZG
IjIySe7X8jIdqpalpc1Uq0L9pbt+ju/1YNI7UJ9se0t5uDgNjBs2XQSaoO3lwhQj
1kid5m83RIHizUD/Xuk+4fvkNlMybLcPCJk8nzPgyF3IbmxNJAPpGWB5isSfqT3O
TvPD4Iajv7sxaOJ9UymDCGA5vqj24ZQCll7lRLZQ/sxNFmQRJCTladNigq71OlwM
yRuoImpGBLDKA752i5mFyx19uPYV7ptksPx8dySrhd91g/waoieayN+/1j4fH1fi
77zGCYKj7mjD3nIxYdVFKC7FnUyPXAk7BoSzmgFwQ4bXthfWnV8Bm46/Lu/lE2rm
r/WKD7taXk5n2iqedF84TGvr3g0HCeWSpa/OZsMdyJPmkYGIHa4utJ95LQnkbn1T
M46gpvbnPyW+PwIamOiYjvh/HlmDxSxvIQ3bNCcUUPfw+0dMzrf7tsOhb/IuFIlD
XU6/A18eaEFRPXjB1az6zME/dg9njJMw5eRI5VzJPjicbguFu9nx4GCeFRAGX1Kc
lSHWcg54Uy9PZJqMwDO0E8PH4ZZOvTUGt15hhnp05dC3dx9EE7Q6Of9GWjrbn9NQ
ALMv7ZpCGRiUpCB3Aq+31GEGb3aFt7J6HaviMowgIE7S7qUVTdpdWz+zU/OUtjuc
dzRI6muF77Yhv0Vl+Ynpzlc15XyYK8N84rg334Wbonzpsr+EcyTwzweiZLoeZWfs
hYQZRRta93nxEKhy5K4rHyrbq5qAIMTv/1MSuN7HXVcIsDrqUlJQPmT1N0X9infz
1d0EWx4YkPvKVy4cdcF2RWAUjCLqiiuYNrWRFeHwrCPIHQJRpiKg1E84sxd8Oiks
5Ei7uglJuRIhjah5D5GamZVtNCYxdTc+WTG7kXHpaiVactGYXjQdfafBYmxlTuC0
6+i5iac70ZH59LLvp1v4xAAnRvUwWL9XswtvsnrEVl68jreRlE/Zy65lnFIynf+z
NcRVq+Gig05ueiSAErBxQaEbxV/mJJhA6ZBXzYexehHedzyGCBajHEBmVeD7V29w
KO2ipRHsIRDRJKfY2GuOCMcW00q81IhhLJMuc3z3hOfULqTEarI20/oP49ucplRm
/AD4OC0TrH5BQv1FxIT2pOytSpSzOxf7T1du8V4nxuiM/LI1FVcVQ7P6J/ALONLG
s38FzjqMr+GY1mICl+DJ2knDNqNUjUWQ9vkKbHXbXaPD5uQQxtfmVA05Cuu1v+aV
Dt+LQK380FOpYLNW2dH5aYU2o7i9hxAXEsMdiBent/rpXscvOhL2RU1262E8ydEy
d08FVw6oxUATLLYNSWshefujoghYUJ3dxwlhTgFO/S58njt5csMZ8nj1l+Lmd2Hq
5vRf8BQp8HOqZQqkd+fl75yx0FI453//CIlgN95Lmhm2sjn1O7cZOvzh9yj7Qd7w
m9vvRBX7QfWwaMTjzkeyN7/yWORMkGA+AswC8tszGw/hknQSO+nxy9PnOV7SYVmF
Px/ZJg2kXcLCy7LfGrM+2MHWNBMEwkqMd3iELz2GfzHVnT666VzXhqK0Z6Y0hLu/
Jk9/v6GV5phf2wOTmYV1b6YvbjwYyZSn7AKzTVRSnvj29EQEnL8hXtdCWVHqp7JT
v/KRjqmvqw7pYA9dctQqdBjvhdOiuJ8CS0u99yLelvIt7w4VGYh+bzq9NcXfoWay
+APZwYuwKccn0IvN4lsvSmAQ8RNQ1qgCmcvwPjtkC0tv1eGbL/I60zVuPh8RA2aJ
GNokOpiw2a8ijDONJIE/P1sKzznth9PsSaCsXln7+k1BQTDUngkMIhe6SK9qq+D1
7kd30VjLW+YI5RIOQX6KoJHgImcIuI9ljVb+wsnwY2X9yux1Uv/svuVftvgfp8p0
nWX7+5H4YFIJxBCSiwbavatTDXrO2j4lk7VjBXLOMREHAhbuDb1qWHpFAOFVjU9x
ZZHVFlxo7FaeMceg2Aa2xe4VOH5LGLLSkERmU1XzIXOkD31fisEwDC8VgVdtwAhr
PV68RoO9AUhdCiYa5MHBCrOxUNMWJqCQQFLINagNXaU7+IiV/9CIHMl7TIwrf2o9
dh2xbyWQH5iDjZJKNSpFWVENdtLaTHCSlHOk42h/NUQVyTBAdMqyt0PC3g4K+33Q
0q3M6CVlVlpcECPN/AA4Hu3gWrjw7o/uxwnqzuTvJf4uoDTNuvokkQWMQPPa6a30
vRo+dA4rt7tMrXJr0hRZeceE7D98hm7RiBspn6YRoSbEzIBJd6+yIJgytPw0ATW2
TpiFKN5/TapU5VB0ty+rS042zq+yQjy7hc/DG5+43Qcp8n47NLNDXZxQfXtWIl3n
ar5xUHMVvlmqBMg6plJqX96l4bsWwMVbi9gAuhh601qlzsVD5Zf3uNV3bJ7irdzn
iwa11BbS8WzCL7AKVKAyFrsHh3q4cMbxErPRe/nDPmHnf5dw03qk2UqQ19KYaZhM
9oTa6eJ4HGPjMimXeWmTP63HA7yX52WHT3shS0Ktt6hzJUCumregjaRTtnLrqtxn
v2krByoFqg91daO53J1wYtPPBIpbOmWQDUf5omHKzdYAmkX/dzc7SkXBgJP56K/p
OEzDTUK4+RXJ2KR20W2zpa7O+Yo7n/aX639pxOAQEUJJd45ts6/EjJc0t6Bgeiox
wJXHrGsdhFEE/BUdPhLaBqofEccyDAorogYsHDHCD18zyxuiM4xzD8bZ2IT9CcJF
bihqoXnnID/GEdYi8uJEfeWr//bq0DeLkWWRik/fjeEv/8Rl5RLepegHz+lGP8WI
U24thHzLKCVF9qBAPQsmg6sLoKFeT/i59ReBKRw1wCZgl96Zao0CcZYmeGCHEwU8
IguhUnXxwnf4JsJ2IlY2M8CID7MXnO+e7iCrRPCU7tVxuKokclgkhxaxrQ0cKX4A
CX2IV7iSQ8qMrAkiPHOSECMs1UsZsLa7nrGxHiaSqC4buMTJqFcK/zF7OKmP3SqQ
pHPMXcR8tp1DYne9KE3tQGjzyjc1PtuZ+vqWQ3HIEmrDAZgUjh1v55D0P3uwnqp7
XrUxqWZKVfsXPEsEnHNgokx3itYlpHtwzVZ0kD5INANsycxYFi/RlFLPGUyNMGVW
Hg+YN7F/NL1gK+lwE+iRI1TQQNFfZq32/MAEdB24vA29vbUGbVhDwcgoIoqzSON3
+GLHQ4CXA3jgnp9HbcEjB5nXGXdoDQm0gFBqG/bgsh5E8Vtl3Vnye1nJdjJfxDvh
g8gciF3uGKq7/eAptGMYQ3Ld1QnUx+MM2OwiH7O6zKjDJ7vOP7kEb64ePU2TFACM
gaO8344uDgNIyqegRJmSP/VbzVz/rYh33uUhF9iLfvF8MeVBVhKbKtkxYZAupzBp
a0KsFJOsMvJvEuXPkX4w3d57+uTAEL/XkYCP/+U5MF4rdzp33SQfkVzt/8EaHnHM
4U7f+GMJf/RLp+9v9ozWuDlY09db/Emx9PyC22l7OGMQ7ovYIBpOtzU3NdBg43N3
Ci81XU4DbX5yMZUiTDCJCe/qekonYuRbnTlxlTYtC/8Hc347v/A69G/XehYr4+qI
+MxBUnfKkQiiiGvrTJ7gUyURSzApWQs9vCH1AAibOIRlRAMSI0CubkBtmbHAB/+U
ETe+A/5X3g26HYZkzWfWPxpKidRjMyL6WYvcqCi402IOVJEaEXK29N5jl6QSyrYL
amtDmZoR3LRMaunq1CAn+Hvi/pKn9GLdxBs7pPBunsYFKHIDJXHJglFOnaDpCGON
rnu8am35xUwfVphwssucAYO+fgEMtTpT9m493Br3aAFdI34XXrkmlPXRbNyJl5HC
054xnciJQsYKsuOQmNao6qeMqewMOEcR11urRbRQs0ycwWcisG8p1hnpr5jpD4lv
K28U54Sd/jjH953nGIC09Dh0LHtvXkmCXrT6kLpclaJN7f/qMz6ecZE8p0/1UpDW
pV4A7F3clKV+6OMbsiyOwfR0OFy+xlKq2xUPaDmKhYba7rUg+KBx7iAjlddVxNYI
6+n56xnTKWWqUxGwv7zt/qKJELJa/1R2NlFVC52bCfQ+nkOsBH9HxGfqjKYSj25s
niZyoI9apgYTqgI+1G2zVmtk0PK4m5+cIdI41sqf6kRwQ9fr04t0MHJpe3c3JnSr
XG0S+JcjQ31wq23GSTskyTwAnpDfLVEqs7ZK6PuZqkcG/wQzUtqCUEBcejQ8u2JG
00qictZhquFO22PqdE4cRS96qi4WMPaI50fNHmgaZtN+01Fx6zpnWpteWwwk4lGE
HicGaYNErs0BSdeyiuujrXkg4QX/uardzvAjqIdO52JxpUsIh91HDgImF3ZRlOTN
k9gSwcxo3pEVGzDgzMxWTvw50J3T9MecrM4q4+x+6bIGKw3fvbAUtsWvUB/QLWbk
QFqRYm65Rd+oFwnu7Hikyy4wW6QA0m06YyFBHM6kTlHn+8CYs+GTZRj57OVkEOpL
nAJgD44FcclxNgoHoA94vQeOkmD59BjZVHw/n4yLl32k+KRZWnAm3CtRBqEFr7vd
+JxJYdDeRlHx6hXWVtM5tGrLw1sGhoelKvXqakcq/OaYXFF7Xz3lacxdoP8Xe3A1
8i3csTqbJzm3VmDgRT79MT6onzp+dlBkGQSnrv8C9kumVyK3+rPypVjtAARgVXbO
/KHEbY352tTwu1hRpqv3hMlmC2b0OPRfu3eNAtX70l8COcFdTfn7s4tlN/FaXCWi
MVaLGGwmHXG77/TrktzGJXryh67cl9iRaxZyDO3i/HDrEpzdGja8qE2yA4w1aX5k
c49Rx0s14OKj3cfc5EOuXbpTiPw+rUoA4I99uakju5+pabKWjOJM2V0UbB7JbSSc
WizQrllXC6C48lZOs4+I8d/VXhfz5jSl8fk3PvlVUrPGK/LmjpVzpc4M2NC4aOVc
DJuVj46Jhjg2jJt2y3ibF0bwGOHZZoR2fZBBuHi3gRGYcXJDtOZO/LqCKjigehyV
ql4lST/SyV6wT68goyVTnTDBCP/yNSYpQ+xuTSiTgwqQELLUlDJLBqKdd6zX0Vmk
hvAppiJoE9DRkabC5iWV9sHcGzDI6/kNX2NzgL4s6w3Ivo0hnzdnOeaWYIzHYqzL
Yck8O4lXXXcSGd1dyh+DgpZmD8vWLAGbtfz40ffL3t0ZmtiuWTnfWgDPVLW2jFPh
n7KXnt3R+COR4cGGyzoO9KvPt4kxifmkA1mdISIdsaIKV26QfthsnhkA8smidyk5
Libns7Tb8a95FIw0LXrp8ppGYFza4n8sbOOVBswtHeG/qfEA5nNTIFr8lmKCa+zi
2k7fude+/7v7gSn3BSdgJ+zdXtY/eueeYRbAnYifYn7NR8tjDVYhOvj5nUg+9gO5
ugS9fm1yYCK68htuyFO7+pYFERoGSatsKyyDE7gEaHzhJXcoxcedgvvW6umI5UjZ
haqfYth8+KHgGR8Fe3fhAdUyVYMmtu/DVIn4Fv5WkgluSwcCuUWjF5CHCQDU7Hh2
8rP58qjwmqgOI4X6Pnt6+zWWB0btVNoJ2Xcrs1GtCw3/PY7sABWBBmreBa6oOJPr
i8LmyxvSQv0RVG5wsX+jka68Xi2oQhL4eXUThPxrH7h3z311/39JEptzJdsK/vLF
VN74oXd0o3LBiDHYmcQEqgEFrjdJUHuqYgP6vDb9NHlXhd54nvR2HNefcQtuTbXP
+KYK0LQiQYEF+EPqwYSgqpF/0mxMcCloqzhcCe3Jjl8fqMwZcAv/gt/jQ1/+xC7C
Vx+Oyhz6g1bR+C/eCm1EvJXiiHDPvLQsXfc88Ka6SKs+HiSOH6ppw6ZmES16V9MI
VNQNN8QnuDV7cDFIyVdVaABUmX3k6N6OCow4UQIuqaenKEK0Qtti+eQ3+3IzZg5B
zp1lF/rWfI1qRW/rETqHHdfr//1oaj/JfOxZ7xwrIKnQ9XSbA7qEzHyGECMmgaD7
IM6aMuw/EyJkeQL+He9L+56fukkHrxG62LLwInO15fbfq9vRrKqaFAh60VsOZNKa
CBd2LNQWKbqz5IbVelK+3hHb6I+bb5FsJun86CLIclpYE+/4O9MfLu7HkLUztZz/
3Ga5+sgjHLMlEo5p6I2EN4Q0cJhpq68cp/F0MURAdEZsrrOosW6R0ISLpxpAz3pi
dalnSHgs21RM+4G1IEOH0eyI7HT0aIXUKLVWwiYUYZaEZ/QcB1n5m2X9ftx1i1eH
hPnT5U85i7qh4ZAe79khlKvP5RQl7dagrLtb/NDMQcwdyN8YtbwLWsDvaoJ3WRJp
WACeMhAfad/vb+kXP5FC2kXkpRDBh2Hxl1IHp9LIsasiCX6xhD95mfB7HWy7HwPH
T8JKIGe6ZD26w1XZp3wRRWU9nyQpoCbTQYN6dfZsOp6rBiHra3gZ6xnXngXp5jJp
biXohIMMyJdjt24hKcz2b0HLTBYaZig7ONfBV6XPsHIXQwNs8SRPMAsYLqj9uRWh
zvrkf8Zv3V4xlKZRlKMgl9G0OygoGVAoZNTtWF6WpFSPdxB1tdCoc7BIDO3y/sYK
SsmURtBPjXwSy+MdXaUlM548b4Hflxhnp4L6VZtYd9KG42rHL8WScNOlp5lUo4Ms
tiuFqgNIhcGK6drMaojTlMzOknz8LwYZlIssT0mbtK7v3B+gAx77XeDeLyPwraQd
aXNyxIJJG2F2fWi8zYX2no11N7V4EBFYFMBav5+b+x+mNtU7QTIiE3V252hJGDF2
/5Y0DqKP6XA8R+jJt52YKA4i5ED1rfdYa9envo++HqaK0zDCiCRBms/cMULMtBlv
4RnSq2VUjNHk0kTW6ea0m6ovcscDBGETJ0FRGA8Pf3Sfj/jGE5yCvGt+4K2BgOEo
jhVHWgxHGTIdhHeK/UUP5i+sZ4QDqcXRzSVeh7mcYcA6owqHiu1lekeqdBGz7/yM
klSsH/dm4BPtDE9LjU/7VESZ+UUTGmJ7WZTAU7RBpmxBOCjQPN+Te+BxDfWgxWyy
vWaB9Mtb5rzBCNR7ZbVjI4Frzhyk+Yrr4tnpIU6/2QETBjkbvTJZjB3Htljr07Tp
NlzGT/swd1LaRF8hlkg/XixQzXkjAlkKqw1xdjlx1QtMfAhlNxo0L/n1cmOrImsq
/wAA58ZN+Ffk0hVUCpidz4wacR6ejBWcWbcZOE2o2cZJdNhlQkcHz8uI8GBcTzxK
vGdz9KnC8vYSQxpMuHFLpE/EVyitbw96R9RM4usYEGBhtO7ykrCCk0UZffNnVNIq
hNDti5KrzQaPwH03LI/x6909Tp+Sf961C/HQCqxKacuBS7miizPG/hpTmNtl5Vqu
DxDmES2jbAaAlttqBpCQb/8lgP4L2a7j2vVtJiIg6NAUFXmC3qMNmSyS3ZP6DAPl
fS4HBi0umnWbJj6XAmAwa2kBk97DtWXrpQjj+HRkKn2AXU+GZ1oHYk9FvQvBGmXm
P73PX4OKDOwUx/ksGuIKtHl7m0VvNPcoUPPvNwj6s6tecoThiSncMCGU0JZoAfdt
PviQGL6vvQKfpqXQYIeF5INctmFPW/IiwUSGOUtgBGTrlSWLzw5ayV4oBoUCAHQw
7kk7vhGyD7+X30jg+Xa+qhz1tU7kfErOiC4rPzWkl2ZB/IIcUW2kFpPXZHmvLdBF
7KBvsLWgmOgXGy7dUv5MomG6p3MyCUb8QVOnl5dFrtcmAC0ND0LQmysfzDiGwgi2
d7jWNVHq5t0u2J9iOaCxXK56IIabjMAZk5TzStcPrKkqvVP2sG3e1y/gxlfWvmaz
gpwFJ+2h+lGHZ8w5veR3rxF/laaxWio7I3hNIZRhDILVx7j7w/qmB2DxCDXrvUh8
mNC84KpQ2/qncePJFGDho6ZKN3gqACzlDtdpC0BbYlvcgUHvNe/rrtUuWVSqxwh+
3FLLoWHSdaPzZREN9gtTTy+lVDif6HjopRkDkJxFJbAv+vMO+VGFG7q6iNa7JNAY
Xtph3Z2StHwqjw7ypLlZVA8HLPDGOwbhS8PwNQ/6mKijBXoKPeOBUSyL1ZawDn38
FNPPPDHd0R5RnR9qUXz1gdQgmY0cOYpPF4phZgUGnzQU1Ex0QHszvE0r0LKIluCM
ZrvOc2nFOR6GexBJOVdndRe1k7c6sYDl6tZc5rRt9cRtMD1GX5NnQEvfmmBcN1kf
FNMjJ0na/iOgvmezfD96WCHyUq3ctlHnoyHF+tbrbQGovmLgoIZTIF4pMrDSNhP6
eTI2yhTaRmRIs05Qyq7jwjhOUPQBnSGZWTu7Y4wLXTgt60OFfb5GFXvzPQwj7YIK
XXUgeMtinKTAEe7hJRtxXgHIHzgZDoo+yCfB7PnGfuNZR54gHxvZdI0hHqDapizk
Bww1qvOdx+T0ioXy9klkq2ZmC9szGemiiD/ys3LxoLtwp4Q9q2U6rTUhwAbqc+ZC
4uAMVn4GMNkz+yuud0tVz7bKMKZ+3+8/JjGy4qJdaS3ylvwLqHnmA6F1tKZtZ7yj
aGE5HombuDqukCVG71XPNedxQBM8uCT2k9+Ij/qVNXjeFozJFl2vBUAkyZpn0IsH
zI5zqLIojiOH0YewoMxFuVkFJNpvgs5xRW2qigoPy8EC/Cja8H8YJFQ/OY6J8xTp
m9EeMLgllb+4lfpEHVRThezQSoOm8ZWnuFxE2/WLn35oLQP6I/JXEdqmf03oyBbG
fhT9Z7D+i1tHt7HmCSsme7XSTp7IN8FSRhDqjHNiVARjHmpGfmwKftpLc+Kdnjj+
uOHgDXel0f1B6xLxGZIBtv6Qks8WDDV9gTVf71kCb/B8aB8gmJ/L0Sk4bsFx2YX9
YmPZfx6z0MqK/8nDc+bW4yXbYfo83fUzG8TDX4WYuX3RrTJEljgYTtEzyUt0fSwh
o6f14pQKbFplPpr/l2RFHmlncf7XNEJSZsgwhT/DReX4HwFmXRj99X08oHxj9UDe
JR2pSyp5D+KJxJQNRnXhwoGiPT2JZivW2Njfz7UgDGQGr5QPTnUGhJipo/wRMzZK
aJkFpi8na4Vy65DEKH0frkaxZnxP7wWrsJf+cRtUKAG559sc/LFDlAtjnCmIbWk1
eVJ9BQ+0js3kBCINHTC1PqCLeSzrnBF7V7q3IsNZ07Y/3zxSWbNH5DU+BI36tb9a
f9L9dVljCgd0iGT2OgzwebH4i5co+Oi7aBUuqJXZkVi4I2EzvcMSHy2tyz4xSbky
y7YtYCJdaawcegxcj/WH2cGqM8dUpebyur2oy1pjmus/Q4eaOKhq/w4wFpR6gnF5
coQWID/xdFvqFtvY/FvtpCojcYyX6JuJQj8qV9uGOuaWXxzJ3ny5+/Pvvhl2AynT
heT28ws6NPTqI1G3Y9FL2kotJ/h0couoOSWEcUAIXNdfhDZAhKD3Acbamr4ckCxW
+uheKZEilaKr8ps5zLMY2WlXK+TGm2mxZzZoa4Vdg/VUsJixqV1IsgfNC/uVuOMn
XPq0RtVN7ot6Vmn43sRSSNWPswIvlHohJXWq1D0bgZrI0MQGxCax2NdZ7wq7DVRM
0fu88lkf9mfZttetGYeqX09DJiDO2Geh3uOfjeNOcYag+n//XS09EqKLZWsN+k98
3sLXeZcnNUKORkx5gAsVLlz/nKFKixFVN4Ry6Y3yGMaCWTGFpTz9VKTE1hF0JuWO
eazMnIQJzS3i440MT2WAEl4G0/NbS1w6cYU4eIutWSTm4ejcIseRW/GbI4FriMtA
Pv/4OeyDc31uung+zKpNWj4GADquo5EpvqZrXgpjz5wc5T7xX2APxB7YqaVcxUxZ
zTZ1pF0h+kipCExvWc6+CfQxUea7ZVs3bhw79oYvW28Hd5+v680nn32s2XjCTCuz
SzckEQp7XDU0Vn9r/f/7IXr342B9Ah//R73bz430k5oPKCIhW+IRYhmX4Ri5XA0U
DEKdFUWzkHcHwGg4ooQft+S1IraaPO3G2U8oluzyzWxXoLDWj4NYv/v8mMsAF40X
KKN/35ZdiaLLPEjDFIIAJ9w6SfnnriR4rGiGhmkdR0ZRH20u6sSMWKbiPraWWDQD
7MzCOf5KCbJ5zt2rx+3EfRsKT3jXDjw1PxyIsXpRKw7aKpuzqzIBLQOF3P7/I2h3
OTM45O2PlYqzmc7awMqIIi6UqcRISOrgN6uTdlp6yLincaoeb/RrC2uTeTc2YOHv
pfPPYonMwZoxMKRFwyDuGMRO8s4lPLTHNVn7UvVfJiwae7e/S9mQIO9+3xRQNzNI
CyQ54L12pTTZaJsopjBA6xRTZY9kWvpKeYKwHfapG9TnGeH0ITO1BKodxYv+LmZY
vZopYshI1R0vx0aIUqATqOQN7JvbP0QY7mj+lOfdU95Ac2hzzMtwHgy7vyZKNLC8
GammP4KfBZ8eiQYPlffKOzlpxpbMxsYw5b0dWIOQW005V4Iw/wKkvZtzMdv5cctC
YDJuhHYWI/6u807HxMPQvuSAW5pk5OoJFWuN3SEYcZ5Qg+gWH+y7o9IcLHfV9mj7
3ySWkDNDXaTrXhGlXVhzCIcS0nNfivhUCI3VddNiOM8Ji1Mkg+bQAj2NgKm2uJ12
pRk5R6+VitMxBrSRU6pUdrf95OqD8agixp89Q9xBiy7jla17NeyMvBsaLPN4b2Md
Lb7ehJoL4A3BDjmqcZX2nu/FgjgaLqCpPzgQwkWEy918Gklgv3A8VVkD046nnovS
4P0j018k3ZtFK1zsCIYVXLED9mQh5vavv6bG9TjdBSwTr4KM86AAmcrr8+/r1nPk
Hbgl/n9rqXjGBLRVrcN3YsJQFsknMoRU9QkYpzoNYSlFp2YLhFwYUd3LI1VIIt1Y
L4Qmt7YATdCZKfIscrwAa8EHtn/Nq72wtPcTstAl8C5SsMZHEV7+nyGrDeywetXO
+Ru0vBqTocHxQqwHbJL1mhKSM/DxssKjtHH7uJ1b/VCyA2ZykWXRnqYVsW2bCpQ1
yZ2iluM/TnsovMX43ATVB2+W2JPyOc8AsZCAKETS70fO7Nc2wXBa7xzLecJUQYLe
9XYK8VcoKSw5tiszO8HoEFK3Rn4Snx///9VSKAATL8vfF6eLWgqyqkFp+0n9tFC8
GURDB1vcq/P9uvcfxbXnCw7Cx4KeV5TFMTnImW9zCGH1yB5Z27GRzJcQgRQAMsnf
Wkejqqc21D6TjmJAeSFT9NzVuI2oOhv5rH1758Iu6JTmI5SCDQHzMuNcEex185PX
/I1Xi+ZvnOU7e0jx3HGSCe3NzbR0rOvf8S+ZgZHsiRcyRzBa58omIuhhd0fFHjYP
ieSMoZBByJT4+6yXiApcz8hcXYk8icVIDwpVPBXIM589x0RVGMGqfTaWEbIBi3t0
Apjb104BOZRU9KW3/HPvtwzdaNssVKCQPf+sks7xg4XhbVs1tRHlnoo6hg9sy047
YLEanwM2cOtv1jRw0jd8Zh/XF7DAe6AqDflhEUa8PCmIrj+eTA+GpiPLtki8XEQE
YZllAtLki5l7PO6LfTDk/h0FYGVUu8H42J/WTFM/jYmOP3QkjhalIEjWRk2cmr8i
6HoArLfJug+zhYmYQSOvr2gZpum5qXINQ3hwbBcqpIvnT4jM5ZLbY9rlW++cJLbo
CUP9J+zhdpB2WZp1c7+F50IzFdzIUa2WqIuRq2428Wq6kzNb4vetI6C4lek+FZYf
c47jfclXGapGAYy7ctGGGHztDwA3UV0OlHoXtmW2g032LApKU7019q6F9A+aQXca
H0HPA9zEYd4zvBvLLp3oNlFxzjlXZPkVm/Hw7n/ttOBB4TK6vT2IczINcKG6B1FB
QCJMRGfRUOpif6JZbXJ74aBkwOF9DUW+1UoVHfJZtLHfDeZ3jY6riUXmrf4yq9rS
y4hFjmEKmb3iXocSBIuDZdNuEjt5OfJyOKIFuvtS7g/yL8LtwrSPRP5wNxAyAlh+
CuuhK2zAKj/xfGOsRtMWDlHah90VqOIZkp7PeFEP5LJ9vLRH3RuHM7dKB3UMzbLB
xXfwYsujxFOZ8ObzaQKgku3uoy5VIjHrPvxyqTsRncRpD1OEf8qXCfW7VsOAgLNa
xehqo57CGWDKA00LOdzg/OF1+gDSmNDqumKI3uhaR4VKRmZdE2F86C+rcRIVVJE3
3weunjTuWwL3je+Lvk2yNcXuXEuCAbr26RmcckKFYxStIPEBhvxHw6aT4AS2tjGp
qdfE0kCVJUeMERA+wdEvFLYdg/nyffdpGXhq8vQICcphqbZ8wGA5hRXd6wV3WiHi
WARfFjDLof0xrWrjmX4lR0agym1rt1gz8kw1SQymZwJ/zYtZIYXvKcnzg3WnUtfS
scikpnyyhOJQzLfc6JbXJkXyOU2pHSWxT97FuDztrLF8rhYWD6dnoVE2F07R+/m9
fKtV7DuO54Acg65jvWSpLwrHO6VUNCUPWVLq8iLYfJ+7pqMHFOHdE+GDKQuzOYiI
cv8XgIPTAzhekFQq8yguskbQ/CdjFoBenVSx4BdZQTclZUr8fR1Zvjmq8WLBqP0t
p+QjAPgWYTYsYgipwzWQC1cZ5P9BTGSFyeCRRg94EdjE5jk5U6ADNy4UQVYpAeVy
ob1NKv2T3Sglfpyq0OozxcCyFLkfbJp8iHHzj9kGdSvBtUdgtjoWPvjPREQMKtxC
Lr6hlE2Lm1rVcRdwtjqgb30pMIRSMMGOtLwV/60MpY042mSav6SF8xIuNVAxwEgd
O42dkVjcHdWP/AfLQW6J5JU17tJqSaiw5e7wDR42OxzmYYp6fZtDWsVwCvM/CvE8
ofHFkCkBhHv1Ie8hJwKeXkAVBPczTdLQzNN91cmUkr9WPGWxEpsaEAS56irDCbj8
O6SVvY7qYL4kjunDYwin8HFlvSQBsc1ReRoBi4yKGLV6iVKC/U82NS1/EhrvmcxY
TUQ8kqwSDtVsxVj1Ff7fymv41ENxXC+6DVdCTwXKTSwP7ok2jKFAwd62fyhMO1Zu
nvizayuWg1Am0s6zapuojeSNtQ5zeNCOvvncnJ6AmGdzQebw3Lcoa6p3zbTC4Kp9
7S6izJktWbWT67U8JAwNXq9lakdy5tGV3cB9baKndI6XClzOo/3JSqkpEDZO+Xe5
bPKNlQndVhv421bMNRxMKperc/UKY6EJ73TRzLOmxk8f7FHswIaiqnp7nVln4kAS
Cbb6PLu43P1w72s/hR0MM1z+P9M580i6zfZS0Q+LP3TQRf5pLaszyFfWSIgZV1yl
9jijdCgjHYLaMT1JS2tfgpNJz1hLPSO4hE/oV2/ej2d5AXzoUqwps7aoo+3N5plR
fHbNzj/AZdZ0MXvt/DFRE/0hMBxy+0sOkxN0KsLIl87//PFUyrQUeQ5UJNEWf5Pa
8OGd9YZ+AeiW83I5b/SggAFg//Z5mbwwTaSsEGzlr2OTO4oOnFYQ1/MaJbIEUMv+
Gcbrem6zva3aa5U5sgqtvaxIHwtigF9Tz7EqlyO0oUmBiIaL1WIQfeyyQj+Xifv3
aEtdHc5XRx2atYb3I+70qgVTZDMX0DHDD/PzXboaSj7Yr80mRhAHh7qvhlgj2DCT
Y7wLYI38ULgkdkASOzLVR2rJs2omYShTcumzRl9trZreaFMLy3WPHGoxOPiLkgPn
DqF8ubgqc8aM2szOr6bjt1YKyRoPiyKyPhRnMu78XT/9xpxop+S14lhs0SSbROMj
zuP9DSCL2A+etofF1I8UrxVTZmOeqHwzV9RttLffX27ot+U+YDk6TbJR3yxmbv8R
IQSJ8AyhHL2TC6sVn3ZHFVo4iIYy5f57oBTeziWDe7wywAryhxhcISBkKxGF9BdN
9sX6N+wCIO2QG609TsPG8IdXaIw7w2bRxDEPyqtZePAIDoKRY0MliRodzMJJcR4u
a4ZPRfOqwiKMjjuFZ4X/9m0pTktgOHn5/Gj7JX6ikkj3nP+LuFtw3r4NsEU8NzM2
w3vzpbch0INzriaTt1rLuWlH6eep4tMvWJwETx7suRCJt8z1YPBRD+ulj1KY5/DP
Jk+RSS0NLTHjBKPLXABS3rj7uvCDfD+7FaC3xN24CI46lh/GfJzZ9GTtVyxtOEjB
OdBv1jaZhpGftMLX+aGwviP7z4GblIGaGnBmK2IHeosMLEHIGBB0MizvAx0lR+H9
xchChDlYnEetQ9zyRXxKhxosopbqTFrQSUc8CLPSpwNRf3vq4miquZFEbWFzrM9h
bbuSWjZOBWcO41mM+RYwlPASTHNczMsBgHdsqA3mfPUM4ou78b8ZNaqIkKKfdhrQ
OR5CagwHfnSEdAtpLcn+u3TM7VZhflktp2hTE3hd5yEYmv8eeLbHFquwdON4Nsz6
wDYo/XndY0Wct2V9+ZzOmvY4eut6kosHEFPG0QY8aeGj1CZpZ++Ejj/GY+KP44ol
2ekWFPV1C3/3TSW8e0DUp6kcyVOxzur23nd33emgMTRjiGVyatFu1gT4z3NkeBqw
52HE/sfDXcJZmhe0fcO1TDcIF+6PQPdBJO3hDkLwdD1V4wUmAHzvkLGgIu0CDLQ2
y/JaNwXUPS3oUpoJuYBNeEDvIIqOegjbg+PfKvXmihMhIxnitRl49NKKzJqOMF4Q
0aI3q+MfcyzUjXBu7xPjRGALWbfU1NKS42m7GiD0IEKbCh7SQnyNlE2BVW2WzWye
F/yHF+yT8KoOncgIiiwSRD1ypshzTpKf2e8BWkMA1n2fEZPdfrCgJV/NdNY/81qm
0AMwupm+Ky8emK8lMPO8a9mdhibc/VVTae+w5C5TeVmmnv40hFQwNV5fxxaiwKIq
ByJHGmNFt/NTUB/1lRrKo6PkthiByc9WvmjnFzQ7qjuaGU5FDvNwuafDizIK/V9v
ER0mid88lhFCq2hIlrxNoBfdtZmyXBVEjqxm2MnkBOsFzWrgOakb30TskVvFscw5
XiPYK5V3SKpaVhReuAKJ6pGntPZQfIztdUlYeDQzQ9fIa8Xf9DL83YlhCUW3Cjjs
jcf7QKXyvLKKjZChJ2U5QHwsykKNPqhDyMGbWr1G4IMBRR0edLdeHxyfjwYmEr7I
gZDD6VFeOjFJ0g7CwR9bT1ozSBj6kaVu6GbNhZ3jHS1HIFk03OpkLG2loBAaxmLg
M9IEmPNfwUHKL24EAIdeKlRK5tGn05WAa0cPoz+uSiNZsUrwzzN+vJpFh4SxXz/x
i2M1JptM+dTJbkBssDib7UbBwa7j1J5eOuiliOSV546suIcSb56qXoDonfdJcbF/
4tsyN6jID5nPc6lAOocNvLv4EprvtAsIwiDh9+ZtKsmP2gU2V6tCdxPpBirv5JQM
GAKv+AhtCYr+PfwT+nuKejAYgPVRo7HsGTpTncBl/dlfr5EXqPWxeTWwFzT6Eztx
M5A5EWOwYszYdtYNcMCRlSCQ5IINoQFK6HO2YV7C7Qzai8sEdgeUuuzLaJifj0Kv
LoKJk7TmeDR8Kbi/b2n20GB51B2WQR2kz/uQK58B3F+N0NtkR1IHZs7XKKl7HJqd
moocWLwN5XUcigD4V1se+8VbbHBpM/Ds5266OFx/zwknPo41rLdGMEI+E3S1C1GE
ZbF/yOi8lvSrxtXvwIkSkD9MdXGi6F5zehU+aCQz2I2F6zDOztK9NBvIIBwFd/k/
gtRy5RqEeXur8LRf7034fuFhWESg7vurq4sSmQkOKSc09c1b5rWSxboCDo+piCFc
Uo+nHB8vrE+VP7V9NEq0nI8mFSNrHnciGiMMwZrQtWXMJE6/AxEhztvrPAP8kuLb
onYNFsr8vUOInZsqpVktcCqWT5BqNNCYz0qLRXfGX+PPZqNbgQyu2gXftwidpCfm
+0CPMsvLA4pS/h/KxoPh6bLPaCJpo3rYeJkeZ3lwDLFvwqJU3jVQ65kP/rNsWKeN
GoL6gmDjlLWvx9Voq8FZwTJ8cQLNd6v7SfAKYyn3HLK+GGqehkDm6PyGvLLskiG5
owrrPJt+wIN6e8JtDdeMnJRskI0lJArIVfK7pjFx3VURQeNo7QGEIXNeqsXCL8bm
4vkBakbJbHmqX7hb3HPQQZou5ZS5tOf02v7fPAXmyyplJkooAe/R5pDRkRQ3ZV5Z
nKvKqNYDtP4D89xp9bxuORpNb2blvvf59YYfFyb++LhOFee6cpKYvhGk4PgvTo7/
plVZfy/Q50x4t8968UmrGqFX9PNqgvGgqXKI2hIZdhHyfvTV3z4COsbqyDiL3Vlb
+3lSwxnnE9SJL5tSexcWkGGHyWkhW12oxeWnULGDo4OozrSdfTCOh4mRbsfPd2sZ
xKsfd4hZjj7F0cjxzAHgy808wCHAki+gs95JciROFF8FxC75FZZeB5aI7UN0mjH2
FsVOhmwV3pfwu9l3HdlyEy5De02+CZ97OvONjkNgT6W1nlnJo9+MtJsmfDzvtOiS
XRrljPP/JTslTvQQ7+rdyKQFBZEJqKyj3A9Cd93Au8WuD3KIm3j4PKRKLY7ouJyq
38E66E5ovsbrEnVBqesxGuOtmiZjozi5UhZek0ATgH9f/4FJ/N5smBHNfVjAVH86
lO36D0ZbYKtHI+k/LZJqp4SnlY0HQQF8I93QTpmQV2TlaCMX2W62he2Kztl8zMVi
PComNkQoh8j+cVqHdi5ONMV3z6D8dTOy+UkeRpu3wdJeGpriM6GZxODQ0c3aTfxU
23brSUNhPOpuZp8X6ggDjVZkvwVD5gbNqtgb1BZsfrxwzMSPYihafEk31mLFBzak
eiQNH3Q3axbSnkRNgpHi2a96nllk2qQt8zQFBrtZ7xwXxcGhanbDcGgDcASjtjkQ
qel2ubpJtbiw6OjmoEFPiNI5X1rG634hEMgefTnkitNIStzIHzmH3+fGQ+DbGWt4
DEMxAKLDcYPX6JMajEb8nQX0EOFBGBuAGFKNtl5p86vAWHHT6DMy9We6BgNXldp6
NwJNyN8C8rGKXVcl7VLIw7n8uoI+DLKPzrF3VR6KQW7bbcfjhrSJH35nJ/pK72Ti
WqvdsA3mRetWQDvssunMF4xECgLM+HmL1syaYlINplV9vRQdtEFNQK4TDIDdiXfD
bCDveESTJNHwF9lrlpX2EaMBddIMerdTPrzFWR5/wD+wb5M8946a1MQE4uNhrqd8
xbOzLMl/y+E9UBF7lojj7EurdRgAlzQUNJihXVYX12yPddLqdWcsy41gUV99BNN9
BXWtvIUW71WQAz5oQHlNN4Uzu7J8Oz51YeieEwty6AT4dmJ+n1Tm9UywehzuoMv2
qxej6cAqczu3US9kJ1gSHbVpmLHe9MJ25CSApWTMEJ3KVOFdX04HblY1ANwqlnSv
+xRh6CSCXSLPN0liWh1+GiYNjJEVQToUPii8xMaqJbiU+A32lkVdwlGPvlhEXL5B
6o7n2/UOUXDhlnk90howpe1bH3xqz+VuSCVNsocl/EvE8DRBXHMuyTijVXzyRWms
tb/8OQ+f4kJ5bC0YgiUV6kCPdxlSaGZHqxnAQLy2K3wqj8GCSSVAkZdwia+6ThEm
zqMs6kOGm6kvzgTuG1Y0gT7YOAUJV9pt0dPCGzrcLpzvBH5A8mIrzvDhqTi76tnZ
9i8wBY0M92zt2Ii2FtmHKVOVpZULYjDQiignN478RfU8zEdN0JYzPHzNJm4kAq1p
Q+9cU0XYFX4e6Wyf5fDcFRPCvUhNyfb96aSNVdjIxzZNpA4LnLzIQ2NP0PrXJKI3
tX+4Eu09Ck/dfktoGjbP1raDo1KAMQ6FJiGFcKmQlSVTBA/xHP1qPRPtEV+hTB2Y
/7KsqHk2MlKwqguI9YTnTzHu7QHGxe3uEZgkS56QmkQBUMr5/Bc1hfR65Qw93RGc
hYNEu7cLfx9XB3xV/QoCQAQ62bulWX9mITQUI+J6qbjIPrZf2jG221VDHIDREe6s
G9etcNH1OTLeCKGYuwI0xzaOayJpkU4qNYaNp4leK8rpmENnDYsLzYZ/Mi1onWuZ
kmKQvIV98xu+ZWm+OYEMOElYaWHupakx1zQlkkQQqtsgpPfMJsaDCwkNFbozm8De
R7VF0BqjHZYPylLXgXE4Wja4/M+Aipwvb/gNG47IYGvaRO3+0K+sFoeIOjJJtlmw
b98TX8B+es6HnRvcXqGUvcPfXdIx8QSPndbWrGE5m/VjfS380huVOqodV0Jr0bsJ
wp6qjvMijVeo+neWiqTw/FPFw1HYUFN+DSe0oQn0eAuWrHCbfN40zVqdnW17R6C8
hJI7z34EOa4mV2VLJigESWx2jhS+J5yIlxlTFK1+hKgOUamB+DuCSLfKypUhI6Ao
BB3o0hmpDdv/tQZGSccdWJgFx+B2dTIFLgA3EHmEtkUAIaasvbc1EyO+sq0hgHce
dQUsCSaiZ3bR/NIPZB/wGTc8f3Pc+2838RKD3leabLe9hj4iL1voWuA/eAZbTsPe
/9OnIafiFbBXO5vAfytugNKpNVcKsBPI28Jw09IbT+3D1rb1XNQ3cU8IG6tL6e85
b3uXTZN0D9MnVipnlm/fOosDmBJTqC71h6cwZJYUYOyyrY6tptdIjkvJ93O1/zNO
ZGR+4/mKeTi68poR6R07kbjZ2elVaYxwi0UJTNAXhOfkt1Z9ZM1kOPhcDg2m6k57
+WsOKzws0YHdVGDqXCT7khsf75tUPYFdxzQFgvUkVPriJh1B+K9fW2T96lDOWqP5
nXU2o5oMQmdZu+GZAbZIgkjoHCkuqjVVXYwp2bNbRps5/3ylS9z5ixMF/xtXkmog
7fW84x3IxA+LI0hj7XNstgW4pt3BFjFk0MmdFVxKKZ/+k4qw2S3OuPFizlC0p0DI
sIKQ2xR9XGRB7bD0+L3QuqpbyhX8xtbr0tf8LYbVvNEyjPfw/w2/V0BV84w4YDre
sZjW/e9rEGRWzBVyAiTk91+l4D6hzlgpI3gjIC5U2QYNZoD9ZYb0ERLhWFkzawmi
QXNcO0thi+ts7fGXgcIP5nuSOwxeKnSO57NpzX5xXm00eKi3+5mO1Mp/MkJYDG8A
XDnfHVhyzrKV71Xgf9EJCVOZ69UDuVm1FOxRP0UC3QOoXI9Jch+Izt3RfZf0S6Xl
7UeBU1LaYKFp979pibI+pCMgMCzKtT1puJA5ujSfVpjTfz8hp2d/rTJ+syqqN2Ol
780oU9FU6pXK3vkTSywJe3wsVecVaijX+porzkhRuYLEUTlJ86J7ZnHY2KUvr+8e
ZGeBoHuwcIOcTD/6bMsw1mL8mUys2q80y7oemPpU8KD1gmsmpofUhILMTZjSdC3/
XvsRBMoDDDrxKNxBhn6UJ1vcPHTUq2ZBB1WC0R7+QwAP46yUJP0TiPkAFyjwa8Ux
0pPtLQMvwhpvxYALMgpAHKCklYwH6qYmSStNpkzepl6CgcqHFLoTSFcABoFHf22Q
A5FY9izgBpeXk901EPiG5l1N6sQUWmIIG3mBlyiUWpYYcw6n+2gqbhQorMJUYfuq
ky4aCG6IxFWEpaexusKPTGjNdZ/zksoM/YcvY+EfRzSYVzKRGYGxkddC5pj4DuBn
keSpru1/6A1Di5E18s0h0zhbyEKcsTV4BD4SX+nPPT2FRcaUO4ju17KkKUtNy8FH
gIGQFJm8Idw4zrqXI15FUtGwsX3LgAtnN21Om+nzQhQQvUsLG5vg5bg+Utx0BeMO
0bl5weGiZl7Cf2kGD33xC3zo+Uf7/YUYvDBIPP4TpAPq3sQDdWhGCGHiwhSrF1Ue
RCafCy6vpIR/tLfXGKLs5/zzqJylkTYvYcvKaQcjSLxB4TZCzqyXZcuczgsMHoqV
DK1FKTBr0/HY8gqvlvPcNOBwl0kakLbef8P3r554UxuKd/I8nhA63EX0i3ztYBDe
WFkIbFOBj+M62xTCmj8Em1JQ+DVXk4UaNA4avn5GcsoA+Hb+qujIantwsHuCnADr
3chE92p4GOkkpGgpPgGdrCobGhOCMcw/4qt+ugcCiwDJhEOMGC0u/p+gSdC0fgRw
I1ypo1QWGCMDPF2Cl87SlMVc57O4W0zKD3WPLj1RRgboX48s2xYnZ21Epdu5DGaS
3Y99GJ1S2W0b/+sHqkCXMC8EsoeEQvAbBy1yjG/mYS3swJ1HlAFEq+GPkwNNWGV5
Mmq2jDthRFQmVuTP1tjxZXO1c5EniNz3gtbq0gBgQ4lnvKd+24b2ylLWPjuo6wXe
38o4YG42h0FgQHOb2GbGXg+++9LbFX17JQd8fY79zjow6c2fUiBtspwJKYPfDJ//
5ZJGMVixfvxjzYT84hHwPYT6N7FVm1fctJUFvuqnUHCt89gkfyboAxsXi8zH8RM3
5vT1a4Jo7dpvqePb4FguOFbL9a5EJPmQyTCnKUToFdEJGlRlup+ikeSZjbUwrb3N
FpfgcnrbVzaV985HPX3M5pVgNIidxIornLEI0L0LgLmnpCbcochcugojXKR0IU3y
CMZfPp3Pl74iw9OevqJnirXzAt8xQuAg7OoRIGbSMO3jHFmp9Vm/yGqcAd2sGqdc
noocaYPOWGTLKF6unxT5J0UUV/gCOuZNSUCRYZvICrOXua3UuOdquqQCZaL7KxC0
XNSsIVwkSFRbG4W8SPCOpLOcqIY353Bzsou5RjdJlMnUUPoyMkdg4WueOVRPU0n1
9xUgvi5gVNVQv7ksB1DVjnAOw1iLnnGFMxl4BfnlDAWnY50EKaw2j7AAqT1jSG1K
oSzyuDQ1P1RGIgodW8+/qPlyUi72SDUNLApymIhRYoHV4qZBm/MBJneYXHATkJR4
wifGe0eINevMIKvdBS7ERp941Q/sohBFfa7LWBmyoQxWZ9DAvm0wRBc8H6EVrO92
yuPoUA0fphcsJw72fXgbwfU8uIWjYxrAWFgPNpgiK965pCKHA5WRSIVnWJKtig18
cNNd378zVZh69nWNmuIIP6HAPRbzLF4GmntObbJx/J0F0FupxTy+k1t39ZLRHX4F
MJOrGZEIIQIUnVm5nQ1t22N+pewTIsrkafbq6GUD20TMVYH9cs+Qr5aMcULhaGjJ
BrdSQ+Z2YuPDgXcGIT5p191wTI5E7fWqZsSqPr95roySNAXSOKFQchchEakoaj3P
Kb0CXjJ25DSozNTqNf6M/6iVMpKZ02VO1CrVeo7al3aBDeM1BTzF1n4R4v0x4cga
96b8OCdLxG1+dpWQhW7SFOkf/1VFSKrpvXZ+eVK3N4yjk/nCgqn71FXj4Ha4kqvn
ffQXrVCe6fLCCAINYKp690nijra4T5TGUXGFJb3wp9wN510rdu4z/Oxk+6G5xT4/
Umfxd24UsJoz5HaK7hc22zhCvz/s9avTcq6UiPdSfZKBpE8xvmq1Ay5YsJSrAg33
z8MOMJfHCO3QmK01APUeymBdm3nBYKKYy/aRHSpn0G96oW+0bgiqsyONjhkVcABW
z/dSTHxhl3zBq0hSNvqpQ9NRDBipf6qL1WFhbVPw7dVDi5KCUv7p+AGRdoBnWhUk
JC6JaFTBQxRW6KtH6SK+UAwrXQAE9lpTmcbG463EPfHOptxkIjZhRZR2g/q6rlwd
9Pu3Tb9e/ajrizzIcV+z3RExjipuOaqyNcZ26yqJFUW6GNdESUj9N6kOsVvFq3pP
n8kcBOFtEcaloGPXt3gkBoweJbad7ToEkKy28DwUGwvW6KqQeY10YTTE4oeCRVxz
T/JnGIEWhO7QwWGd6Ix3zojA0qIbPeln9AHCrTtBPpnGXKauHb5rFWqzNN/EZFXU
RUj6iZRTa/lnhCCV1Q9CIxkY/88wH5JF6SWqoi/qARdqeC1By71fvayWkquWqWrF
T10/+eo9AhNe4MV2BgNf0Rflz1P7vYtjNWHx2bbEPipoaeC0G6z1ti1Y6y2dsAIy
hoxmO5mCVQY02ptAZkUix4ab9Gv6c87eNr4/wCPe0pOskwx4WVX1G6o1TMbuvzBg
jLZx0/Ka+YhKOXDqkjDUEHod5s/9lw1yQpCZmHuZHwFfJHILj4q/VSDyPfoQLzvD
tj3tqdDm/kogpOICPztzWkCDxwzQJEV3yDRGsa2AjKNjLyBiH/Hvj1s5HuDKwjQv
5fjC66bzJyVKksBBMzb5WcEQTEipcOUE5PmDYgdamESniYzaCicCqjJzLcaFKUiH
6XYbd9aB/+VyyW0EPWsPWI+iVeS0vvvCKtzdUgP1WCt9UCAj7OK4SQOTlLvWg1hT
BzZmEXmUN4sjpwmL06Ej19JOHh2Y2RCY0U9R3Pl5bnUjqdXRcm/Zz/gE067hrg2S
y7+wMGYE/u1m/+ZCkFHOWIvkZQ3m56oD1gLChDodGQQq8WbZbtdiHPTRJDwaBCjN
IgzsWksSLbg6dFCsmyxKOVt9Ef+uhyNUlo3FMkC9ZF9K4nXhBkqC0SlimGTOPiNm
fUKfN1xtTximM4iAETeEATgqz87bma2CPE+PQ8rcK27iBijTJsSA7vaBRGt7nvH0
SH5aw7hpedJRzjqEclUPp1AcQRZ4i4gow518iqejLzdtnwc6IaQQIUui2tWqE8HN
eD5t4MXLBpK2ISsVCXFFNmQkyqKq8rinqwRkg4UROKhfTk2OR5SfhUmOAFc46JHp
5dcdW0y51WdCDs3W4R3ysHMPxMeGXSKlIPUPryAMF+Y2bgZoPnNWmPPyOc3gfEPy
76b7uqBkSvnHL+eR2xn8Hhfsu6v1/UlaI30vGP2Qney3OpRWwi9Z8NwM1dUdyNUf
W88VrqymrnJb6fLIwMGf128Rvh75HJlAW+e7K3RJRd1DrLVyahHHP7ObFLH5+37m
aNOvxKWvzEqaeR4T7MFV1JHybmh/FgSoY0ekiALhm4cijm1v7xtY7VNfM6+9FCYQ
BQe1EkaPU3/GQewVSkiCWEIJ50eOtiTdlEkjIJV+5nzX6ZNaLFggXm1GO/tMoN7A
wQZWLKmorMN/0P5kYcfLWrIfQqLunYZdPZyc47JODK//gaeeUH6O2v8yKygGVHlP
YPM4pEg+z91itIHIs4yth/BLVBExV+TAjAvmEpsEmZI/ME0ga4X9/buoRhW1tJKM
75HcX5lxWy60l+O3/IGeYO2zcJRzzdC2fPqbXXY5LCNEtKiVlUlO720v/4wMzRjO
m1+rJi0/YBcAWXwhh3w12rRYKIQ2WqLG3JN7SSd2ttUavZ0bDf2hJPcXIDxMg+EM
Akpe7GnT1RzJ9+4mcljJDyJM1pcR2qPinQ7TEuY9USYQb9uudsii5BQeitjrF0V8
VwyOm5iQLtaSGSsfi9vAmSq/tsGmX5uOgWMKX2NcjP4fZW5NjBg1XRNyTXUubDsB
7Ip984JhO7nC7yb/Q2yZDidiVU8GDIsCIadJa1pvB0tgqhTsXpl65C33uqtyaIyV
IwUp8necXfPDy9Jxv288z9bKLjV6OfDaOa2NOJivzRS9yFZGKvblPswiayccdO8v
HIdBYNbQ6yPAJ3jIOgqFgu6dpeElEHYpvBXy85nt55s3QniEThCEuPpO+x2w1YhG
PGyPnJaXWf7QXtkC3sBLvB17CGeLFohw0F2tRMwz6M33lNbXtKRpJdS+HZNBLpsQ
ivSLVK1cUYoHyPutQpCRD6Jr6GjI9Xn0PsWj9IMc9dqOqDMb81DfpDdHNwEiIqvO
BNf4IIkxQdQIkEIJt0LumM7H8JVrir08i7NxhcRorOy2WhbV7ImQzVUVO92amPv8
DgLTPv6rFP4/ts28x0Vp4Z+Yyg1gXOkSt2FDuab7rBn1V3nB+BedQe00ldbNTe33
+emWSbf8uwxcVZFfMJ8LnLEbEky1PQpTU8fvHz3KDOdwzjStV059NIYBoDfLqUH7
ryiovdGJTRpdq7sv35KE/jWL6IsSpJeKq3NXl/zaJEI+QwaPeVdfu8ExEsvN2KS1
ycNTtLXqQ4KRgdXZS8dOTvEcMbQFZH86YCDd1jKiWoFz6xTWycSSywtcquDsdsMV
M19TbOs/icNe+BgVbY+y4OpfT7pOc5HNQDztOdrTM0LuwSw3aKNxNMj6aPMkgRxK
hj9tWkzPzu3cU4kt2JjCSg4/U+l50vjJDO0tELQWqnebTCoYpQ08GreGKyflDyiC
hgRgyfJ9MwW1fUMrri2xZ0tPFNslixD2axTXmtK6Nf8UZNEXUi3pEvqceDKgrG2V
0ijTbYA1UnErJBfTzZnRPRuYlJhUwSDOTfBv/lB08Qu3Kg9iZMxqnvAeSji98ZbM
9uSYfvVDtmmzz0rvxiGczaHSDl0WsYhVIRSxceIEUPWoHrDPDUGBdAuh+ocFFjx3
tHY3/pbyKKFdzae9yCHPoc8kjt9ukUr+KbDjyWcWgUrN8x2beRMGCSxMSzPXvYBg
whYETciwXiHHolpqgzViDbtVJ1yoZSKDrK+PhEGfD0QEc+fyiCIhMHrSez3R5T9a
9rcfrQQDaMz8zQgzz4/IX4MxUeJysiT2ctIu/DQrV9WptkmVcr8xCRWt0JeD8TjC
GGqB0AbDM3W2j5/A8f5tIhRLFXciov+Asy8yl3BciJvbd4Tl/WFRIDjZYcwtQLr4
KyLkIohhXYqTTtbNZOMH+tRsylnmBodMlBfPXOmrwdnV3d937s+8XmyDa85YZQB7
JndgbYytsJ45bNjy0R6qwrNsF6w50yVLlKv6OF3cImsuwfM/4I3z9mmp2vS0oV7N
bsuz2lcT6FtO3YGCy1+VCqd+9VaYYpi3uiN2Qx8C0cr7pjfna6OoltOoIhbBDfyY
4y8YLrQCtgty0Ohx+wuK65y/NDAts0uNLIAtNVAPCQws3XBVYm3nOOByuvyDKrTg
BS5SYWRBkQLAnjq8kTcm4g2VnI5HY5Dx/MAPH0vTOHXsJQbsVQSacaJZureaIjI6
l3vNLwcZepB6lF5tnNa6I3gXYRM87Jy0do3JEWETO+9rMoyXmKxhZZXQWdWYOxvh
mrPVLnLfZaQbiWiYtm0YrYsa+nqLTKK2cMboxUhv/4/5xzgaKxg3HyLNP3DkcQ6C
vshzzqMwm1o/8oEu11FUcldcMAe82WYtScxaHP+OdBuau4X6Pufwgiw2KwQtgtPx
12m2TkJ9Nvji5EyQjPi0QANdkFN7Fyl8wub5vDmeloReKE3q3Pf9poNNtGveAsmj
gZEGYd/new3NdRYBSJGb0OisT5tVxw1N9alFUakK8OFaq9TTH6nlLzvSaTmVAClk
0aniKyFiH3Ohvibk6LvOmD2WEjFjjFkZZE3jmlJ5Z0RtFDZfXe2KiigQ3Py+t269
4gC8KpI3zMNr68pYigZ/AOy68JM/lTb5njf7KBREJxE5kV4WcvsphEwofmQkuyWn
/Xhp36fi+rNgakCm+bAexO7i1b2Ef9VzW0jqtg95C8PBt72CyelRiV1a52a6tAz5
asjKk71F+3ekBXXCyyvl1zOGGQEHqhqWtEGJk+ejiqKOLzeRjcBD9fd9b9XgSkdT
ruJcrxHBz72WobXclOnc7cU31I6M8TRb5elUkMpDmm6aYjQn/jhsUsQ/hAD3SM2N
FgMOdSTKQTHjISk0ndlYO7LR1liW5suz3h+vZQAmxarY4+AgQ5KbaCFp73ZTb5JI
0ba9gAPtsB8qKMqpD69pyyE/qAid+oP5DEBLsl1sRXauKihPyVZY8PB2h2+0fpG5
eV/4GTCp/Se/F3L8acx4Wo+NzdXc92PhtjH9a5WH2Pi9i4/8ZneRNpeIXj9/AESF
icNOlEPNZafrdoKQvxLK4vVxvziiMMFKU3yVi9BV1Y7D/IkhWNXX+MfIVkZGcCFn
noosSxZxLSCbDcT0BNmS9epHfMRcFwQhVSrpLtkn9OWbZ81kXUReZk3M4rteO1UV
i00zHJJYGlELhSTKQU46PMFQo+TI5XcLsdPzVQmcw+wlWMeCMpIuftCTWN3eBbua
DCrBX3fkmszN9OIDCC2a1XIqZ1wdQSbTrEjBHhS3PMWM3MgbIjDxSAwiatyXvgtS
hgTtDPPAzG0Hxfh12LY3zBAvgZM+ZHCgfC2BuZrJJ1K+A5GruLgmde8RtZjRxgYw
cSFfGqHKSJs5XEzCyGqvF307wDCqXquxL5WKhPszzRRgUJW2BY1ymh7FcTz7W7WR
RLUklonmeU4XJlPuAsPuGOYoa46uWJequXi45HJ27gOyt1Uq2iHIE6Sp4fJx9VHh
I9sxSMBhYBs1ErIuVCxMfnwRpEdw5KQ61pQ51Y4dN1hkhK2EVIwjdRCK1m37+SLc
pWXygWGxOBfcqR/LPuF5Va4mog0DvEVAN+iz0bBswZFDIYehnfsM4BNHJqZajjIH
xkxQVW2dYOetrXqQQeiE0Bk52L5urm87ri609sPAeDZ/Kp7nVKI+UIUly3VaKuZ8
i7NyicOEVJ3Cp5q9geAN3s+4XzNstIIVnR+ubF7JFEuYPT9MZXjHAhnX5MexrrHe
07+0MRhwLctS3hKcqCoNVCYTB689zTEQS/iqupVHTp+WwQ+ux+2bY5qhTV93olMZ
1GlMFTqz6a24xgRPvAAHqK8TOc6A0Kp/17w//7SKgBUcMgznc44r8wcxL/jIELy9
HRzjaSUWJLzVVCDVUPZmLejsxLnPXmEi/EiKTGDFQzZHZwNDTDNS962SOfPEZoZ7
FYp6o14zVbrHyDpakmOU0wDpLCE/fd9an0BEriA8XrSDwXvoziez3JEN5FW6nGJe
Dn1OPGjXYf/I0ZZWlCFFmOO7J0YojuAJmF/q0EmDHFycEGawpfzMw7SoiZHzpKGa
84Wj1dGbhhOjmBY0AS1rauO4jGlpzY/3sCzpN/nnr4/2mq88T20l9NP5uI3EIgAN
ztE+gRR99Dy1eQvb5uoKOmCiND/p0ek/gi9aPOvqvZ3IQZVAB/kl6cOG0mwCVJnQ
qMPMU0NTC/0QvKKCsU5Fu2GmVkuTEbBGqcXq8Iytx9e9WMef5rVmmnBWJIuB/eP6
4KfSO3y+J0LnDjcyD5I8TplPNuRtpn4TKlEz6Va336e4ceRE8ptuahZPrs+IZFv/
fJF/7IN1MPHlHz8Eol5LSDQc7NCgrS3N6txCM3uowCTtFKg1ClfU4xz0PLLn5Nsw
ayl4h+CzUB1/smu1E6xN3b5lhCDS+jdNWeKjTgzQmC/OjcXVM38s9XxOnE0WeFgz
iLaqzfDGicoLkzqgqyBGWgctYXj0PwswrM2FwcbD6Br+IiWT3oi8qzJgpgIuzTlg
1ksPn8gemUGschuR0OG8zfgZTXph03NtOsknZfu2IRLUl0KWLA6yLrK7bu9YFRPI
QodXc556s8ZlqwGZmtTSsjZ8SOcRCVlB7ea/WJQSxu3yW8cXZfD+Y/sWfg5JoQIJ
6Hw/JZqn2iLi16770q3DuOyihG5MnxZCDhJfhQRQqXJ8I03UmcFqKpS3oiKT01Ux
v3wOdPTjJd/yIthNqvyhInUbO281bJOGo+JTm8CKWr5uHSr2D3/CDgz3qnXsZut+
5/SEqfpUt10UR0/qmEo1xYrQZD7XC34vPJ3NoxceES9UwFEc9UGNrJ4TOIbJEMjE
Q37YZ3gugX/02Ff73pCXQWRu+TWp82S/vpEMS+ogeNMoubdyIsqOX4fUAXi/4Dn5
ErGljB4nZtHQ+avrtAQ9QgjLeqE8xtJA6J9Yec9TIA7ILqSqYjJcuVYWYp5fQvFx
0kkHE7KpLsk/ykd9j3M5zdO0ET0whd9eFjeRcWOjH/npXJNuARkz2GNuV0JdbLLz
y3ZUEhqO/Shi0WjY86E7fZFhPSZFGl7gSxOgckJSQbdxaLtTO35TSfzXludaf9P6
dfx5cK/DlnpL+AVUGDUGpcBGXCAo2VVmys7OLsAF5EwDMAulsxRVhZB95l5dTHEM
IWNT6QmbYmx+4DXkWRP2muP+5deCfm9z7pynoWBaGjBZOLRf8PWX8tfZOFqTgdhn
YPKvApAoJUEwAeR9uX3jokqYo9ZQ23y+grCiELld/TWVAfY3t5wujBPhMLHMxc6X
bzhmG2qjY7EvkkvSJKzZ9wYkQnDLBVYk60cFU/3K/iPFm02fs8Z4Gk+YZQQBGMNh
JE4aQ0sDxbDMY/waeidTWNeryqVyDT5wuDQs3DAWjiwCiXGntjgD/JB5WE1w8lkh
MejrMW/6n79u26MqlTvbvG+QNidBAqfyS5DtTEcSHLSeRPclbMV/yaQw9DsrQXxK
1PC23d2VBmy7CGBGtj8bAA1OdRORuvTOasUmCM5c2Ww2IrPe90FT0UXdjGOZFKkP
3qriY0e19rvWQJ6CdAz81zsDaWTV1wCgIw0tPz+laLO+IPevyUjM2YTC76FLn7Aa
AJXkDMJyU6BNiCpX/a3GKOcjQIXE2Vr2vlkGZfwz+rVbgHyVZ0K73MNtoWFHdpyD
Szmj9RVcl6gaSQ+DnZG6xFlopFcpRAHPlShNogH7Hl9eMVMzfZOJpotrsOTtt2LT
eEEA5vC8oF3JkKkGIVz9D2QwZCAcfeEf3XJN+bckl83PRBlhaIcb+ZMS394QIwEV
+WFaH1UklBdeVAYDm2L4ijWil0Oum1kJYFHX2LxPAWesW1AF0MTmRCN9Gff4bBub
eYey3BcerfgUTb2P2lBst4UCYpO+VpB3k6Tu1t5BRIfj+f9iwOknux9TLvsIoEvN
yDmpgi0nQkK3aKfxFyvv7W+YRrJyJIayyHepaBGHEuDjeFS5EJC3gpQ4rnnEyCws
VHsWfjIBJNpNbEOryuD/MnPb16wokgt1Z3e+z4FJcms5vJtcnhYY8WS0cdkwXW3r
MMBvIvnNBTjHaiuD7euLDxMNJJGSuWDHAc6lCPYDgW5oJfIYEzRwWV8DFoQs5M7O
hQgS1y5wwkXZYkkWQ1oiL00GMI81f4yxzapJ+LiuOZ2md6DhVJ6wL1jrwdol9Ain
1Pdaqy/bboNfkybv6+lhnKxd/HV0gN/Hgv3lXC7NFS6Y6P8aw4wL0z6CP++E5Lsa
rGK2vQGjNW/RWW1bvsEsxWNtrKsU9Os7TxkZMsfEjQMCRDXucxAY+uyqxCVnnDRD
zdv8qPBVZCCkLam7UAOLKdZk+fEvh1Nf/AeBSs0GM6IvTabHCKCLZV+gtx13NQZ/
5HYLZhr8xIazRYZL64bVp/bepny9/IKrCzB0xwKmnz1VQKR2S30104P0L5fOWWVl
9a/71762NLsW39uqEJvykdvk+l1Oww5Fx2GARfZmFCGfwIuoa8GW8hHg/MQBsVJd
MYGN7VwYjN9d9Zanb4DEJQDVDtTh55q/UQvOsY0MCYR3XtbrN0MsehPkEgGZq8YX
l87t6hFbeRh0Oxvz7sH2LMnpXn1BIZONNvjudded2edIISccGpdDociuV3fslUx9
r1kbd02vpfvPm0DBORFV8H4zc+xo3ctS4+EvSZlFqbM7P0mxACmBlL0igTz/orWI
B9/G3KYAMj+ICuk1KNk7T+Zj2l8xfODEC24bRVky/2mOuMzSiKMIYgF52notaA07
cox09HYW5127QCz9aPMNH8F2+qfhUVfkRFdFkj/Y6LQOv5uRqroM+iJR5AN6vRtZ
9KfdhKUlDCx1xZjrzqjLvs4Sv855rAXQN25oslPwHoi8yOlyLjsuP0U1TvLlxcFW
4KQOs6sH84x6lfvY7ysY0MtXOMYjPAFxj0XXol4PJoDYK9aUEdacXmQ1s/6g41kv
jDm/Cmnos0IADX3qXqFy/xpij40JImSPsgfPU3aFNX7JQN69M108RyK6gFscXJch
2rDeSPUQKixRitq7ZUo6veNsHlkgNlms/CPyq2me8fkUKGad4AVMi+wP3YXNwWYC
CDEkHxrv4NUmEAoZGmAlkBZ9P7j7S5qNVY+lv5Hm2T6EMqR7NKMBP4y86x/4RpeT
t67UhdcfN8NMTNs5afBTGDsESIvZFpNA32bsL3GzCsfDcuDABZb8v+/BeCSGxATV
l9Jnaz836ubrQJxmReBGHYYfbWk2XfznPij4tk7BLohGq2zgpPalO7Uxez2C4sG0
qpzmRyx4qHmeSEF21KNJHdck3aelEb0qGFKAYDmYXGmAimep+3Th2yf3tmkHTFBY
Peekur2nliAvuyiEsxxYrtbh5fquoZCQuGmgq3/FCXl98Z8+vwThOodlj9IxfVr3
ZpC8GIbS+w7JgAkxaOkCpTUggR2xYy/eJ2TvYbMVWYv4MrVTp0YdDE4l9ELCWdCC
n/QUYwEvoLM/R/YZ9k2FlDcgqu7LxlvKTtBAXJuyYq7DoWqBZis4vZU+vxKx+t0d
iLAZaw0kGeOaBD592eSXrpaswut8mbM634qLaiSMnAvL3mXqKGvxRdbaFd+Oi4HD
D+iz4oAMRwauteFZJN9CiYvwfI/fZjAqyfmkhZo/j+RvLkw5AY0WImE1d/8Z0dmk
m/2+E9fwGcvwXoKoS5uVfVQY3cyFgkXkybeD5YVK2gtHNgShMRvAbFYne+7PsCy/
8pOZi899pRLRS5616mh2NRJa8zbfzA4ZpYK7B+iIGWAOnpqAmx+3FT5tOTbKr561
SgjcSFvfCqleBuug4PgSjsdzxEP7elOhlKn5jG20r+8MrorBJTh6tsaHtbydeWDO
R1MBdaHWCh9e1h8SC+TSugIi5WKdq9UP8fJQyar20xcZGtsz1OJ2aUBD8SM1sn6+
ctA5GO59CEfVxB9Nv54oR2ZjSIGv0dHCJ8OBrjiSALPRMFYxE6wiN8VbI3ykt/yB
KymPwc3bXZvjpuNOQSp2jJZYIOjnOp+ReC7e33Ok4qiit8LzRiCrMnWw4siU76Z+
G/dZvB5u76gyvrsb6B850SvDS77jxJ72wPFoQz5u8Gc/RzJ4F+DFYfC58KgNYIDY
2BptZAFuroG0Ek/F8ZasvzsbuqFPm9hFmBRC56Tusf7E02ufex3GVgEoM24QuYzq
m3qzi+B79scB8QQ2BAc6s41qYtjl/bj6cL1CR0aUAbTT0iBDITRXe8dKxAtSBDks
QJJhUoK5oBCz0I8nHzOqmBmURKwtKgJGeiGb7+PYikp+VHLT47dwroRQbqAe9v/5
aJm6WXW64IdfkVW6fRKbbfqSF6bVkAilq8ApiKOIdS1AWIRxpgK5fL0cu01QaPub
Di7YWun422JvxH6oWVQR8Vmq/nPNklNitKxssHazUnqovK2IUwUJzDY8KioTtc3W
kD3xXKrHxQg62szX3u/iTO4N8yYwALe4D3y+q+zVdLxmQKc2fCS/khq51gkt3QvJ
7oA38Whoc0i59/EQ+7Ei5mLLy4IRqqVqr7jDDqn0aQ9RmKbRgtNbIMDTiR0rqLtv
XiUuDpenkBOIEg92qXq4xEO4TuobRw0tlf5pe7aB7tp4RB4a/k19i/6gFTtgYooW
NtFt4Ocz4n+3OnG+mUgaE3/Vm1U5ajZLnWvztoArQVRyt+97tNnaRfeL8EPJ3QLk
Ob15+FMi6xJhYKmy7MLzI//XEgMklsVXbyLl0JXjxVkVgtvDJUivYszWUZRzh+gN
CYQWnEzEjXc6Dk11aP5dTna2YKITN75qTZ7PGm/KYadtMF9AqGWluqFxcdvMmsZ4
P9gMgpQxgKp4CiMExholyRrkxMUd6Fxyh8ipAyL9VSR4ujgwTtATMNNvw2/5CjR1
qMZO64nY/4Hn7AV7hUqK6UZ0QtzkHKG2r5WfuwnhrD9C1J4rfRFhHa44+2InUbHx
Rx+0Ws0XHKgoZpPAy93nOofjnUoF4J1VIZs3fEFQklwaXgi0/6Xz0vGXMgAbXKDZ
nii3ThZlWcMQpy8p8icHClWepB9JV0+o/6KKqY/fiQQnMyMFTAkUU/CxVvOb6hgm
h+aMjuCKc5d0lYEpnJHp2kD39B0GBDH6Ffy4d8Yei7HhQMuu2tXX0JPHBqCNlAAa
zf+g/qe3y/+ZNP2YsHCsHRs4jTIsfEybfjOzo1EA9Kp9kdEiFsH/VSAQ46YGTOh4
Nh+MjQu1aGxwNgPyWsak4ma44HwqYhwrACbhLl5zJ1XBXOfoy5fuFeOFBWoQiaLN
CQnJaQ73Yu4My/9cFgPfyiC4EsiG9gFC1JHY3GiXig8gRGoMa5itduNZmIUSZieY
3kEruli85VmFfPrbwQua0Bnrz7eCwm+BOcjhhBhMJt8CkiIHDJelZj6Mn69K25RW
JWhRVeU2vJ8/F5BSxA4W9Izc6+p83RuAFXozPV/5eRClDmJmqZS/JMYVs+Xko2IB
hfYw1GMZDTQ3s+A67SbpSC67EDXp92Q3QIxZrB32a0hrpzBh/D0776GQ6vf0h9Bh
0KWjTnMxpmNmNpu0ILobTlJBYMZiBezk/0A2mWOlCZ2OQ9vokwKxDonhClqgp/32
atq/0HJRrOxwGgbCOxoPIPfcz03HebW2VgvuThKWTH5APJvFqt1nrX+qg39KKF0U
LXZcldslaRevbSyDwx78pPHmb+vGL48EYyp5YgOg/Rr1pl4qU3zh4IC1e5aL+lqu
d08eDIMyZlH7+fp91YHgQ6KWhu1MsnJIbXMEi+lTv51EfdknMFnYHTFOEKwGYaQm
t9ACUZ+FjTTKUX85ZsxTX2mkMBNfvWI13oEtNlg7iZUADsKUAsbY5tQhUgxiiqgM
cZ3tE8SqrDp7Tjp3T4cwDOO4sqTL1vTY6F5sfveePAg0ABGOhPFEumnM6ZMwmKG6
YIgvrNPI/eKmjoYimva7aFR4Wr17AZ7ICuVgyWGRyd3noDLv0ua4bREEEd9RmGgU
THzI0ED6mFXHAyaPYxGgih3HWpxqy8Z/IrezQM3PvIw27378CW1sCdC5mn/2WIS/
hIngKJOt6x3eD69JOxPZ6FL3IC02HbtFD/q9t3DWzla6Fo/LTQt8/6AvRbzsUM5u
auOoho4u7Qksl7uvUrUvl/BfOeAnS/bMcjB5bVFRzb6FRRTD/Pj7lTmE39OAcvjt
nsshgAB0ytyUaLcEQT1rCmfRWDM7EkoxSL+D0oc7ja2ZZFmxqG/76q1vYCgzrufO
J7XYRB4GRJlIintmbDhLrREHRkHr5iZXXEt12R/Sm+GEUj17IzQqV1twWxO0d9C2
2VPjPkTpDjZLMmDd8M5L/liYYBhPxykQVB3bWJxEBVUMjt4/CfUNjZuusXkOeRSr
pjxMFhJNotZwyb+ysH2zzOX8TwCsVJC3xl7HWsdy+VeyW+lCfoSF0gj/RkG2jeSs
jg0de1VF8tSEbMeNNvOm8NNhTAZO6bkGqq2mP+4jtG1Ry6tKqHcJs6UMcI9nWz/Y
fBUBJXTWbj3kxhXmnFw9BaX9dX0i9OK/TmJfIWtRdCvjdNQos5/Pd/7CfV4klabo
Mmnb4tH6SzA4qnaTQdSYmXc+49bMdb97D3+fzzhriYYjY77EjoDx7LGOjj35Ncax
h3xEU5QbhsKcpxS2z0R4CYHy//ziTH6p6JvJ6iF9ZQkLuBG58IJy47HE+Mw0fRmU
w4yXz5y+Boh+t0iDGkrq2jNDob5mPL9vdW3Dtn+8Ic0Q9hfIVuGS+bs1jROXGxCj
+OtGbRQzICCA0h//KU9S4OQudWyzDT/7gofn6YFQOd/avgKFAX6apN+5QnFZ40y9
u0ZlEhrQh0EtuBffjBibXGcGi/rTakJ34HAxE1j/i8UPSgKwZdo5VFLaOMLW0u40
iyjypuunxA+W4PU5GAtLfqiMr3A//wfb4++OBhT7WVkcPEXVJqaAC4sHTbMnfNpc
BYUtjG0S6jkWFrrRiXKiWrnzX/C7VtsSgiPAmGFZVr7wfm9jK5sAlHVLRsblLn5x
fJ5G9eKjo8jaI7eBP1PANpGDIfwPYH5oYqX6gmYbx6cYxDfhOysh41nS4qU60+MY
YENyNV1sAHhk16Iu60UfAyUyhSUTS4mPgwaVHbWTILXJGeyufQTE/oZotk1z125p
+CX4XqkYqOjFftmj08DxuyvHVM2ZTrItrkUbTsGos29lRrF4Yd4gwMbwtteOpLze
k1J6EgMGNh6tVq4VQeSrJQZf8k4vco4GNQt0epRpBtrLyzkRR1nl2/5RiNfLv3nl
tcFItOkDs+fxiwthJl9DHXrB1XmvHfFXRHSFTO+1yY0DMGRiqsAq62IFt29vl/bm
9c9QjnJg//B2np7MDf21/pfKIND1RairiX5UhRHM1gKc3IcFMxOBCq42hK+iv8Bd
bowKzuxjTpYqsWAgWA1aF5R/DL6CesqxEkBqugLp9vEVYaA0XFGQYEO/i2+IFodG
y/8zW/dcdwg3bGh1q6WSBWmNFDoB+2wj1d7WZ6zVFCL557ttzLMZ92uhwDWkEjRs
G21UhnPt46+uhuMs/onrENvm2NdHJaG/NtuaPBoGB07/aSYTiYtNIV/t9hNdbRNK
Kl5BUWt6Qh93cvkN9BgJwSxT8AGXVvPWaExJ9DM4d/hEMrX1FmvI3odpaq6knx+7
0EtZ2khURzdh/d5PmcVUs9q81qK14Uv4Y5JkFldHfdrK3RiPqpqiu+iLszPW2Qjo
hkb/TejMNA+vb6Myab1B3O7aDCPjLk5W/UIJyg0zv/izd7jzC0TFp9oK3NUkwFH9
2ZXl8mdg84N9CeDah/b9AuR262tpGg9cQxE4dspD+Qvp9rxM8JS3KYg3o334l8d5
JjEZ561ffnteALq00y8uLUiDkQdsMpRQ504/VuyK529M9HZgA140/IKjz7zjHkne
qC7VAxi5DU/VKaTG2FfZI59JOyJowz93e35eVPwVUfQNoRfaC+8DhKGxgeBmnUxO
5ZMyJMBEMPuOrKAv/81exMz5LM/+pHgsk4EUP/3nUeTYY+4+mbYavxP3MFwR5XAG
nvRvAsJQF7lDDvsSPYJqgpSifPna2weferM/3EpeEWsGDwKJSwqNn8kO1si0NDzR
+IOc9iwczh8x2xDDHPpp+ochR5hbhG3IPqIxZ7Bg/ia+606NplO6HBJ65Z8A4iWs
RA/vYQ/PZUso3leLuue6FmEeMPAOnvlI64/rcPjmKmH4LR8w++oRcXjFMf6iw7s9
zbtLDgckdzPLvw4xfiizJVJQfqChC4dUc6d8AhTbqaIw6g5X1oMVMDK1PNqBdwgS
PfMnY2UyqZCEaC6pZEIJUW/U7f93pxkBZsaUvCI1j9F0ta5r5g9A8v1bEEB9Ha2K
IGng5vN37CSMeSFkRQX9CaV8qz8jsFGNWqkDJ1lbH5rNoOlemvLrQ62tpq5W+NXm
dRNhTu287u8/8TQ4dnC/TgbSQRVElIl0m+p6bWwY9Ci9pD+qp9phXc0PFDZBx4tV
GdaPqqVx8YHVi1YTZ+cKnXG28k7ZzPoALjurGx7pOcSdBTNgJ8U9mdkFOpQ0MQbg
8+Q6rLclft5GJqmdPNUzoea1eUpnkWEek+oXVzmyVALmQPHu2F7Ie109zWGt5cmA
ubekmew0hRed1TbLiiyGh2eSdf7t2NRUM4DAOs3c9wOaJWZsoVPA06+5EvsAVzVJ
dsDx1T4VuMur9fQsS8WWPGMPhzt46c0KFNggffbtOJ6mYF0AW2VuMdnsuH44UhA7
LiEcGbMQzLDvInd14beZXJeACP0ThLwlRsEKuLvuAEVOO3qvbDmkFKKZVxS5xTQH
wx+CMrh3flfDtRSTSP49KOVZFIVJ5h9sgZGZixQqzBBohriVDTiJLvK2yqPjX6nD
QDZQnaTyPLKE9/7n55rmFqUX11Q+388AMPn5qeeFcAsUSToZoAprez7qQjy5iGk2
uYWyDC6fRWgPJMAU5r1tZaNbOgkSZ9j0+/KXI6FPQRc=
`protect end_protected