`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 6592 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/9huKRhRMtvnNqb3Z+UU7TahEoHV+T8U3P3ufru7l1O
3DlgtZzb9QxCbOjthp9+wDkjygH0eUfDrEl1ovhZG60YTjH273PSjMhddiNs2jf+
fHQ4YLElvb8w21FYc33B+0jFtcaRia4XV9OreHrqfkvQhCfo0Qt200RYM0W0ZtRU
AW3W03IvET+34l9b6zwVCevdD/BIGlZiFub+t1c9L63EvG/Y7w+zKVnoNzLSAh//
n+WJmW4HVLCoBnQplLkWMYNfHvBHoy8mZBtadOVJksbEcs+MBK2nDvGa82WqKZIQ
rI4SdDSx/i4Xq4aS4mXntoTMpYQHPuWqnDSAD5QNZ99M+ylGzT4w7AAyx7MFr4e5
IynAuP+4ki36TlqgM4iPeLdkRAT7Cc12LhJcfCgNbIVcZ6tT2DkMD8w5lBqop9Cf
urcNVUbI4b1yFxxCgUdPqKOnDCJnexU3YdymqTrP/YS46YbOpEE/JN3fb6eY1/DC
4seumWBVB0e+MRGjQ4Pr/p/DBF1XECZrO4qQE7ovFmAAwPknALSe0eMuWhhBL5Rc
dsMqGSf6iWNmY/8UrtQxRFwR5fYEkeij3xjUeFAs+Zw2mso6esH4ltQfzCzBAFfY
4WXcOqagqolBKYRgPTsV4UF8wBSt2CNjDpRRNi37dZtNRWbtFADvIRAFpWFnos+n
r3Jv7YuFTJuaK2QYD4ETWvfNBIzrQaVXJQS5BLlTKSQdRf7ZiE3zpU/9HQtesE3H
QNFsVr7/x6OZZqBz5qui5/0HCNqK0Zo60CYSMM48sbhHJwiG/MNochIdvN49Njty
vqdl+cdII0GT8eh+DqylX/H3CH9XfQN4W6yBJjIWQ8sNlXNcB8XNkUGThe5BvelN
E4WCRKOHKprNd7+Ac2L5AB44SP5o8zWdEVihN6UVo4/jbtj/iFHX+j9aif9GXNLs
Rqlo4sQVfT7tpJf+E7G8ORHi+X2IlJ8Jyia+NZLbRsAiVHmD6E4BYdDsbMvlYd1k
OoV4CzLnd3u7kMZslDNy1hcwqvm8WsppeneHAUYShb93klYgCQAPJQfOG5HtEX4d
Wu7dBIlAvh+37nlm7eLiaPJz0jx/Nf8aSpNT5q+wgzUwkCQ43sdoK796ZOn7Ortm
gL3+kh3vjR5iSY8q8eeverkUQ3kH9fRLwHOA9ytDVhovk8GROJsq0LrfzKT9+S/T
qKLBxSbja046L0RDbQGWxXPNF0P8US7AsR6t1ko2BP9avcPS16ouwobloa+yFS1D
p/j4Yeo5y5dlaKmqkZabHPKsVzezeWXWdBoPQ3/XBNwOzGr/D8gIVwmcJbylvJYv
LLY22vOjqQFQ5kgw+Sr2BmTiFFOh4nJghgvYHz40crF38PT0ucd5omK3AAmczmU7
6gFo8RXFLTK49dMLg9qcZ1xBlqXqTf38tM38Obashjgtn21CwKBtc9IKgLb1SuNf
hJ8WHXxBRBdI4Qb9MtmkI+tLrI0l8JSN7/lBCDFG/fyPO7AFcD7tykwMdmpUUxOC
NMsQbkGTmga7XQGRwi5qOSFbrNVRyZIFk1JxBMs4vtY60rW6mmEmXzXlGWxeVBjq
NyFg/PxfLL+BZj5rApDf69lez9sAkhS6+UHYDcHOyTNZCOwjDB2SuVGOsKGcSQjY
HOF+pQjA9iin/dKeIH25P2O26lSPKndeC+xg9IYOHnNhq+6Cc9JlcqMgWZt6wV3E
fg2hOTlhndUJLy6eAYDLjfs9JYX6gfbWLDjkzpG3AD6ncW/3amnugSc4h8RbFlVU
0NBbTdhc6Py3V+Ndv4zsNIbvYSfITrg6Yb98SJac6MTphY/CaDCoDqRdNx2fekx5
S1dFTpgI+NwLXA5XYoP8VSL5LnW9F6UqIiiiJLdKxg1qfZEHkG3lLJaZWRrHdP3s
HsFKpdkgmkuiP6VyWv5Ak8QocyTNmd1ZTbdVXPrZcArugTXwXXeNWUHHRs+5uo9d
h3fnon+Vz43TWkCFWTmj7YxuumPgbBrStR4sZ1jFrVAsWu9YM0GUqkCt/ioBC8a2
iI0oNjesarKR1kwx9G1sL4m8W99nt/TsIvkTOkyUZluAZRk2y3VPVD52GU8GRnfl
j6QthMk7ivjZTtz6i2d4O2ctWl6KurzrcoYaCcsnb43kcjDld1xof/XpJzcbsz9U
Vc2gJj5j+SdqxGOvKLKXBkyXQE1kAtgqimusvnKHpePzT5KiVmW4iYFmVOF4yVRP
woi+WUnCoAD93zHAuKOCwh0Pu14VRA8IDUnBFqEq+uEsmUSGZQvlwFEDNIwvR3HV
eRsw4q97cA7lqXo7QvXZBPE9c0Lj9nyiKgupzc2M85n6jhaPWPiCkKxBXJoaBxPe
++CBisV2/zLkKXgSEWSnztUrBwWfwizoMaYWF7PqnABktJrXZ2RyE2FD8Rjk33+e
jX5ceGtLu626TsOr2zJfUWrOPT2m5a6kiOpH9E3zyCGUSfnkQwKqXEbBgd39tfOE
LWpb1eIlOxf/+z+6bax62R+uVTrT0c4kBRwHUwgxMLUR6Q9DwgRKeT25WDXTnIey
fzw+8LBt98ExEXIAr7jHgBwOk5wp2Fv8S6lW0BK9QHPrKjN+TNH2JkaDEfBBgPtM
HHGMn4BSAdp23m0tWHf9Bb8DXwT5WPEXXJoetmPgbCeGBHtzcFQUrKoEasjotDYt
2flUXNjDCmT8m4zvFwOn9zpKfFdPws+16F1cfx2RpXTHkki6BEtK/SMWKgsPDNOI
CjSa5HM6LGqyynRZuwFCHtcvQmdHZFHp3teNWp4FWOzzpBip9YqSuy9k0hD9yJ10
JYwrhDxcO+9B9Z3Z4s0hdyV5LVBuwBTkZF2jTg+2lhrzZDMW1VEAREUK9WPzpdoh
i18vwACCbgGKZV5B3quRyp3d5lfaNwRQaZ7WmZpNZalH82EygjdkAl8C3izALxAc
UBACoyindv2zRCZSn5jEu/H2Ag+FbgiftRwpB2P1n/jPyU0guXj7aq404jS+KsaL
euQXQT41rfHXzugH2aopqXTuKmzootrYKOBEJzFAJ2OZGYb5de9ipP8/5rIvMl6S
xM9EFCyQQ2dH113QNGhCtXegNLrBttgrzAamsXKrfqyPAdAROCA3VL6PQmieHwt9
s/vttlpn7rZh49Z2XKHE0v6twUYtDaY4y4kSvjvlLnY5bjPJ5hQXadS5s0ePe9mA
rlNsKEXDAl9p5JIFshFycgTo9Uctqr3Ko8cEScl21XMks3PWwV68y1BIp3/+sXdV
XJa6hDGMcgaUh0jTJyUwcRQ/6H8DmJzGOn0VF7HNQtHxpT9zq7v+a0jBMasrqTmK
WOlLkaUzmfvtiM5dvk7gRBUV05NiRKgrWIXZJ8vWguxwk1XLns398YCqwUFLWwz4
Hh2dY/JIHuFyKGv7WNvYJ2fa76U5eVcb9D3e/2621dnII+vXQOkWDIW8fxpjdWq9
1Zm3gtqmiMOh98dd1/RkY5/9jlM4KS9N+3UBMnHKrQo+E9SZsvKJyvwhZXHWoVEf
HLZMacK/675NjhBtNiG7swHnTpgqbTSO19dHiyWcLtn1BLmA8JCNT4tvsqvPu7j/
6zd2c8jT/XH+ipWlVmrIXJOOR8I44obBODwfdJ3c0dP0xn2+c18m3MFNADTOhSkp
vPN0tkGvsEqJM/DHn21tldbasWjC7vp+g9Z2oCEjHlzFfA/AsaSBWWdQc0HVVIcI
68NkyVQqesRPmi0zB9dg9Kr1SuXCjBzHSzERhEvemSJ6kPQObvPBaP8Kp+hvTG7d
H6Ewvzndus5lFYiZD2o29zRVUVTc4MEEo2aHOD0PppJq84yUgxR+Y1rsLVqFvfoE
Ma3L9hDIMqYuGCacH/h2+iDVOTJnI9ZLC1OVeTgoWVc/wi2btxjjTZaRXYX3f4X3
z3yYRQsnztMTmHEWRsbej+4wL9aYxf1XMy+1r0pZKeMCFGZep2VuJrIEn/QomXKb
+Zmtdv05b+xkcOiWCS30Jp2/u/3mknjfDF/nZ1qsmGyPHgkUCSexWfTRW8SrdT8R
dkFBHJnDA1iBuweLKK+uqPbeBIu/GygnPiZt1uwhpGXDt6beZyQrM5HjhW2F4dMr
CNjzzS7853RIZlcKpfyywObXgiAj8izAWpvlMSHmGKGUQxfKpds2BnQocFbyN4rI
F1eh3Z0YjGzXxlE7NWMbbJWGAmGvRMCZtI4r+DADWsDhTISgA+wKuRAuAXI7QP63
BTDJTAXmpw6jkFy7TJ9OJfZ/hYsjtcteQm1RLnAf6ZLpXc7JJokH4XbvThdB99/f
tgmce2y9VdEn2j123vOXcIkZ/jVvueYaie7GtKtqjlyCUps6wUwPcwT2eCSg19wA
tGDRde1R4VDXtM1opWMwLfBI8he4auBZCVvGIp46g9odvxon8ZOnTgwJYOqj6Dmy
7lq23ZWLDiX4FW1bUHPbrtwx59hjuNdgT2jPNoIAnxmpHh3oxQytd4v5K8RuxNJa
ZMD0qMbEAmuaz2weaeFC9n+VYtfpB52DKK5tZcITWC1l5uKdnyAGEPK3+SX/kcnr
7tg0SUF4WYDga3bt6S3Ux3G12EU62SNB/2p0Y9lFlIP+H8mA7FSV5tLV/Y8faP8j
Tc+xEviH7PDeJKXzCAA40P2xFIqGbdBPG6eT5U0HMmP40p/5U930APSfBtU6yrAb
9bjCq/laupGoKQs6Tqgrj/1S/ZpjlpIgn5ekWgODtEqR43qMVAkEwb6lWSXmYDRJ
V5zAypfnPHPEtG93DU1PSnk7QmVDBWouAdmPhydbP+qS4Sfl/hS6WkT0fUnCmWq8
clwPHUntzouWlHwbFF3vbvRwoHdEtkYI2Sux/9uJ7nfAKGq2wkR99CTbqs8Gaetl
PQmPpa6hZPfecDVVubhE4NoIqSF3m643JH5kJHCnw02vHVgwOQvCq8yXrK/Mc1zp
2aUY4wafVf7r3MvUeFfm48SRhEk/KPAb8b+7t+r6MyqqmdgCwd2Ui6mu7vaLsZh5
OSblDYOP0joZEMoVDtsuwVzpeq6DhQapIQMT+tn+molaMlEJIrVwvFwebzSFcPgJ
pmtDftVg/2Y+tabyioUK3UjdSK4ztgbSaCe1HJiJla9+0uX5YRtdHaPxX/XMQSIy
GYqUB2K068ueDaKDJrY44QiGUEYzwtSNd5UG/6+uoBrJrAcWNRmBowrtH/D03S/o
8ayNS+A7/4yAeT5PTCe/AFFfFjKF0a+qeU9HndDD6z0kDeLVeFtWSpCebF1y4x3y
3ilaaBDPp8Vux5vFzRKWt3ec2gqgugRf6eQVi36FMki0LpUKLqpxD7gFRQHdFETI
A++OvFEvJCAqg6ThdoylAp6AdBnUOnjHPBCqc3V5/6hWwA0Ys89oDGEfmizbXN6J
tXwrYe3ctnPkWnG6Lc484ENjEABJsN+1RPclEzOiEjxkXZj3cdcrvEdxTF7GFOMO
55MJSKnv0v/dPazcRbuz7CeD0lFH9dVGSshjvAlCTmrKk/zIEbxphDXElwyjEfwW
hu48/9fybZ8P5qaStvSb/Png2yB/lrDe8tg+/DM1dV3+f46+7c/4ZTQMm8fdDrxh
W7HhDohuigfbX3zcOrQWPcH0ORuJJi4NFbeWLDtaqJ4D85n8eR276Pcm0Wf1exyr
rXCrm4G2bfHI6Q8xwdQHoIRHDhgE/zZUgqsTwf9KmMPdM1r9Jx3HtP48qdKN0c8q
QA3YZ2qS059yOrNX05Shij1bkrs+WfJ4mP7HvXdw3G7FHDtYUzRQ+lbNKf409Nup
ybXu3VDW8appyjnJ6n6gexnej9hsFjC5ZU0eeiZrwI3Vbf1txKLd0SF26GRQJbQw
h4Syve+QTHaPZPeAyiMo64VYvq+aLAF6oZcsrsBV0UTXEBcBUXKAMVza4EuMfmOb
Nq0n5TEnOf4tvZA/CazTQd2VjNv++CBKYYPvamJcWEEJpAA1L2TDG/2Gif/htLnO
5ESbIiYC1JeXTTzUc96wWieGX/NLyrh/tI7RMqHv7eQPLmGCbjlTZadTe7Mh49CT
TyvbcFtaaTFCKcOomf5Sg2T8ka6nmlIq/pBouYCbKC0Bb4nP0yQ8puJgpzXcWraw
yHRMpZ+/zOpE+etuqDpirE53I/AN4K1ex7wV2svp3JqJPqz+VzuZ9m5puBDFIRT+
eISh/HR23mNzliwqEPHOFllWQkdz3EdBPavWgQVT7p1d+Pdi3KOXE3/RKUciHWp7
iYG19LUZbtD6AcwiceDVU7p8QCEZcLZFpZyFJacOJk4srlfYA+5KlqqtQP7BYN2Y
3VXG5TtBfeRp0c+4a14MFYH0MI8JjLGJpG8tiqTfvvbWzFRQ4xoe7N+wWAJ6WScD
W2VmTD6tuOIXA0vqJWTemK0JhoPAK4iRfsWiFvI/o2zUOfi60V2pU0g0gw9JALrB
eEWtUsEMCl1TWbnU+2Y9wTTzoyC7SshZ8i5jg6UTJEAePYTdugkJSZjsswbBS4sZ
da2IbJza8NEqURsjLDsV+Ly3rxyUpfkHgr4psS4hNB9sCj+OVIX4eg6mfqZnF3yM
yizarKc3xL7in//dRkqwMmPCxftv5Jp0RXNxGUMDv8M/1WdZ1tPAqD/l3KRE3jeQ
P+3CRjb0F8PUHnlbSWMmxCdhbhzB+ckrWPNvU4M2XRQC1Gf/dbgCjYKuG1DFSRyx
r+2aVqLi1qjjFNIUNIsbMsaArIaqfXfCTZt52k6k/crEBNUpHQ33O4zyLgD1Tc1J
UDnw38QMn6qJpJBWiENxzonuEL3xEySbTpCSuhSG4yKvXbIYvZYDXW8t+7v8qXe9
ZKNw7AtHTVcg2SbMbmaaJu+T4Mi2ZbKr6kCLsAgQbCtakNTh76UF6TSmm+httY0K
5XyAFozyrS5lXuTMLfF1s8/hvt7cJbCIMGlxea6XGlwrwWYFYg4JdgYsThIs7hr3
uGOLo4XmefoK6BB1fS0YW/sB2Jd4/EB2Y0SCAx9wOwtOOiGSezqfrkVLNvrntjAf
029Q41+Xr6TR1zccjZahP6kxBwMOwtqAxZJfGq3zHXZuFB/1YzLqcqxS7XZpPZUX
JS69VRtKMyk6NvPy3JQ+81jHRt6pO52mR+sxEJWv9aGMAjSl9sjByNhzv0yG+32M
PPHWTQSFAvx848CdmSjLwT/gZVsYiKTcyGmQfpctbJVqSfbhgKSWXmpG1nSYTXbn
o35eln2pnXTrhRJPfnj1nFMBkn0dwu364WBDmvKoX+fYWsShJobo9E9kDNg4tTsi
u2u+SQHTMNy0HjQWVZs6vgVqr58bcrCTX/AEGHQLh16//cJNhVCSxjHEISfrLYZn
LGgVlreoluiCmIjFlSyjWaV8KUcsfgImX14eHdINaj1T+r31KcQM14J2Bs+bCDH7
nWhM2MiQzDuzSlPeCQcHtzpVt86Modyi1+4IsWGFZ0pmArKyNJ6/oziXqMxaDJAz
JMQ3yrcp6A6g6owDbHICUATedu2g8nZvUJIE/z68VQHTIM724yrZVuwFW0m136i7
tXi9Rex4oQxdhdC+Lax+i5Y0Xoxk2xwKB2XHyZpyLdbJ6UxJiGwlpgKiugYHSwLD
QkpKS6bMYH7P1cjsx1Yw5ajXqNPSJFA0yP1yVrSTfFYJyXgVwybNhoc+fU+iXhmi
fgkTqglbAi7HGfjreFFaXZDjDFXK/w+k9MznQaco9e0wpIzJDtCb/Y4bLrEeRx22
niZohHEhTx/cM/SKa8xzbyEjFwCbpmFVbkgRJSIFwojanzFoyr03DBfBuUWB2T7j
2oyJN/8dy2P8qDEl0bNVVznDG7LjLezxZ4CUgFDlHphkCWn5JvjBgpKgZiE7TeUT
xWYZy+X/TqszIjQOlmCy8KYGA9Y29ezNrxXYOBKqTf+ihKgFMMvrkwSTm/x++uMF
PGaOMSy6dEXHRDXiYmQEc2PeI5ZDwMkJnPIj2CwLAeDzX48ltltl9QMXXd3BzoiB
m21Rl+2g1kEMUZVqcSY+NBD6I3OMTRqdyX9CqeZUhheYirmsYXhWg6sA/Wy4pm3M
b/GewolnBhiKx+iYpiCIhgMJkqy1k1lB58ycYTOkxI6lMLEN/U9xp/Ii28LjZJFl
yMNOLHfbeqKAiaHUboGI1OsfmopEGAHSsLXaCA10PA/OPSVxcHmdSPU+d+xG3tZG
ik5SNgnuOj1wJB2Xist3ARO9rt8uE4d2/ZvHY4AsgLq2OvhTF2O4N60bP9LIeqAh
wYj5VBqXGOJeqbwvdX5NOp4tDz/4yRx8GkeyV00/jskAeA50yAzc0UeL2qEKEXrs
PRaTdrnhpkd13/zveEQb2w36GypHO/nbCM6Hj68TRVtIDoQ0av23zkG3oKnLuhys
PMVktZIpd19d9gYWTLDjjxoeozLUp3Bm0P3sV9xGfu9ZD0F8otgzn480dQgvqNGV
V8gPtDNHxWEHcKIihOyVsEP/jTQv9AvusXWmJ5Z48Ara72pl+P0GMwvb9qGd+DXK
KbhbTbUzJUhT2V8iy2KJE4uS/vK8n6+1oVHhJsDB3x4woi8LqtrqWsTIjfEuL+Kc
MkWYxdVs5u1KEto2hrla0AbCGPLSMjW0wrtmyGLMFkrT91pKEtqKUSmYuNUSBxNX
yHWmS5dPau+rFq/UCPNK0PNC9Gl2tCboticyn7Pgw8FdVYfPTLR4bjYtWfCHOJ4q
u4cUZO9XJSQLicVHNQUvSqiRhhJPqHh+zhvcAxT1N+r7xxHcM/dB2R3cKzZjPxoO
cZaQuYk7BhgJ7RO+FJzL7fmVbio0tu8oI66lF9aVZHU24LcKZlVdWTgc9NKziTlE
I67CKiBJaHbMd63w5xOHmw==
`protect end_protected