`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 14624 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/9huKRhRMtvnNqb3Z+UU7TahEoHV+T8U3P3ufru7l1O
3DlgtZzb9QxCbOjthp9+wDkjygH0eUfDrEl1ovhZG60VzsOe5ctuLjqOhpaijis0
F7eTtOhgZolho/7mHPdTi3QZ90MY33OnWLYtpRXmqYdAgp2Eoy2R9+2FuHd5nvsr
HuEEKSNPs4w1Lig4LQU1Xi1tscW8bXw8S9OGOeEPc/HSQe6hXtsbLZYi+HlEQySx
63HsaPifALLjKMlyojC08Yl05BF3zODL3Ypqkqt9yM+nahh76bIZdwPHmIMacGYx
hq9WJ2ghdSOb2l8EGszLpbWZUuZtREVbqKZHeNnrXvpcGLqW4ed3a4ol/kg2PwJR
/X7I10jqjN/SjBoTZVKZvK+G+V/mkUQhxx/SvSRLvQQcRG+zXzu9dH9JJmxo4GI4
xJElscz1NYc/qn9CaUMpufX4UkExO1n0RMWtHgyl/SFj89EQRV3zxXHElowHPqTc
mzWTFYGh3CbY/8p/qugRvmcc7SAMJdBFUAvsq7wYd2czA/Mw9L34NCmx923j+Kaa
yZTEF52X9Etp43+V1DkmMWU7LFVKEAmfvOHodsVyb6cGFHSp2kXxfbHezhX7y7ZP
Fxee/DmCg/uuq1divRBN5SzsPyGBghxGlkDIYuQW7MZjZ+lsCogmzmNJTdhA5TcM
llT9a7yIiLlb2pKPPqv5lBGuBjow99DM2mbcmMLv05Z4KjhIBRxNR0KQoodYvg8p
OjvXEZVZ00KjVNx7acQDr6z5m4/zy/OAsYs/BavLLG+nduUknVRNbwiH6UTaZLbb
idikv8sUpunxl8uKlg2xgClq04bdzb5F3DSMt7Q8CSAz2FG8Ehe4BQzMzuGPOxe3
0eFneibQBKSpMZ6F/fJl43oCgSkQ0H7LyDk+pRIV/ZEr0SGICNQL/Qb5/N4eVQ0H
YZ9YZCafT7ky7Sx7H4vlhbfvZ7a9lsIyhs4VcFjDh3573q/5GW0FbtGCjplmfIQ5
kCrF4cz5s8DoO9KA5OtSJVnPaBpS9eAtCrL1i5EP6FkTpWN4YuZ4MPKNRUhm5+oC
wjOT4Al3z8jTLT9ye7uBGCShgvgIMtChhmQ0prWR3fXvHiTlyhMFzYh2a+jHyqnu
K89An7RbDFL0IhM5BRh97nywKAo6++dOFfMYBxdqMXMXbE6cgx6z1NobvWkuoAJh
zVVfU4+zgGFW1m+eeLmrQ5Y7VUHYBUsgwX0tu7O3E7eCxQ7I0kYA/NhLN6PpOwOI
o9+5hRiHzbpxQltxWDnNDiiEzy8xHHT38mm7itRPgA4Jc1X+917MN7ctXhC1cxWH
gm9p3t9cxxpGMX9+kzOuMayphZjhgY5NmBRe3C62aUXq8RQaCiFDzzRTokoq1eVP
SECAIDWgYzBWg85Vmq88Dw0254uSf0H8yxSfDPlalY6P6pKGNUBluhueqyBGJCF1
nudT+HjQWSX+I/aVJ14lWxBOuIksLrw9MRVOfdXQ9zUyLDIkeCkrIQtHNWc94hgf
g3CgwU8zbV8t7OMW6S5iLPj3wGrAFEBURcKBd/D51XL2Ef/oiTA7ScwfoKlMWbDw
VZ8jOHQaKENArJV1PkLJa8VAyvUC16Oa5D5B+vKNakV2rESPJ4Q8JtgOZ9qYbBSR
EnYjyC/9xmynKWFPVb6Dp/pnNwBVJWOqkqSFKu48CxR7K9VVUkxDM1wfDzrOQnCu
5BUZAn11/ByijbjBSWe3pYDiNdPLFw28gyzrIwxrZG3tqW8Jf0N+Qet9HCZAWpCM
XhgxGOiTo2H4vmDyuKafmQzOQtYn040ztEFY/RAf91KHr7EhVYTYJe1sx6Gkr8re
yfdjPRVJ73jUt79BeHlcuVlxsYWryqvIuCvbxHVEC0Kc6e8cGq5v8CqzB1unw/Vl
IwMt+hRCj03vZv7plikyFr3jgy0dGN7alJpsFI6RzhqA84nluC0Oxzr0NzQVD8Yh
yRe97AXK06ex/IAxtC12v34btm8jiJagVl3i/KQCM2bNAUHN5ifwo/JtBXnczIrt
r62VBRACexFFklRqY/EPkZDEUZgjWSepbV/pyCyufUloKKhvwrtUdSxwg7eT6UwV
NtqUKQr4zoakaafrdRVTi2aWm/cTI6OASKSmEJ6t55aTorgZy20SqPWFgYEG6YDS
rxA4uplzXMcWwfF582L1OwIikdPGFqJSAdayGKRwGITGqTtlGx6jQ+UB5H7ripLg
sycBCdO8eU8EziXCg43qkfYUS6sxWqqs59hZGxKWRh29Ym4QLeKE61tOPYCM0eJf
18RUy1iBa5lKLpOJFwDhhRBpSJ3AHQjqH2HX8vWeUJTVpHXu3IftkHsvHm9iwMvZ
8Q92y2tzWJUaw6EMK9Gd4Dw4gmvREfWJGvrXWxizRkMCEJvTtGmQsZUvPGTRrfk+
EMh7pmK0ur0f/vmD8jIWR9FFqchJTxTHcLER5NMLEDLv2VGormPQrICj3PLx+ft3
HRhLX3gRXt6sVBKSO1RLMRhv9vi2ajSfUIQ42FDlu4+waGjc46MR6oRzQ2AYZYWi
HNoEcf+FASy7kxr04vmWRtRTtD/v9WuEbF/cpX/M3VtX7BaSaHAp1pwWclYIxjZs
9RdsGtBHTW6Hjdx2XAEwbKmPpNUPaudYZO+pUCb2UbTG37WhYFmbkD4yLkfTUJrm
QhfCKtzEDrviFHD9VAYLM7o0ajSw6wMW17IWpnPKS81DU1UcHbi0H86L8OowTwfM
454h/2j6lBPMtCCfR8gd5LgXj7C8MszKCnoJfsLG6vNwMImRtY980M0YRRB4hpYV
XutP2Fi2oJid/esRHvj88OJNLtISI0dLZ828KKJsW0teMjywiDytavtKEQX95ZFc
j2edBtSRLxLveeZlgmZRNDH7G6+0teFLbt8xFd5GvPA9Df4Qk3mOmLVEjbF7yaze
rmL25ybyCcGX/rHyBDo4qHquReU6BzRwK6G3av83d/iDkkd2NICne9nD/Rn3cgMx
o6eLKCCpqxO03UGx788ZQ5CaMpPi7zAvqlFLD8nzqmlsIvTiwQ2MQ2WGzr7QUQOq
ZKadKiBS6X5N4gSTDaee/p3CkTatBBSXLu/eXvs8kV11m5kGctLU2WSIKMsUWm97
jTOK64yMV3BNfyeajY6C9RstQHKywwZRMYzT3F8zuSJcERZoX77UD+CgIrsFoK3/
zzoiChdk88+Nkq+raf2ua9iii8Hq00SLVEkaLOE5eAV8B+q0l3UVvirkIQA9LGG2
GG/dT1xKVtO3l1yMsXzk0Qk2tLMmhU1O1+Phjb55fhyH+xUPYT8QXikamFy7Lv7s
Yo1VUTLX+WbyVySvQFCG3HHUGgJP45Mjbysxai1Echh1F+aeq67OGtDD30/96004
Po/eOmI5Uu7tkvcFOsi3yQoFV+boa44ERG3ALiuw5YAdvUsnJlZqyylwuJkRlM1i
unz31WsQjMJpX3A2FGEoPpnWvvqy88c7K6haw4T2f3F5pJtf2qYwRiI6Dyl3WiMp
toH/7PDyMPwnHj6bqKP0vhX39GGkOaHibpNvSDw8JT3vZXcymKBKNoy7oFKzAqRi
w/TfVI1kZ5ytW8gXj7zYFht2fgpwHdLIZHAOpGUL7zr+e/1w4hs0rQ2GhxVwVd9y
8aDSGOkRppjUaC5yfgfAFAP0FTj4seCtHbQELwd1rxtqujj+v8Mk6Xk44LPQdcJe
Yxh1xIiN+NvTd7JlJNKuPqeOepYB1dxnMD8k+zZDEfKtOXKshRzpYjGEnHqYjimF
bWeRvfvfd6eXjYqXSMxmra80p28BbR/DJrzKnE/Hm0ymozMMr4vOqH4It030LfS2
mCvNBx1jxhV23ZHW/av5MeNWW8NtsfOUHCbdJ8Zt8IFaEQ2Gl86BBDWkJ9TZ1UjR
bjlY5IiEO5vQEV/9MuoCVQ6g/gAAdPXa2Z/JsyFYNzmsheHSRR3pchjTXLZ840RL
Q25UwATxHsgy5NsEvb00Qvig6kOwwgHP174rLMGynFnzkk+nmeghPV5Eh52J2q5j
NI3uVndmAE6o57+UywwHv/E5xnYbmGrbN7VyU/XINIWwcB6pgjUT4geC5bAnVBjc
YD5Nbq/Ec3DTrZ41AxgVJD9g48Ca86eV3OJz4dnJdMkUo11jCB7IHWewPRVDTiCS
c/yDaLkS9rR5e6Osfjwf39QsOobgFL7EmvcFUAkHhmkzRfLwvdWrSkqoOkP3AT0d
UNpoh11L/Ii85kPKQedtOwafEISHpBQbbClxzIUT3fmHcg1+GSAEiLWH0hKvGah5
quGAqtyUM6uG4l9VTarnNdSkROHCGgMnfhCSSTHvN4XiXIh2VJiO8a82NcsxBG1P
tq0QzYGaLaNLrUWih7qkzGZU1eEzctkfi3BI7DAP/6EWqxgsAr41pSqmuRGk2qDK
gC+17TXSXPrvjeDZv9dvE8rZS8bpuy9cGjuFDcWSrAXf2ub2u5KWpfxiDWOawTdX
I/N+qMZ9dk6ybzM7L2YlqNRvR5tbgq9W09uQ0V7aicqwd+rJjZCR53EilskQkS8u
ouD7+SzjghqOaZGBy6cBRIsEQuSReexiV8jX09C4aiqLW6eZGST+D91Oop83WtAY
UKF4I7gqal0fxs24X7QAhcW+wlCas+pT0SjDy4WZcVKhcUpqDQntLQiHL3C3ygof
utMXnxNesANo/06Uhw33cbM+qBfmrXjVL2XOy9JON1QVUHa+5aRj5PMLkBTM9Z2O
SWbA7J2BTZ7i6aavJtWlo34pwtvy+JhfdFSbwQkr9+l61r2Oo8X0VExz+Oi8B7Sg
Uz44wanYfuEFmPj/sNFaNYaccPNBUw0duG7KXI8hUSnqOnRN1gBj3ZNX18qD6NTY
nlkFyywzZIavn0m+yLkRSNKvsU6DX4VjujYpItCuhNMLwT7Hc7z0eyYSuofJ0u92
FBIxNwyHVC99ZtB57O0pFNm0gWebM1FifUq4q0yPrR/k5+jxuFUCx/J+YYyFrspw
bpiUI4oA0ZUz/BIUcwQEeo8t8VcBTMspkUV3TpTXPWQynifqEr2ezA5CfUT3jrzc
oHzAvFUYAPYWP6L8JQD85fa8EZaElVSytwFN8IzOdrfzId2lHVXs4y6qZEmabLnN
PJ0gCjx9mpOhmViBPXpeGJAJ1Ucs45eRkWHUdXuAT2aEUpPjfI3kIgFxfv/9JlGl
dz5nDx2YmJcIDu+y3fKokjt797T4bSavYKqcnFp0kvmIs2Q5iZvettHNzSqgPfu8
6L0/tqD6IwEN9+ZhTeN/H+02h6Ej3QNN4CqP3oGTKfdlxyKUXa7jquk+qRlbAjSM
/uK9Cu1r//pReCiRWOzS035L487b1YwezYVMxuxY+Nby6C9JTZfsV5esQBX1Uyi4
gDF7uP8nts7PJBei2AiXgoExuxL7rA/ozjjSPavq7NyZnC+r66UO+R8ioSmffyEh
mw+49pRVkxtj14p/6A8ZPx3AXaRc2yMaINm9HWbjSZq9bFz471h1OwYa871CSzAk
1s+eplgiGJyVKaKWOZjaw003qaQez3N9gwwu7ko5Nu79+qPqBc0WIO7RJPFxtygS
JjheeYfqI03WVKEIeVOQHK/FvN+VgnKzOvsrp3AiOKTwiNSo065FlJVK3kCC1l7H
sqlBL4nffuZnMlewAqlik07G3xEMurKlvdYW70hPIEK/iFf655ITs/HrL1lKO5Hx
UJnvqUUtU7kAFJKmOjoyW29Esnd/GPYHkJDliErua61L5seYADvB61bWpgHqShY/
LsA7FYHbLPY1qnw7uxOUEC+HNZz1qUYly6wL/fgr76VoGNOqyiZlX+5rBxMEPXgE
gBmM9qXgxCoNo7R+qx/V+rQp0RTfoWUoV8sfnSilau12Sl+slolHCxOJpiUi097q
g7NR9jD2HKRw5UG1uCDg4NHzeupLbsoVn1hrk5xJdZY1iKshos3VDCovp61xSjJP
X9HCAZgHXfC2U9sbUP2Q+xVebV8nq0KiEROLLmU3o4TsP/Cg/haPl00qRiejsINc
n8TUkzmisRB+SrQBFRAq5vhpCA/cCCaQVr//RkNK6JTCFWpQ5kN+Pc+bvUdBy6A1
bdUg7dYP6U1RxkDii586Xj37SHZ2nXAyV+HOKTdSa5XrbSVXxSZo35oZxzUWfoLz
+umLaapXt0DEtmT+ZpAG71Yn19HVjn7i/uGOrkqhemJXKQziuz6N0bYeKU2wMIGo
TZvXuPf/BaJAqRq53fo30iVhfKMmsX5a6AiKx9UHKUJ+WUolyvAvTiFdf5/pvWKg
5CJUw7QDNrZ1znQs1NM2vRk7qUq1Wmjkizdhes2mV8Zhq8iPELMbEzT/XggsDJRu
pU6ojm55qOMdqFAeBPZe3xitroH3Y1u0n2GQHRKyJQ3M9808QVNsPYD319NNvPyV
bZVAbck9jQHuoDhcS2O6n9TJeSSqoDBKlyv9bwqRFCJlgVS8t5j+wBBzMeflkK6g
mIg5lFl9j4X6VnZzLGxr1BbvfrdQmfmX6y9YNsy/sP03N0jLZwpV4qf3T90mR47U
OUG/91XeC7SGCt/HaviNEa4Q4jY/qXLuU7UkIHRHFfxH5dnatCs7pBPBkDJiZ4vS
VcntrerieCNnlh+DNh1PfTdliZRrfH/W5ShHmmZ4IMe26ZBKHZ5iHf8cKlUD9Bay
4Cu6kx7xo8/jVJll3Sqh0LjvVcM0PvVTaPR/0t1Df0erMuloph7TmdM12XCsCH7x
eaLQD1RAkxWu8IJLbUChXIcAZ8PVhOv6oaJJ9QDjPTJzofk7DnYW+0q6sk8AoLxA
h+uByed/9oqMT9Vty4jo7tWunzf69Uor+7Cubib2ia3UWHal/5C3YdDqBAtlOf9r
OrMixpUXkjhqUYgEzsy9FtApGBwAUlcusmWtS6KtWmjwRBrK3MhQnArXITqOFp8x
hTWdpI+HwCOnfkE62hrk30U+em9hi+fQ3hiYwXN6AUtATYfr2v36Cs6ieF1kiQIM
mA5EI1zpYMfC8cGoh7gHYPKcvv+trrM2grLZXAcoSD1ceJIy+gWWP0xuIgDqS7bP
+G0MQdePYEnY9KyD1qs6+8trgHCPXmRPUdeAxNcADKhS8NRj2nQ0yuPcwKz2rSIU
nWBvAEzWytv/33azODfsB8tg2SXKab3LB+rnGqN6RZXOoZeO0tIlsndNMYFCoIh8
zjBLOvNvO6gE5yvt/bnWhYzMEcSMiKDdxvQ7NGDAIoNExXlk/BV6S4lZpxjJoq/B
RdW9WCcUl4Da4sGtGlzx9xsPffPIAbK2hkGeY4c1ogGxa2+QMEM9Uuen7PcLP4n1
WFr3ndZq1yYGqcRL0DYE4wiijmr9l3dYQi+fq024yBc7GoAlyVn/ceadWwEUJnhT
fjzpJ8PwnpgTsNSL9ZCxy8ZJ3aM+4hcNpOaSCFhjfFawdRowZNQNLPEfo2d8DZ74
orf/9xqw+xeuNvJa04hEA5RgsZIEenjKzJTgIqdu2Ro4xlnwklllwNkD1qo/9jiH
JhBrURQNVXUUTBIu2Gg/JdGc5TmwJJZG4UDVWeWbncnk2d4hAbzZPufj+rRywmNy
K2csso/8B2BQBSlP1ZCV/orgiqCPMPpwFlJF4NMypkuGqyaiEqnNwobCxZ4mpI5N
L3ZjN1BeW7AYz4Axcjoq3DiVW2yxXizo/Ui8UE32tVmSsTOPTOazFkDB+vGtK4zz
Pkuq+BSR7nPtzfPcOxlCNFXM8FMygSwdK0bR5eUF4rk3LNH+ZuNQ/82xxKMF76bH
1/qApvvHfpzq19hZp9ZEiDEIz91jEqnj0mtRT+BaVctNWHIJbdSSARHmsoa+mtuQ
IO2FAyYqal0BlXaREjlb2AgERNypoHYgdQLll6zdg1WxS+UMX8uXbt8ygd1OwBqj
R/v6i8E+lfdNkNwG5W7yKaYaT7exVshb6yd4kaQmsUDAJk/5jMOrHXkxFexNaJ6x
+ayUBIsmXO0eceoYQZz7cVeyX38o/g26MCv8hDHgccAPFXaMkFcFEiiKh03FNGBD
6YTg8eXQ68VNORRosn0DDB0phvQeaHdFQN7sIH4RpaH81ldLuGk5GbVjOYAAxDUe
cEhlA4Jo3ZtnRpQ3TEF3Fd4qllyA470NYwDHYSfNp6/yX92vjXM+m2+lDpdVLfs7
QLjC4l3ZLTaomF1obsnSxB2XA/Xd3KHSOLSBJzIf6SlWNe3ZtJLUXCs730z7H2Wy
SxcstPxESLQhHaBEhnDGn28c5ryveNAKbsu8kTH0X5b17ZrPMwP8cV2Gcr8Eqi+w
UgjGo1FDykcTsh9LgfLIHsrElYK5IJL5YeqKzIaV/5GYn5PF1cvpWlT/rdTYjIT/
FHv24OYt8GWoC01jPUURYEBVfXbhuUS7n7BNodJcuf3ylPYBqceV4B8+Vtc1F3Di
h7IvArCbKu5Rk6LL4gLbQy1eP57vMuWLfl3iDy09FKy/k9ksuFln8dHNHkYuzHtd
dqQ9C6t9b5elh7HYbGns67JkDiLOuvGnKtah9qnv48B5OoPe1SPODoYWWVdnzNd4
ihiN2+lkyelLs1e36b1OM3Ho/g3ESt/W3wK65G0HCGaZ09w1UvFISnHC6wevAM1T
8Po6Kov4tfhgiKON1jaex9ZDQsekAEejMGMP507qLqLUSQL7hgFB/8G6wjJeecdP
/AUa5WCJ2uJleNkE28SvqsHtznxDbdcDMQyh2uAskFDdsn3jigsGDl0oChJHE0c8
uk+zSoxU5yXQfUfXWe5wINwNLA85sr3eubFNs/xcmV3B9c0vRWHrj4rHya3cZvJ/
WgRPBu4Vgd+DzHTbRwT1MMY32ABmnkgBIu/zLrMJvNs+7Y5ZhFmtr5q9+6yOhVpk
R468YrHurMzsDsEGQyc7/Y4V+5C2Op1iqqK8gCim2bnj6gGdMZi/4wct2VtJWSkg
D7wOzu+I2tOHRubUmB++2n5pNkn6BpFzCooyLcdY5X+7F+e7UyznWs+jcHJls7Fa
P+gDOxJ6aJILVANfqntEBsXZjdBBGHLXGn9C3wEN6fQVc5NjewzEKbixDaPePLFz
s/IGgkoGTlNExWCKIXRTGElLtoTT9+9pLcl7VWNnPvlGYzmneUCQAN+ukEaT2pSh
mz4rYk8Fco5egoPIFeXPw4VzqcA2MoQn4J4++kb4vTK9CZzkdLHsb9+pUEaF30ug
iVuJ78ywpXbG9gq9I9Z0/hgPJ7+AUu7E7JX+n5UW7F2H8GVToULz4CY/aDiWKhkl
9/tXcoSPfIeIbPBc9pcsvVCMtlPGaolF8h0NNcwzW5aM+VB+23nh0m2Ef+cPdcJ1
IrIpfSzShhhfasiv9oe0YmL+qwfSNzDf8Q4kMTpBbciQ+r3OXoBU9vT8u+i6DV9B
P1j0J02UUmT7Rh0J5hBiWv6EabxyiujYnbWMbB+OlvoKHbp6ZH/BtR1DgHGTD5Ri
6L7fdqGWXqzT48l9hOWT3qFIPVMM2qqVvBV9pXrCIu8H2qyqUCY0aG3zh2eFs96Q
rPa2cXT7F1mfP5hIm5kfFh3tDOd0bVSUFeOtbdh5ILLh9XI06ofroGPQHVzCOp+D
aLSLQ/mkC7aJQXClv9aLoGjbZ3bURWfrKHBxD+HoKTcw7uDnYXAzZ6tZwf1TLTCL
h4yyr+ipWf0DM8ONhHyGCSIeu5japVxx4tD7HeSYkZvaEfnzEh3rsq4lApX2Ii0z
jKNZesLBlYASC2lxEcj3EwydOr5h1+fmhvfyfgW4L2/wGhiQncwuKiYk22wrdJCX
yxCgv5PyE81qx3F6SpoYGCIWM/lOhPlEkQS6PI3+cmHskXDj5uuX/IKaUKYfo7pE
tSLQX1eIEYzQJs31q7sUdxl90qCPOQldO6JRPi3wr7MRnXuzk6gERRMm/E8VHp2U
qfn6trUm67kPxsFrxF25OmTDgsrBuqEVeuFYoYMPChzTBxLd+wT944I1VNUDIuSj
74Dy18mgBpa1QBUyfAV+Tm715I3QB3rLnRu6sj52vCNSdgquwwS/AvvVn0EIHynD
Qa4Vx/pVNYiE4zph3PfAtZUQ5QSOhUBIgjmM2iftgV7AWAk6dOHHMVZ1f4mUv77S
Cpa+jJtcwmCaNXI9+k4llSWSSGq6ogtOytKv9cSkA9ZG80q2vVweXZ1FU6wzM1uH
HVL+OykLMHHqMpUShsrKu+GOsP886Rl2uPf++ruYOsGXLROsRy2pt+WgDczgXQpN
UHS873QO5rpe2bTvBLZFp6C3a+nnxBLdPTVDDRENR4P0vthSBbX9fvrLI70Jx46O
b4FF1bHccpIMdT14EAeATr7WFAwZsMARyYoOVlQjiawGDAIdQiO6IGLz32wo9EhC
HirvYiedoSrugV3ey+re56HZZAnD+UKUNytQnooF6C5/GYvOE9dwpEsu42fuVQO6
5sxKGROX3lkLnTZJAcAenUdAYaAlc/lyA5kSkCJk4USRcDbnL1wn4HBgluZ1HoUM
wRUNYqIG6lzAxGWCBp4/l5/nFOPeBw+uYqVAL6bgyvsrkNd5mlyIwLjUAgC/AQFd
VfJ++v7w9YHDfZu+qanEDr+Aj3nwB9ygP4jL6I2Frm2/LfbLmT+BGlzTN8ifca6r
Tfy5zrpGhTsUby3Y+h30Am5GNhav8fc8A+mGGYq0fCJPnFSg1ffHdKTYAySNMRaf
PWDe9YsVMjAVakVQ0VAbG1IyGTuAekZpT1JRVY08OM24d5s1gpjamH/CON8m2puh
FrXwYF1MY3V6AkPohZgPqvwRdVTt6qeSIbmjWyzz86ED7QWtL1wwQd9Rc5mjBnLF
hc5T58mIwOU+Y3pLPOj7x0Tf5sKtqXKC/o3vWotC2jr+5fiT0NNnoHLeP285US21
lrvPew1MnFK5gycnInE95aJjDekhmTyOahhZjFli17PcerK24jF47Y9+RWtvTicA
4x9owFAmiqwaUK4Lt3lIY2mTrKMAZmgXhjAD7I6KwiTURW+5Cq87kLSUulI+R4jR
fKogNrVlPJBo0p4BPbT4orE6X48a9MuC7w3h+JiutlxULMIwZwaBU7Mt9Ok38ZkJ
SOXrkt2SAJBLDb7XXdBFaKAxnRfcjYZN7xDPOe+IaA2fDaVnSXLp4WKh1/8mwYCY
izWTLZeXPrPdxF1KcGtPAst8AqM37zHchOdrD0rBwaZDrBuvzEdB28ixzOUhMQXK
eIg9c2+kRFZSdHYPARNLOkLJY7zrAG02vDVtiXxlPKbQR/bFWZGKhb7TkklZc9Do
t7woUyCgGtxmmH+X52tTKtutfnBDJPWr8bV686k16c18LuvKr6Y4L4Ze73ll34dI
LsZ7L+1ESwCbwAWNG+yrXPhNwlvra2BzpzBcBW8Byhb46WYTLArrs+jsbSVFemwg
7PJSlA/mSQMOXwsoiVa2DPbKbAtAjNSmyEoCNicPMWOlJOz/DXZc4nM/9Mpk28hz
lGZtzIIp1DF4rqylXTAipZxWJmqcxJxFO/pIE1CVlxs3sf7URJXz+npdK+93l5E2
UbqvueEOBFUJ9j/t8YBXV8UrA3UqQEq+4Br8t1TCjf+jM0Bcdsv7ZMd7m8U5mjDN
0Xvj3DA7mQGA5yw5DdTLVdqERPmOLkzIhB96ARt/GvZdiB9F25HhAbnBJvlGFg4D
x6P+Bq7xxuK8yH4JYR7p8q7rO7PiCdvzPiyER/h4yP0AUoNgI2mgn7A0Loqbc1BB
rJdci4ET9ZZif5VmrTTCNRn++Mpq6RBsCuNLiIl595xUbhQH6dLt911rzQMzoLio
5ysRxtZFei+lXlOdwZkg2GJj7x894663Zxp7VAVx+CxrIyktJop1NJWu3LUmGPc7
7UgEF2dJ73vVAb3Q/20Hadg/9KtOEkFbMcI09ZxuBzeE42UVvkQBzDtxtqiddcVN
Y8KcNPLb+6Pre8aezAx9gfats/5kuul08J7QVNMdU0uKAvNBkadPvK83muAM/LuY
a54tD67vuIOe0Nl6vjqVUnpQRfMp2/xoAD8L+xKYbSPWdGFu/xH68Jyair7l/R+B
VCgP5WBDAuach/vm4aw7wxUtax0gJD3GDfwoTq9mrGvAgkvY7/FMMiC0zHefHT4m
96btAZ9EMfH8XV026GzWB8TZMkLvKM+w/YFShw164vUYHCqnVuhtqonxIQ3DN7px
477qq5ZL/T6PSlM704ghwcEqaKDnvU/3SO3npjgZRo1W3hyfAvm8VEskkvnD6BeP
tQzrL1zObBhWZmM7CxWF3zsckshzAYYpF94u/WXm/CDtbQxFr2CabAig47BHeWJW
BPHBovM37I2L3hYsjiLLjg/Y/AnCYJ5g4BkFXmiC3q7fwMKsHnCw3tSXPJV4ubQX
XjLI4TcJjG8rAyGdXaOwvXk0HVn3g01q7BvCDJ02XZR/fOImDrNNbwek0l411Gq9
iKz4ptSUYXJVNKLaBkBH+w/C3frbor5L1IELTTsn0q9e/FxlCKGG/5VFzPZ6OgBU
EBy3ouCiVQmKQzymPsrJoy7VSGP7veeKqzG3DgyvjlgncPP5iJ/vGoKEI2cnnR/W
Eb+K6Rn87RdJAOGHySoe2vt1rKf3t6Tm9JLyNn5h7EKAiojvc5JuLj1v8asS25Zt
L83oWNJORM/+vYFCA6NIyx8bhWJRfBaAAw1/cGMnoLZw6wWY+IeLR+O3ekjWYNFP
B3oz8BFLQjdmYyzQU4YoRWzfpqX/7Fzh171GMb5d2zPOtPhP2XYMQY3tC2Wx20yX
PxlO4rNPX/F+jCMCswQ6Jt8U1lmrExrvyWHiHlh2P7VsoZgt97cdgRaSaYb2Llvu
49wXqzVyvh7xjkV77iPO61Pb2ZtXh4Jw2BoA2YO/mTBheRoefRnO8ouWryWXf+7C
fbQmKbkstY+k8aDENfHA22PUMGJqYijO3e/+9+oOWJ5ayu7IcBXyKTs6zHQL1FOt
glr6THwdnXjcPU4/R1zCgcVI+/v1+uKE2ZXSbKSf1lmv6wUCGiZCyIrxUj99XrS1
CdGCIqHnDX5iIdn9x/vnaSkvxQHcySCEs3c/o3KhfBOilnWJtel8vlP49zNP262k
jI2GtN2L3MxkRhB+PGB1n40GKr3kiclyvbteaD2Ss+8ufYPBM/ioF7lJD4gNqSr2
96xz0uNxppefPJtUWHVZLjCi5ARsKpM73uYjH/3+xlTFopG6pk6PBlGewN1u8AYS
y8RBo4LBLpenm2N0jigHM5Xn7S1qDs9lcKsbtu5y8On7P69SqKmOMt1lnV5iWdHO
yP0FEK1XUEjrWlE9pz8yMujgpqB6ONPtUWGsyYAr6y0G1aNLrF/X6VVRuhyurauS
OjItvetcjaNRPOTW7x4ctwADZ0tqj5PKHu/E2iFi9W1VMhqwfrEQxOMVv3A74As1
hcuNKAx3dH0btQt37nYiGBqpSVVhIOdTaRcJNaUdtyuKVXixs1dXfkeXEoXOPA1u
scGNpjCzxodJOdrUtRd0HS8IJMyL4gy+vgkJGHcPTpzixMp7l5UrPdKZ+tb9/ohV
olkE8dmBiwlD59Rp2gdh8SQo1QPAmJYAC6xSnbFcC4hBir7QQDH1joLNtvpqpBup
fsCx0JG2IvX5zRwBKuuQjXWMCE3691EfP9+JeJT/u0UWD+6xHXbet470fGXEdy1j
4eGY5t8VZFSm2BjbnBia/Zi6JbJdkO1B3yfVVeClQ/BWmBzMqEIvgpOcDQKotxNj
kT5eJ1/cGMs4sUzHMMyBO+O7zu88QImbgRt9LYXfyfaTpI1vvp44++825WEY1Y0F
2L8DctORsdJXxVgD6AJbbgiJnRozH+ozCqWy1dulqEqygUbs2hLYsaEZsOdv0qKq
Y2z7suM25E9ab3QMs4SbISCF4KDMXf2LGqV36E0EwFYxrva1zHbm4QGq3W8E0IkZ
WKAfuN8WWuGGUh8ZWABnC8TS6CdA1HnFkvWD3+2NoA58ydoNjlgdNKV6ziDt4Ppk
Ywk3Ft5mEELnNGjk/n+c+7pSOF5bBhVII0Z0dEVD4b5JoOIR+i+tw4ui/0Dekeyn
1e6UJEpxeZHILFnVHXeN/5iX3gIXP9s+Randh8t9FFiBhragxTo+/oIWO6aMh96P
bTv2Go4MFW7fLT6EOzqgMUN177GAedVquigZ4ue29bsDbSpd10HGvnUTnedFPoco
yerNkfMdKEIubPOCsG7Y/9waihOgXNa06+if2T+t3IZgqzm1o6ZtitCvWwc0k5ai
FFJzsl8VRKzZpcE0eXd+W/aFi8tAt6JJP3A6KF1888U6eFdEHbJ/s3JdbNSoX4YR
bB2czu832X1PrsCTWjtUrtf/YmKNfoluU9F8iarDcq8uuoC/bjZ3nxtaR7KGN/sr
TNSuIlA5PG/pGzhfKkskpsBZIxZAi4cjjjHOTiHt9741jaoayf4G6l/6ku5E1AQy
63MIJLYZlWW/quZB7XWh/hl06vAlx/d6CHnzwPvkKU3np4ew0LGBaS5Bb7CJi7jw
fQ+VSbOLYP9MwsWEm0TysRR5bDHgW2OtHT2Jpsz0aYf1OSewhvT7jrgGjGwYzAwg
dC41wqo8Noszu2a0T5iIIOKBdfBp8u9furJZnukLz9qa6Rz77GPVhi2PRx5nkQfe
auOtMbITr52xSBaypwTuYz9tGzfqz0MbvtArb+ZuLFNxEPgsNKINjZ6x09vjhVu7
vKwJZqQQEU2c2S7SKCMoaFTLbR/XqvHRtRdIGSSjnUFQ3whKtCgAxfmkwH8dfPbX
FvCSeMvvdqiELA00PD/ufqvMCliE4IYUd8JdjkVdL6UGF0JHh3+VhWPkH30s9BsR
Q4nsFuHFbiQdiMJeoFw+IqpP6mcuQRinYv/V+Zkd3efuLI0qEjziPSilijF3ysCL
Gmx4U2sYVOErCq/zX4ixeOtfXPXKjbcRtIjrzFTZ6F+N4oXj66KZGYhj/qgpiF9m
q/tWVdur9t6QV4M4XEZ0dq/k0X1h9KWLcAZlTgiPMUW4EQ6AhL+MYayG/OOoFZ0p
EUp22jabjzAkh/cJpfXOojhbl7tEMF1hmGit9IfC1TsHjDhjOVXoaFqnKFNJWdn+
/yTCiEWM/X4nI+wTUsRrkmXMo8RbcM5Jj7rdh0SdSNuwV4YKFrEm9eswIB6tCj8e
MqDlHyjtxO0VdYiXXgsUdbA7CZnlWpu6tWtYP+N0Gdyt1xLoJYGtxvJau9umWqXE
6Nt0pWEfT5+FKlfYkw05KjHbo/O1zMcoSYt0aEuQd+4iPDcMz84XaaXWt7egkMT9
IfTmuO1zJcxrtQzCH7gWSBZ2exItV30rQL9Kk/64D1fHpMXIt0Mz05y61y6sl09b
7IgFFbi72WFAWGcSrNe2ZBNiZ5SXixWrLKXcsF6tRWscMGsSzT/sUR0WXCfn30BS
x0n+MvkRQI9Rr5fmbyvIe2ED56BWDPykCinZyXAGMrxsLUigwsnG4cfoLbbz6PiR
M7zyXF5RKp82WlC9n+T7DRit/cIpgjkBFssj0IsTZ14Ftv4tvkZkFidh1wRfPYNx
5SXUQOJpaBUaa8usKzmjJ4DLjNeI9n0FTyaAnUrNA0V55uXseJChgXAYnuEcLWjt
v3U+GoSEaNYUI1ywCRYHbIBno5UcFVKMWP8Ozyf8Av4pIq8uexjjxQ165mf4dn+J
zKvNxvEY2seVqTsOCeRkH4V69dHtKmIZKNx4yK1bu+BhWxVIyH1jwsJEX9kIOfWt
xA80/O0NJOAs2KeCWGSAeJDqGMTpjPoHW2liy1lzZ64iGxURTQu62Ci6YfQI7S2r
JQQ4+DeWg56UGRI6Xfm+vbwvMsRAGwdgk110vc03BUjktepHAGurT5bwOM4optCR
izwn8ZA3vFeT9Z2PqzhcR6LKomiEkeGb7oKd34rE60KUEaFX7LMlogg9Mdmqnnp4
iKlz6YVUyVAWbFkATHeVpzE7BxeET5Sk2Q685JXF207cyBxmp5+PW7kP69DLBE/i
hYv+/gB4ymA4pPWKxM2CjYwKsNyEb3aSGTl+6b1irfNZ/BA5/TUl+mHDvDj5sE5D
6lzyFF60IMwwIvrMJ8muVjNZ83HLr+e886k3+YhogVB3F2OBgP2W/uGgBi3NCS3H
09xTQtvJquv1UOWLBORm/hzFGodLypkjHGGWD+dYeV9RbcSHhEKJGzUzaXAz7Nba
LQqHKOfDNJEC/LuPFu7ExacHpgfr+mY0L14RxjTlsWgPH4VRg2Os/MNlyOzT3fXH
BWlixANWLL5zlGe9XN2qqL30Fqlw0GRdhlzBgjxA59G7CtICTNWSAOJxke9f+aV/
hL379sS6bX7BAb42ifMXcS5sr2k5E+asPwv6VlQrkEB92zplXcFTh5BWsdRQsf/7
WkLqhyJkBN+mkI8QEkyjXnHBl7mAyOpRKx4calM0I3USR/Ykjpqqfbr4EVzV91zb
Rc0b9QBcYZWisPicD2cqxS6+04eD8gLx3xEis5Nl2yWq5N6xXQ2Eb0Zl+uqZv7uI
e7cEKvbQTkK/na1eICqTKF6cAw3itmGLN28KAc88XvyakM3p8aB8A3g7yi9hyN8z
wv33F4r4ZEiJKTmlMAXsx4ldlTOB2Iz9jMt73iaigLlEzrX3ob7snUb2sCxps99p
ypyE4twGYrMQXKfrZpawozFIWi1n/s7T3AaUNx9oUBSyqPIFaw8cHVOBr3WvJJ1r
FdIDWuvWNiB2cFrxyv/PNqnHpMcBG9eu4PamqYn/ZUT+uGYYxlbypu0x8oTSuklf
g0HcJ+GMh2ps1rvx2K9kC+81Gh1zFy4vT6rywIs2YijOXhxr3IEFpcmSnKtE0YGR
5mGT3dQ+1XXBr3L0t+9s+iXReGrxR8eDQYZE2qvkjBX+oW8CXG4Bhv/i/9xm4wAz
vWEqBwpwzYJEgU/H9Qb8D6V5QH6oCtsKFhyR+xL1z5rSxmwzfX49GTOEo8uA8+U2
bb7KMV429MW/a1l2RrWmK4+j0x2gk8Um8RxS0/TjkBFa25G2Z++hG/VFDRzVZiAA
R4WKMofRTC8l2EbgB193A81QRU7lD9pwcYPeqoW4jTUlqIU4NDvY8xLfrpB53g0z
0InH4gM381tKesWvxyHAIvbpcieGNz3iZjvaeFgWyHEi5XwVkyuUvcjMXDTaGWN3
Hstk6A7bXXyUQd1JaBMS8lw/JtaGCP2+U4FcuQ1eQq6LD9C0j/PnnocqutFDkbB2
KtI00C2yT8cR1NogaLJdyCKZIskvtgbD5T7UWOz7lXsXKbUGXTb3U2fdm+uq7CyK
/3SV3WZDwSJ0c0pwIWBq5R8IgZZ7fBb8oM61NX3MLN3haLN8+tGVEec+nMqkXLnu
EPMcd8mVfifK3N/jKXF44RNZcvpJvcZq3L0B9VOnRPJXkmYRvzfeWnVMht+lqQbn
o4jGWPlV99oJk3aKKYDVcfAtaMfrhwjh8/oLWdjEdZkaezabbleUnzVRxcymJPrH
U6K/yJj0gTrhaKT0SkggaJNMchQdxo3dLCrsP3qtZ5qJysNKWc2QqrYNFaUGu0Ee
KYgnLErDY4mAuji0XbEcHdRB1S6GcR+xVIVTnEeZpCOLR7g5XPznF9PDHhYawsbq
rDSvt+W9cGEFiAGrEC5QbWp6Xo0HP3ca5ShUijV2sSqr/5VMjjIMi/CiyA6yccVP
eVSyDxuDwuz69v2J/ejuXVkS1RsfOP75WqMs5Dg9mMCw2qawTz4/z7NaQRv9X59h
JZrbuuAhU4+sIE53AUSZPw/tEoUYTDvP4vB/liW1XPJZXdEM04Qg+RlLwwN3zmPW
XQ3bpzIzdP8wlY9+Av8v7ZqFtabPCbOvPcNtonjtqocLuDAQ2b4z9V3fajficqTV
1iWacBWO9b2iRiu6i5N4NYDVq33HMIw5IQvybctDYqOJRLr/n7sZUuVfXgyvoFtE
Xz4Ny4AtJC3rAIiXWQvZ7695xKdHA64ohvE26Mb4TbN/YlLreKXsGoLFeLNiEDdn
9I97xQsO+wyechJ1c+ODr7jAqPZ4A0aOBD3mLyCwhrFnNLAgzbeBFuC2aYppEUxm
hBWs/Beu25hy3Ed5ttzBmls62ZxqFwnp/0eJx4aAd9HSH8nt7PVUBdLCXP367Lwy
YP+MU6dJkd3I2zLEoKL7mO85SW+hnM8+H5uBZTMo8XWc66OrbyXulEA2+wXykoW1
ig918S/sQ3AP30YCUdsOobuphNn1VzmmKRJr95ux2MFCkYPHNNotrUuv1FEE3jYC
z99v3RcMe7jyzFebt6zW0maBucjRTEmYV5P/LF5pKtkkJhhNgLHy+r2uY/McJWxZ
zRo4s9g21Obf++0ag6AvDQ6SZKQzBi3ox+9923JWnFRbTsyLtU/Z5fnrEZRMNTnn
6tClDe3gIz2/9fYX2q4FqKpG0rNdAKr5E+nR8U/VU2zmbnMOBeM9R7Ets7iuoOXf
GIqUs4ISPjFiyYtABSevw5ZdQDyPRyut4/dBN0mVCLGI8C5zcXOPcFcbyHi3G0To
JhT3ZleaTsaQy6BynTR/zwdGF0uIra3YdiTL7wrXOPiJ7JFDWxj3T1DpO7FrO9xB
5ZfhM3vRo488Wytso2/fLCLaLgR6AxpQWv2SRLX+Tgr8HIMxo6JeVHCYK7IqZ2Ww
3PHGuCek1P0CFPbRFeCJVqSTUr+58xP84esdxcst/waX1vu/e5jxOU3IcmLrYGYN
Jp2tiyO9pM6MhmbYSuwyEcSwJojKOI7/A7OGMU2nipjfN3P/Xuxgzc7hJE3i1URN
T94THpCLxK3Mvh9zDnAVq9pY91xxSvzzRRXGbYf8olNzRM1Rs7tyiwOJb5H1xabC
80GWPmtdVl9pjyLFuzcKy7XC4NpZhDLzqS7ZLMP7Va1NcG4DrIuQdskfpbwhHrPX
JzDUQeBx3NkKmR8YUVLu2XNvrQsMl5AOAlJleW6f7UU6h24C3T8i15r2cr/oanat
T2EcAG3P3sYNpMLa0TIm7WZws5LPVQoi4MM3LR029KQKSqZIaTml0OPRHhWk9bhz
dQZxU8o0xwIx9WNUpu8iSz5ABLhmi8IDsudaU1QqNF52m6tdDVKbbsC3UwY2WAu9
VenheittAHN1Dwk5l2shSIQtbdwBwY+btSgzgS6NuvkJljWzMTBpgkHsaGSSXmi5
T0MaP3WVVmnzzwKUnvQODx9U21Mrtj2irBGYlgZoWWGxx7hQtK1WhZxxRMXRl/oe
rcGaPiyWIMzuveimd3U8iQb40Vdd9D+vsRgJJZ49vy9sMPBvGPTChVBfkHXpI4nO
jwrnvue7DgwpGI4HJI7Eh6/biYpAC42g/YcbU3lU1nlToUwyzGL/hN4NOvB/gBDp
v8rh3PEkO0JZeD3bXzl489MZQ078baAy2qTRoRmq+tHkDODPHRDWUCCwZo1y6KZG
lMI4VVq3k6bUjrWz3ezAYjH6/MWPE/MyKwXTiO0rTdc44Tte0WwbVzQE9VJSBo9g
hLhZLR/1pt6gYY3DkcEU/ZvfGp8tX2rOTwO8bqFI0VON1VJHJ8b4s8LempKNa45p
IGCxbBywLZ60lB9UgV3cnnlAgA4RP4O4wN4L7tM9eqBV8QooOdOAXMGR4LXrzx2u
NbVnBpAWChmp9vwJ4gcagOeAku7uFmO1zDuojDVwUys=
`protect end_protected