`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 8080 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/9huKRhRMtvnNqb3Z+UU7TahEoHV+T8U3P3ufru7l1O
3DlgtZzb9QxCbOjthp9+wDkjygH0eUfDrEl1ovhZG63SKernr0nUlWkFQ/jle5Db
xgoNzG/6lTnJbaXWCF1k2QhD3yR4jx5X76sOF+BF9NEMxnax7Ao+n4woHEerZbH3
Ne/BhQUlmNlrGDYGKDQ3raxnpxK7ScuSb8Of7lJ4GWOtZx+VBKtdx7APjZaDuTed
W1oBS0ychfvBYolohjkKs37ytL+xR912fbd0VFYk63963jj5JP7vJ1ZApvF5NfcT
TwLIS7KMkf3M0uQSB8CZp8doz2hNTuo0EA2xCKhvS/AxL5j0bam4kDrHoQUPcEmG
pIst4H1F0+E+NEFdme9QJ7qTEopYaRChWUiuywK19ZRcc9L2tqJeYrvI/U8Lhq0U
wZieZdQZN6b1IKccQNr3rQs5gV3o967D/c1vsdvmQyiGFlso551o0Npy3St/L7+i
ZXeEiQ+WiXjSb/yYclOoaGAuW0E8GiCfz/63AShWuoaoPNe/9SvJrYpHcG2GXKE5
uw+0Nw7GuB8jHkAr1+tQ1VXfs/4ti6OOKq0MbNBboid17FHF9t9MMgTX8oyI+jte
xY4xylFl4dAoEAGLup28g4Xqlk0OqrvxEG1xEI03yPQtFTIXkfuMZKtf1qeW5Oyd
G9EfqeXJwwc+uHpxQkwnaifZykzdWS7NF1dNRhK+aex9//UuPfx7X/g2IddRsrkp
7Y0YHGXCRFVlDgtZdVg5La4m0A0rb0ZxklNFa1LwRdsw4k79aTVs8Ixv2bb8oDt0
tH6JvyiwebHGHXcBkdXE29g+xLnPPpPIYpsuryyAje4IGROg+hGjKZysZ0HQM1Sd
javtKq7lWDxSMffadr3oBMJaLJpYeRQqwGd9+hDmlOKIq1BmTH+6uiuvfYk3Ewx7
myQq9Eqh8fLogC/B0D+TVVcwshamx7699/2FPEjjrxBTgvkr7ZalfeSJt6ye/5AF
jwqqipRNt3qmvNSTky9Ol7crlDAJn7HQW4bvFdNTDOqMib01/wvZMmca4wj9Ts2b
RTCRss5HZA5OMwpoPbkpXD8R+25WbjbcncVmtcaDeJ1QIRKUHJuSAcGoNsAtjQcV
FKlP/xuwJQIR47YiaFIE8Z8U4oSqHgCw4if4NqyxCcgtLx28OEUcZ1JVeVBz2NPv
XDlYbV5aa4f8ziNgAScqhmRMvQIU04FjFVw0f0a8IDbzYvaVOok7J9DHVbvrvA6N
7LDZfyMbGJAHrzIlLulSqKhRyme9tbkmd3BJvWWkvw8MoVHSnzRW47ZQl02y5WM1
V8gMsgVp3JpbOuVakLkWfucTztDn0bU/3+Olv3YjWQiole23V4SBQbAodyeKLiqJ
5vQhvJ8qKxBdL/XK8GktnaigH3gKnX4QAfhivkxhhoBYwrGMVyEIVr5KA5US6Z48
s54CcoNhED1Ns99eHxY9NN4tOLAtmcRukd4YtmaJVq8FTg6PblJ0g5JMXUh804cJ
Vv8ugMcvH7s4VlpRFEGAB/YNLy45kp4FDh7zy04cgXweqJgqdc9BtANZDqKxLQ43
x36OieJK6C8++yN4bLkcQHQfXySNf6oNKIp9zfJiPDGXzCmXG9AEvREnJkG3D9cs
qjT26wD+tEPYLrM9AyywiRviLOSTlfGUYgXyJXePBtWb5cFpilI2SD2wYI2Cgc/L
+WhzjYpq/N4NcI9i0mchE/FOge3mSBSp5e/ODh63ltTogooZgWGnXIweG0lNss1B
iDqcVEYEHfpx67X2vWyf2vnIEXha62FlPAI4SxRV+hUt5D7up0aY/zFjKe19DG1z
nBDPiSUnUoeb9Oo2cFytjkNZD1XD4v73rKY5VMp5lEq0UY+/XCb9bYZmaPCDzqnH
RmTETsNf3vtzjYPZf5/uNyIC+OwvD0WXkrH9JESypGg2Uq8LkEsZhqMsvML70zCw
sPgV77LF1eWME8bJGAB1yhPzAe2LB/eCMTMcfB9hyifX3Xt53fui1hRFFRdAWe+B
yRcY7f+mdERyYaXzSAA+Pt0nsUHKJywUXd1+oKoXgKw+VBWg1AaxgCjtH03c9/H3
RcsYJSnl7m+m8g5i2vDQSNJRe+XOwTmj96zI4vd5dAsJdcnYrzC+UXx/9EF7xsiW
vCafC3AxSvhaXaFvi1m99EOSaJT/Pk3k4seifCSPO+IiPwWi2HVNw8P57iKffhyR
+IXQ3yrLpDJXy7ru8Zi8udmuzbxolUedGqeqil2B5h6VkuxsenIPxoKkYMIHZnYh
gS7dtdxAbIFbbmhVwM8QSn3TcwdZT5saG1J5lsIpkB0jgpigNhg+t1iXp454wNwR
rEn8g82+Zn6GXbuFR/f/t/VNuPsXAdEoYhszYXJssweIxUgrcp7dkoFQwUTY1Dij
TEuZOHMuSgjPf8cshshaGGRBywDR2H1CL2Q4IuOxJYxlEkjJ9GFN3oKgc9W5PrOi
gWLGHsH/hR8UHzCc8J91vV0YKlNo+rV1HlvJjAku15d4f8S4S7szW/OHhjuOLwUK
neT42ahsfnT6zsGryD6I0cOQy3nyuJ76rbVL5J4dhR3m0hYqYwRvsZFQrkEJ5ZUb
vshbc1dIFxH50UDp9Yd26ug2yaNhchLnWx63hHzax/6aG3fPrv0be+0+IrJvZ6rI
xbgTXWjcoEtd5EIyvv4fDu36G7RevyEfWRmLDzmL55iAeU/St9fpWJPP0ecWfvSe
MncOkwyi2QXWeQLhyFMqF/eI13c0/bcAwxXC+WbOXifmRIxl0WAl+i9/R3eN0VV4
GyjMtUh8vGPlT9IEMp9+ifSIa7BX4KMjdufoQAYfy9P0obWJFpcC6CHW9619VogQ
99meJ7xRrWKTJt32UnHMJk8Rt/wEG1j7ML3HhnrzxtHF9ujlwGL6M6+YLNiYI9CL
isPnKaj9aH4yhfv3VVvev9P0E/dlrMtpGPOEovGxoIl3n/1v5/j0y113dFb/rPYA
znbpHE0VuoGr/JOKKNEUPgx3zv1fF51ojT2ZfxUQJkQSMqyAOsXaSMwO3PgdDHOi
G09niwlsd9ylD75peG+LqxPvZYpmdVz402ROKSqIfxuVc7bIWRZGmAm1fe/ofZtS
XeR90RuHQ8QfrJNfUhOlY8OHqJmpkICUK/91c7Z7yPgdHXJjJsVNcjnUkyBkhsDx
s2w1lmOwSaR5/nb74sjT1fk+Xiuw+o+61lUIWlOvfo7qZZYVFtbFmkTltz4sPGao
A79Y3UOxbo/hL+Y0Nkaf/71sXzeg0EmJecWLVICqqPRcfZD/MHRrcVRrYkEfSIrA
ZC3rPZzzYXHy0rW08ZR5w6sfTM7qm159eFu4eLUCAZmjlOjgzbbHOuMRLy4l7s4S
ZevTTgBuBaC5gt5RJD5ymIGv0zWsXWlka8VhwsCTIcuWdkFw64P2fOa5/QomAUkY
9z2iy5f4ryxBsrqZZkhisnVJJ3fYLDpycr7qnT6lOKrUV1//P64G7Py0RFATBRHv
+ss5amlV8X4LtbVibfomKChFZqCOE8F3xVvEjeKjEoTbzTqmxOvDy9Q7S9D8dnct
YZ/UqNnbNvQ/pOEtSei47/LDDwogdG4bcb0+ay4iSrrlt7tYcXR1phhbECrpNxOe
g5MIfxQfv3Rvk9XAaGcA9AVWwuXoA8kOJmcL00Nz4rTXw7IOMT5GL2e3aLsF6ElA
N/s/fOkFeobMJ/kef4EiUo1puTYjk3mMlKBet6CoABwM2eyJudSjcUUtBg9b/n4v
mcSOWagGpp5svF0UwyOCGs/7pmYVLzUrA/2TvvqjxAPmR87XNhqhSQMCzovYO5DV
iXvyjnr0UUZgeVYBIKYOEnCwTWy39drtxweNt4sg/NYRvh51pms2IsvQV6tm2i18
2a7eO3NPo0cQMnYy57MPQPDwQA+G00T9NNy4eFuwTfFBcHjCX9gpqdzB1cxuJdjy
sF8hTj4F9A5FKyloCZkauxos2kiM/ftIgSo9JYK+8yF2hDPo96DAlr6ZAJR1LkGi
kIXk28FvobiRUhsDpTXhUhYdxHWB8wAVYQmebjDFPvAwU8UykkKMbnSgSA3VlGRO
7F9CfNqG83Rs53BfCFuv1oY5uH81c/XdksCiePQtOhhG4xw0ypYipdpw/wC7V5fD
sXjUp45vmHKkK5Ex2DaTiHCY/qvnEuZXkY5PaWdq1dQuk9eTY7KrFi3zBOJ84CvS
yLEktDCs6Ac3/QGig0+iq05sQDqkCPA3NTlcYX+Ol+I/h8+V2mMKVxTRiCJusBvt
eZ/3gm341IqDRB7daewdmOlyoU7b24AIXiVQaoCGiS6u2CMHgLieHI7oJ18sgTxX
PpljFP4Wv6nUib6JJS4KaRklVDTrtwAzE5FeG/sTwuobcPkIXPSgesaGCCdOnHlX
iiIn/sQRe/V7xAdlKCLULTKmKk/ega0xv9SAbsswNzUML+xHB4wM04sSKHHvJEgb
PCHM2j22ILiie9QJvVjbgRlWQRO2wK5ZNj6jCJ1+tbJ32kN/QOpheZDVQnY9efjt
tZEDVHuLb7XRbh/CYLcy33TkvIKeLfWxU3iePUvrFpGPEbFnxtoZiqKDjD3bywmO
kUZQMFKJV7vMa88fs00LkNr2lLgq4cDlak0QVhfgxLaZbXjpT7cALTLP2SpqYmyU
PwFV+8szcpWl+9ShDw5Ge63wADJ2dZZsN8UDZ++71D4SPzx/J136udhY1yQLP/Rd
S8ZkVYkltkjxWzI6IwsJkU1lmkIcjrnE5L1oC4+jiSmPZfIPfFYBKXOCPqSkqYrL
U5khMojD53E5cV7ZtqXtuRlYklrkpfi/aejrDdJXqsJ7bXcloipBeSmeffVTQoCP
dVg5fraE95uKMpFmBpV52gU12vfXIFTKwcmPv5lo6vgpDmHYOiKDO7GfOZo2RV69
ADvb4bH7xbMamD3cz8eOp+DhPxetns1ngTPfs/RXdZl0/TgvO6K9Iiu+4BGtIq2J
RJesozN4Jn2a9HC/eKLGNQB2elK9JX5a+lnrVPUKParkFDr1EuZiirvI4mCQpEzU
2QZQZ7N8A5pnHpcQvCnml+YcL5H3jC5XDduz9hQ3fYsEZWwGLqWhCmJT+zEiV0Hq
z6F0JNor6cYqRMSCWFTmCE6E/yGcsnUaHeHf6YBqtCNfaCN7PYG6HsyXqgR0QaJc
EIWK5dF0QNVYF3bIbifEWUrurhxV+8nIRgMXBgljqz2v4998SVciNPfYWy7eZfmL
JO1wuHydQDe3t2iJZGJG37t5bmmUIXG0PzDmEhj8s8CkbTrPW1z9Ukx5tRurEtwl
RDnkiQIp5YUYZmbc2dleLiXJAabNhrecPaIqFNZOGUzS2ebB/pLLucbEznaSqEvd
Iauiq3hbypMPOYuBQEW+ZV1J/0FMYNqh7esdwV98AF/ATRs1Y2814svB6E5fqDJ2
r2fQ9ifxfY9lMM5aD6U05XvpxkTtTB4c4fj46fPCfN/l36X95eIJQxvoj66YbZFy
8rxNilrhq1J49NJ0oQWwIcOUIDRZZ1vpuvOFoRfRKz3bF3Oi7Oh1yBMcVDKn5vpG
eep3zHRDJOcF9NJ2ikZhRbkfR20G//4cxoMWGr7AjL0wjq/ZG6elpLBf7yKdTNA2
mzRDzFgTslD6xWjb8+5hrxSEjIqltH0DuuWqy1XhG7WM9pRv7t5BAuofoqSKXH60
nf4VBhWq/+8qLjOIup3moBYo+c/vo1dc6PZW/fQqCs3SD+oxnvuKrmWMTefTa64s
I77JZ9cZpTHwdwcBUxXV4/W36pK1eFtO3wTYUeAJeypZ7FPWejYapt2Aeh9Zk9TY
6KQrk4feFCiR6sjQjfpvN6QBEJ1931YkB/lRmYYbB+s6x01q5gBmrnvyzJdDgIHf
xFsGmr6Ilwhdqe8ccLBY3GqTaXLTXJ9X8qfdJAYGcJ8DebwC98SScBzh4o49Tgv0
qxmx4CeJDz7TSH+uJhIC347ZvM2KUd4/Q19BtIzWFDj+4LvBdWSMTlacTz0N+Fzp
dn4YQnf6na+uueJ9DLwGoTz54oxqlrTdTjNxTGtoeUTInJGCB/FZ0Sxubd2BbQhN
Xz37CcuPKCAixOSPpYOs5/FYVBevQ+YoQorgQbHN6HlqqmbnKOAJoGkw5Ky38als
73EMNwfqvV+5Atqt2Wz/q7hghoX7VCO5NPzD9pmStutvA+eojMjGW8v9k+f1N+ve
eIaRHEDg0/znIzq31LCmXgb7Z4XE8xGE7GnKxF5tGZbgpt7Xku9dvVJGyQS5vYhP
cda4Qr/DcqBRz8SiwMrMfAW3v3C9uBZDcyRwXtmD2z2TdRKZG/W3ipN6GzKDJRL4
cA2Wo3D5YnRf1yM5oQmFP9DKes6o5/hxkWCYZXe9vhKSG3kKqKh5jXczNU8SUuj6
ulGyW1LjjAspAWgOokeGYodrNImDRW+JF2VbMp1wdNfucbGClgZ5iVInnvgOKD4J
RnJrqqpWmS80Bue2gyjcpuZViBTHxc1Xo7yBDgCzBW5lDKZRubSBLmqD3yd3OKgg
LaYJ807TJizyy+gD59m/xwO1BBJegZL9o2zZYx3AohM2/t2zUtuWa4UPnjTVhHEq
yPjktlpg2joFHx177ncTZngdgMdf4SOC3cAZbWtJnZJPEOmOLLsE6ndPLS4OzrjP
623uGdw6a7V0QfHxZGLVcup3rTpe8QbqxXgyILxKdeU0aQCbenhg1cYXVkpDxb1o
Wxx6/tzdQWZ2Bi+Ghxjx5Nn2vHvcxin6xM8Mii9/WtoMN4bxX+Aihqp/huNUeLnE
Cea1RfUDeOn4TmQxkGK/jh40gvSHvGhbqIOtNKWvFgcGzxXVd8Msw6o6G8D9dYdL
NDkbXLnudleTU2EReEzyUcJGdTvvcChwaJSj3gJbiCkzLk/jvPlxclVyiauTArVw
mM4X8dQ9jnYiyMfHbaKwInI/yE+ylrue2pToxpKJy+CvS8ny+u33BRKZNVnWaY6Y
nsDdN2E7yyWgoLNv8dUMyqJ7y1vetAcfyjQloBjKwc2qtxvkwUA3KZ3AyET2eJzV
JyAF25YAoTIB5LaTiJhmLHuWi8d2KT9pNsWaxEjEBKYqZkNgr3O2OW3vkMnMHHS2
T4olZVICxLJjUfwFjsQpjzJlwdZR8E1jlhtRRhi7vImdjgf525HNBvpFzXRHY5zR
gaD4RMSCIS0uk/jIts7o3W5fdj09Dk/85RU1rEzB9lTYZit4ozhUkRWScV2tSIFE
PeP1nvztt+mwCaJE3kBeFpMiCl8MAXisXP3UqgW0+fEqdtP5HZsGVufKvA0vmtRj
CHJvWwtUM6aBUg6xgxgX5oxfprQzmAz7Dq2JaOATqlZIGV5XjD+B8ywXZk+6973S
ArzzPNo1cj9Rub0L9678qgJL/U59rG2S2roQihFNENJY3t5wEXPk/UTy8N5kMxqT
bNIT5enqGfsVFpasIMpjpJCfvjho9dLc9LjX1qs8vb7CC0eGx8x+Ve6urshcvRlT
GKn/d0sKUQ0A7Ji44MlN4DJTDsHoYGicbBXgCfK7cIr6O2kXNRbkk27fhSXEhFhi
AYu4urAahS9PoQr/0wMUtzMxTbu9WZEsdhBRnsvcEpP9cIAmR171CrcUh36KNAcW
2DLeNK8H2i/LZ9nKkkIH63KpCjf/VGRicWLfkKQSKzT/Syb2t74i65T/Wqc0unps
mau93gCQ4AsJJfreDdvH4TuDdr+Jb1/vg44P1TZS0ytXgIRqKZmFdBNAuHTFVxtg
9o2vNQWhnir5wm7zuZ/nzZI5pryCsiALYat+xGeQx5vHCmYjpRaaEMV8PFZARvwg
tgd5dx6BTSvVZWqPz7PTw6KYy2k3iTuSEiOTU8cyXLNCoaRnQphMQGRWsPmIMyCi
uuWVUcNbclHYxJRpwRF55qvcWHqwYQEkCxQdPHKb8XTc372ufvT2kTY/s24+syo2
ma8JoLXJfLHxJoBOVv1HjvK79qGYGGnoDx2gaXGlR4dPkOw+4f+fKwNjxTwE8WGl
23e5GfITWGoikkEneifOcVg0HxJE87QLv83EqwhVFth0KZKTEUIj+G5S6MYuNMii
zRyOKv4g6OzbY2Ru1ixUsE6IVuE0bYmuo4McM3QL+y45zvuiGUojrxywJtQrAGwN
/129mjC6YLe8Vi4XE97JYiWLqcYRjYYWij7O8FWb08zNpthNwk0rdKB3gWIZveql
BoanCf/4sIumS7jhIdROstZ7W3Nbp92/G9hG5EhnRR7bl6nDKDDjnoQ6+Scpi4UT
k9IC5dkEyIkYrgQ6OpS/lK+YXPkWnKg7WMUhR+Tm1OAv0UWNxoXkDPsVFxKmEY6H
JIXaZVWZ78R1YuuV/hDzgAwWTK9KOPqGoM8rtoHmE0htDbBhBczdTZPyErYPVbIT
/WL/hIxgQDkYi+Irt+kGEqcfdlvxbjIU+Zfkto15cujryI3r1WcnB153revsWc+c
Dmd39k33zWaJbA3pWoafllzxTKyt/XU9hrpIAuu0i4ATD4e8RPsfJmKBFNNFMMly
OOCBwdwpMCEFU00Qidk2/Pr3+dA6+KfFLt6/YFl8YbllU8/MkpnEJKT0NM6qIyUi
sFAViQJ7QF9vQHqxtN9TmwuUVj8WMnNblm5FaKQcVYMc8w5jZweB0pq5e2AQmCoV
TaAwMh8iQyIHmUbBnUOan5xOALvUk5GpScwNMnAjYSbaV7MYi27Mf09k/qTjKWsA
Sk6Nzf5+cDltAwe2mBtoQrviBsRgKwGdeR6riTDOjLM1ITRoA7afmo9wPJjipZ/n
pUd89mRCYiNUtvKkHNYPMYAJf8RP0IK0eyN01WBmC95t/2Oiw+nH/krUBZREKW9Z
rnTfa01Ftlxwi7ZVAb71Uxe1XyF8rPBRYIpd1fu+X/PvMnXdchiZ4ogMbnacF/5y
GGUl0MW7+UGQwFUSIPvGp/6KmGOr39Uci7JYirhPc/Xn2l7lpVGL81XtIEw5Nu4F
np6v97IAdauN7SMqtii4xo3BWxGGV0vyH+19aCi7uxfGnWspsYHFqIyldPrCHWeW
64DfV4HAI3YDQbkvH5romhaS5AKVzH4GGM2I3l6opigxUVMcQDjA9UiBnfiOTJnG
7gaj9eito/Ia67wXfgDkngyAANyD2DHHfAHAjOf0Zg+ZghlsiUYuhCac4aEylixE
jR/+olrkWKM4XBx7WMIU6RAWYTbIsqLWdmxTNXThNaZarmR7PDBQfqR3/uSWnc3e
JLAI6veEt4sFQZO0+WF2jH2utgBrTRdd4cWB1LxTEIXKaurZgv7/mBVG1itcrC1Q
Z0+QGhdyTS/pI712zKVjGA8XRuWVXvGqr3nyV5+ZKqmOgLBpZegQtkH6Tt7JKVtN
gWziA265NKiwp/0xVQfsncNL2A5M0kSwnCRuV168mU9aXn/r+NteSIE1LijHwOoL
k7ZXXXVmTHvM0zGGSEQjDEmU+mvW1DVx3H4aP1RJ+miesdme0efKBAdcvAuZ9w6J
ygQQ6SoRsKU8j+KufRSg2NUrUHjPP9xyj6zjrb+/4JRUyLwP1TDGzbcy6fYQhuPW
QF4bigg5vqVKq5HiGRRCazOaLY/owjE7thhWZVOSKW14yw+Xhyn7e9wDFxT0FzH9
zVPI8MwKFt44ebGPIX8YmccnV6ZMcm0Vq4CSK0bepXprjw8XfZMt/RvQv8DfKDHa
MwFWWbqsmF2nTAAR6KqYbOaZ+77eJb6Cpb0Fd9tWqZ5YYkBE4HQRe7UCh9jCsh4b
MUPvOX7T8TufIxZYL6f7mDx3F+6HrsOTJxhpvIeDCaz+P9w08D/ZahM4QttYT++z
vwSZcSBApNtQEtXHK4QcxdSzkCjEj2ox5YMWRLNJbruKJTtNpjcBVL3fQsWLXKxK
Pr0mMLXDnctHjnyadwmyP41NyAqiFZnsBUl2PA54vSuQgROWzQfd0zLDj+8PUvum
OXFQq4tH357QWxhY6mUR0Um7pcLGXH6P/+5Q3ma6s4MRhIJo9TO941FC4pXipbQJ
Ju08/v+vnehhF9QPDAmed5y5QuWYbM9bEpmDZxSgpUXm7l8sLnPf9qimE1WA9mte
bYxMPcteYolTJ6OCiPZF0MlgujhynXGYBrLFqIt2/DUnONAsNE/WoMEdFU1hDAnx
mm/nM7smGhMaYt3R0Tfll+zNXsbZ/OcmN+rWfh0Ub3RquuUteBU0aCww0ZMoxpOv
P09pp7d64o6IsHPLQRpCMiuc6mkv+nlblCP+y/YprafLYRf+XBqnM+egqZpKUEr3
ThwRAu4DqLE4idflDYyB4QibTACNhK4bQghXPNRoQYUDdKu6tWjdI9wHaXSsCyEE
kjn559Ip1dnWt2XM5d91sTKlMwaoesejHUbhwAP+yCi2TAmXGT8NGsfsETu+1sMh
TYoZUxc2Arypdqgafa6l0oh7smjJ4Y/hwm6boNS9OlemP6Xfyxlo5noDIUf/NuMU
KiSg+tcxatzRCacyQYLAL8vGGe0vCQNfbAyNx4dqYrDnDwmNi1UIO0r6U4GeLVpm
9mZNNk3lz9YnDPMT4BgMIN292Rba4NrTFl6vOe9nuX2F+kL6f4/i/s1EAivpVv2f
7qgfamy29dUN9BRCn9dA3rnsf6Of5JLB0ZF3tcauQJZVpNmQUr6TcXF/uiuLsU5F
4jTiaval9Tk5YPcYMoBR8uFAXSHvkZoFcutaoj9QFxwzGh3kXsQjOCs0c8KdowrR
NfKPjcyQNNcSApXmyTZnCAINU/GCi3FJ63ucISyNsmRhPHG8bEm1CagfGDV8hXdh
BxXY7IYwBPQkXAOOjIxuSg==
`protect end_protected