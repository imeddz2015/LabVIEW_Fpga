`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 1904 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/9huKRhRMtvnNqb3Z+UU7TahEoHV+T8U3P3ufru7l1O
3DlgtZzb9QxCbOjthp9+wDkjygH0eUfDrEl1ovhZG63L3ufh/q3eXy/cDFwYQ4R6
DN/kHbeXKA8DuUxs7BF33tr0d8gI98hE7IbZ/F6Wj4aDnqx4tKc4KUhBLqu372FP
ouyBkcRO/OBhBjifwWKu0kE08X2TCQWnhuDLB6Dm8EraZ7V/V5cSCS8doYWFHrMm
QOSE0+qn8vXQUeT3Sx+0uVMQTLKhgpuJK69E12rwY3yLe1LmLhPfS6kw9dd6cibk
2jssN971/6Pi5tsUJbI+0O6e/Bv7nC+L8piX77Wuc6+Mt+jzPTtYJCAp9FV68x+t
X+UddvZmT9tarz7s1+MxqUleIX+z6W7fIYgucx9XAPJ0H8DfksCZb16KWljLbtP2
m/fS0Don/PWXGvyB4CYMmaeAJlwHlwHFkO2sCHjPYrNSqBq6+PRd6tOun0Af2MoX
TraZBGHxHg+4hqvyXS/clsmcOhZIqrkTkYoCxVmhFadTdq16Ek2XkeFBxoJkk85b
dq8OPKpSWinypht9w1N8j451C5iUPBe5Qmb1xknFgabOa+uZMfy9SyYLiw6ux1em
Pnu61TaN5B8LEi6dP8/LoF0AvnS1gsursRX/8762ZgQamEDFe28fpYTw/+lU0O91
qkneMkD4PA6Bb3+EnVJ4s30cGAjVGImJi98V/l1vfZhzW572baXf3EZhr6r5iz6L
L4fhYPbxY+ZK4RF2IeQD77iVgJXB3RIjva4REEa19nRCf7eJ4rjOVP8hOQSVs4E+
3ha1Ubgdpfbz1qWACzcd1m2r7l2sPub5JFKe52NA2x5Klhwa+sSeLlDM2Aw8QfFy
ycOGZFALJyc621jmXG6YExb554J6XJVmLXPzZLavXpqWbvjJTMcqxdEfWiiVDiYi
aFsXjov8MQCEIjRuDchL2jlm2UvQHL3y9O8f5/8YPMB1wZBQ/PCn86bKT2AE/ejI
03trolzLOjAUxO630XmU8jtj8R4wMJ8qRMxY46wHbQYLYsk6A0rjkK3tNvYAn4mE
fMYCfHt17mxuZp6DFqGOgoayMaMBzokZ/KenzjkHkJK1t+yM8fIKuBfbRf66xVRH
I8DtL8Jx/bZz5G6PtIKK/enNHmhrQ80cne43eM1Ifzph/CWmCtM67sJA5pxaO1oc
gmAB1Nh8ea1JuEZwaJo5VF5r3CpP43OQB9tbI2WiLmk1hmdCd6XiOqnj+Y/Z5tv6
Uavy31lI720buVq6Fy+gB05JysSsBI2C0Pjjtvalu5uTNpEjtNPCE4P8DwhOT4Fx
kdS3jE7BR9vL6a125YtN4Banx74NtonuzVjLJhXrNSvW8nSdhTeRA8Tt5kZS+57I
GHFBiR2ej1ZhNYpF7Ck8PYjI55UISU5IKOFdzVF3rzYteJjD37G0PqnA7u8Z4U+q
qvN7mA0e5GGA+myUZ8TrPASQNZfU+5IED9PbAnmV336SfHZLLaXaGfopRRFZmNVh
r+8K1ec8ulNm//6nFRSaukjHXWFibOwCoH/nsO9W/oYiMA2rTDpAi+G1pdwyJEyM
V/QmcfyW8jiheUpfuoDVGz5Por4xKsRLgvUMxjknSZZNaK5uDw8ea1ovPeVJr+CI
zmyCjj6f4WOVwFvwVeFjQ1keDz24GavAnv3vsvmgCQJsRkS0ffB7DhbubDoZFrcR
P5Hu631abZA/zQ2mTxWsiXKdEeYbqXeX/VacDSw7kpDuwxtGpgqTa3g4+Nyk9RyR
lYxdYHsefCaPLYvJ3WfYw+7w5k75eLJV7IyrVu8VmwLiM7iLrKNaTucWDKQitV11
aZHW7cEjfItErrxkHp4e6fyq0XVX1wrlTJ4MNYvjcCN7Ax1oZSiPURHRCxdkbJ8z
GA4nc0oOMDL0FmrV+XHOLVqEx0Xtkw5faaHGXNHDsgwXWN5hQkTKQLDnrpBV1e9l
mNxIe+h0O2fwN/Pfk0ct6t1ezIpR7RUoMk66j9jYyxfi3NWhD4oSuAgqLS2wUNB/
4Ix8Vnf+qY+svUVk38KeJEkZSJ264XEtXW9Xa+VCk18denKdbnOBRbcWxhGd8F4t
OnNeZha1oMqUinA6diMm8o1hfc8X1nqpjVmtiKclnQqOJolxcy3yg1sgqhnitKVo
fqzCZkSGTr+vv6Fg6uyHkF262oPYLxF16kzxANj+wrTtE0fC+P3L+pl+LBAS9NnR
BQJF5l2VBtjYpytba8LbWa2dD7PYnRmyWd0kQUArrCO92Zo0ksuvb65/ox1kM1ZC
kLdPcEZdhKI+Rv5Mt1n8K3yZ0NBUK7miQIeKldQnrQYn2Rk0ms1XMQzkz/GdsItt
r2TWSRnkdVeRDHPHCeOR2QCzaMFWSQLJNi0Difg1V8dEOrJt1Ugw8b0VGL6YSvb2
iTBJODmJ0oFqDF+PS28mnPgFm8Tcu8rr8fPCTl8ajj2yWD9bQ69qdfmwvSuUABDB
/ZXeiZIT3dQu2iLkPsq9qTBJLJPMf7u0tU4ZeyxcP68=
`protect end_protected