`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 1712 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/9huKRhRMtvnNqb3Z+UU7TahEoHV+T8U3P3ufru7l1O
3DlgtZzb9QxCbOjthp9+wDkjygH0eUfDrEl1ovhZG635Rsy1o6zwL9isw7JpPN6N
B0wk6B1M7oOJ7ucY+Q+Xc3KpKX5DOBnu39TJpA29Md/EU1G69F7N5pFZFprTHbvH
ZJE92DRm8oNaLn9K8eYDIdfIYOofH5Cu50cIQaJlybVcZOQ08EH79UuBHCjtggb5
jmXQwvIuiVpuTtKnJgh3sOWhac+5S4I1NjLw1lLlXkXmSEjtMkpeuXKWu7ZDiLq6
t+2Q1/W/LH6kxq/C8H93KPrHT/DfdKQH7LBGbLqU2u+VWaVENxcuzCN7PCbARUYc
dEE3JsdBs3HrQ/qUDyJ8oHi6ZVN6/zTBT8ArX81dGA6g0yCoVi1cBjRlBZPfuWg/
4OoQ21Uunh4DgH1TkWF85R01tz8a7i3OWA1lpBCpLMYG1gm10arEXn8PMzyBFsmm
4/aPFilDWDo1Z0AFFNlna8qCHmzXbooVE5Xzpr/vDuKzbTI5tCfUI1VI05imsMEl
jspNbwVwT2GxwYso82jGUfWS1g79p81mIFIke36gtROqFneJByjkSGZX19a+AVoW
qPF2ftcXrwLH2y6huhaBrFFKJV4NXd4L8RxwLVadiBHkfFmQTMHROe2I0LytUUEq
QZx6ZiXyTkl9OxFb4othGC60InwuqvrtW5WTR3oIr8zFDlirk1NBfVbamNSOfluj
44JKyPxL6S9SSCAkIN6reqLemfjFcSGS/x7hU0h69jmKcorqR0LAqXZmSIf0+wRP
KAc+ReU+WOcgARUbSQeHOxn11zohcIut4Y8/1QY7Xqrl2+7ir6+S3TCfCoZEa5pa
j5KlkzAZDWr/HHqCJZOhXajseFM2viZEpkfz9/TdtclMhFVn+M5w7hIu9vnfLI86
ad0Nm+7k3GarldULwLEBC6HPNZIAw4pTeJ8Nbl3MENjsdHKLJ6UX0IME8DiXhzaH
sdcPVf0zEkXFaF/Sk44ciISuYFut7dZ1t4uaYfWFQEt2J8rBpAXSmiAZNv2HiUkd
G0aONqvmZgvMbdX/vzMtK6BR/hx1idCp8WECPtf4JHldbpTU4oXQexQxedefkToT
gofbkTuA5/QiqNWRvaynYytK/SmEiG6Ax+liq5QqBK/lQR1lWmkPO7Hck8ckj/nQ
rZTZskVK8p8Kv8rEYG6APuTCNePJ9xjOifwXo8QaesGbNb8n8rK7koV5b2gd5xQC
hFZ/YCrFRShqcFvV1LLfkYbycSscupbnebvG9WTS9x/QVW/NT/IfLidoP+4kThU5
vE2domzO0R3+HbjeS5f+dAU3WT5mtOCEiNsUsJ+Q6qIV3GEDdpC7OooLDUeE4Vy+
90hhY+TIpBgxfOqnjETm8vWEW2tjO7aOSsEoy5WFgXHuWevFp5mw2y29ApXKfJ2F
1mqcUGdBmjk4U4LUZEX4kdx5p5J/y6JL9pz+NiRFK00RiRx2lduhreICfqqpLO2a
1DmB4dS4O2vou4ATdd9uGimcRPRBcoj4gYaB8ID1zOp9Cbzllu/4nOIAW3apUpYJ
tMFRoeemXc7wHSlHnv1knaFlLL8F4s2V9gHFAtSI08HQPHNqPaB/w+Q8SMiBjPKo
NiJp2/0REqp05XM/v91gYViV/9p/0IX/h9KNPZnAlOhuH8sqp2O1VftW6SdaAmyQ
lv+MkwEcZAVaQVdfgCIKChiVXV091m9OSF92znDVkg6U6lsVbSIYWpKXBRpXC9r7
BlPauEaisZzO0LZ/WIRVbZp+8Ze7fg4Mw/kzfEHTjvvMEB+vsB2Wu21zhnaJXAVH
yCbG4ToUadOfgZ9pC8Pn0ey3nwH1mrO7AXUKdQzofrAlte6mzQlEzI5Zz75h3nK4
0yhlrXblf9OlJI6ZjMgSg4hTLcX6/tIi7I4CyiGoSjG50OYL7+48utmNQ457Ur7A
1heL7b8h3sIZO2gdjpcE0GV9jW1seYGfne1cbJM/T1R0TPOTbliRLLw/yHaGc308
Y4fBy5MtfdrdsU1Iwu3hP/a8z7cGdyvPlOrxSbbVPzkzbC6yQhztAThUpvqypNqo
VhnR/g4YjStlvO/ndhC/pm+K4vaUsI5lGZK89WSXepW7/AI1PBJtj46l9z/OcLWu
zzSDXLBSjCW6OSou56K83mvrpXzhkYJp/JoEk+SefZxQBWJEgsl/OQKV/eay7WSN
Zwmem4lFXDBzIw0L8ErhPGGSwb2HX85X2TW4LC7PbKI=
`protect end_protected