`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 4928 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/59UwEX+aE7FohaWu0/8IpTj7mav863zUNIsgIH2BWb
Abd9opeuBjbGF/waQMI2vMJTwD1ie1YueHc3nSNpEh4OXp8P5ybZFY89uyGz3ztU
W1EsuUnchJoQgbHZ/sLbgtGRgsrAFn+ZoIeGN1d6RAF2wAESJmYP8zw+p00RvjZ5
bq6N2EMRDBNjFRM5Aaj5Pu+xsyP67QAHfOzogMxcEnE1OuDyVgnMhVOKJn5oo/x/
hGWbFGaQNtEFETuB34cItF/DVY9rCQZMNwiuqBSRcxb9ZygIRnkcoR1SGSBc4AbH
daiK4zpzTY/4cpKxYuuNH3cZXle5U9N2t4aqcgRHvOVghqUrUFxCVPGpD6ki0UDY
G4ymgKZElLsjnXoQLE5ihJOuR4uTdcoeiJPps6Y0dHPbbk58NK0QgHT/boE8QBUu
ASBtHp4N3vtGA5y9ddSVLaBEeV5TvqFj7n8MBO81LX0TQalXaw09Oqau8DyPW4Xb
PcsNHNJ9jaftFw5YpOpARfXTk0WiiW9XQ+F3XHQcJ8AqaOMkHbSUtHcIdyitrAMg
ghTn+6Ir10ZM3VffPvEBuKfLkAFwDCVEg99V8ucxQ+V6uehX3YcPQ4cfnf4L9bUc
FnZFRRqvD/4XyEhuHiGruXO4w40vJCUiErspE88ZLPy+1HWaV5uNqLaZ6JoZMDRd
9W4uSqGBEpEgoD8NvclZkTcnQi9ddhua8fXuOG9O6xlBKgz0ofZM7KMH7tNQSuMo
uR5lV/yS7fbFEt72WyIZGV7CbHTQZHJ7OHEX5JJVi5N7O/Ny4irOkM+0zAuMXSAn
S6ryDiBBp/KdkypKAmWkMptqxhQvRsJx8d1a8eA1suL8f5XCnmnBW0Ovhb9D5BCU
vGnyRFDIY2Jmpj7nzbwo3K/hFDD0uV08poUWJqM7U0zmUjSToW9gS6ZhZAPdLGA4
uSupPL1Ra434W3BhSIReLM+oyiRrFqRcBGe1ej86yJVf0KCRI88ENO3/r1PmHfm8
F6hPf5HK5jDfirzOGMgtzMhOzvWQe0v619JSPa4EOrLkvOgn0/2b0Jk1PRD/J43s
VCFnuCQ34npuypiB7KMFWojArLNGpfvvlT9SFR79rDa/P4U1KVO46f9wkbJcFhzW
mZlXVvaZqUTfeFtDxMrCuV/jIYanWn44AW9pBz4bSnmb3rbI1m/R28WqhT3xWVyf
mGc6GtZtTYIIh36skce/Czc/es2w64oV69CjNzooPNlezlIwtzZzPxD0vIMkbyju
3l5SOzDVz06sFEJoSw3+5oRlOtZqGCzomhK241yPtD8E9JQwKG6QDKBbnAbOpmiQ
tmp1mII00jjgBengalV1HSsKKtdm47Mrt7B0nUXCGrElYx2YN6gTSSB4+9h7Nk8a
wFdKeggYc5xB9AbR2HLwDlwEKO/rdUhnERYzQhjypIxla48Rq4mzBQSV9XYfgKnf
YnKhcGntZPS0sz8P8VPlPKwoQ0bHcDoPo/pgKXSYCL4r2o/ueKRsHl4w7xOr2NFy
4fHC5TWOqiU6BK0sD5DHU90ZmX8Y+A0OFbWwL4F0SVBdi1TBgs+hUIekwYPi8+uC
Szf2T2wXi78tWmrcuuFIv/hgJfYLEFB50nJhB4o291xvJWJVZTOJG1QGIylKE7Ds
RkUvLlAwMznp9nWQYMKKZHOXt+Z/668StnTeEDmM69gCdXF+mM0REGR3ePrZLWuN
bxqOtaZ4bIS7hR/FSwURQ2Sxmus7afHDeZsKrYUOeq6oWMT9xuZceytgoEMZUsKS
syEptNm1778ug3W2GsM5iqtXqnXsdAF2dABFFTjI+HJcQNuIffuRpi0z+rFVkaJv
KJbButbFgAN3N0FyiAs0BjGWZ22V22+SvasZY9K/K7UPoq9F3FhKZEuwXQkRLdPO
0B+EqPOKWaaSLngb/X61269bBPl2NLz/8GEWtZsfImQ+tm5MkMgRU3PJUaKKhvzR
O0Qz1s9wwfGefb15FVb4wJbUDUrZ1wodl1hQHo7iqd8MJMgmeNBu/wBNGanixCHg
nBlBjNDggrpELy4AGql96P9hKztVtaaUGuyDgcLfOwPqaGeyJ6NonDhCr3I6T7hv
pQqsvgxLnqRsi0Yw3aSSsEM0nGLVYb5dqItD1qSEqoP83vPJ7XIzHOA+WRWqdaYQ
/2PjeZMospAeN4UyLk3Y8rTK19Th4qeQ8z7bewY2pRyIbotV+vSinTU38Pef6jrd
AmQGcKD9ZPqj/SpQEAaMQEj2Q+1aexxRUc1LTSCUEUbw3+E3lZL9xv3XAUNoJppl
20TjZLPi6MhBOtodyxuSJlPIZO8r+2PF7gjcPB1/Wy3dhYqiUAfkf4PnEd/S9xul
5dCNLBgL3/oQhxvxwv6NCy1hYiHusCSL2qFLEfiUBkPYSWvhJtTdWm0F1kQrd8sM
S91hWt9MdMQSg2s3erWhgbbdiFyRAr+fLjVUuf+hufOl7inimi8JmLAoVC6Sp5F0
LVIVqn//4lVozNSiVmvs9970iiKfspf4iui7v+nymADUaQwSJQJWnJ2rzA/RjOv5
caZ+ehzOmgC0v1Cho4RHQxzekF32P0L5nMfcGFpWDT547wFMhCH/KDejBUmyS9Ps
ZIqfSmLRCtw+RU1H3KteOZqJH/2gv/rQolnoJTl82M6IYvXa10A8F/ONxumJLjsB
uL8AD8eUyMalNRwewfQLaKg5SqMzP328lN3tAoYFFGZNQToyDzgV70DkuFwOiWwH
uh7cbscDq0e7IgsSgaPyZibNdL3rlgrIxosZNE6CkAf5IiNZuTlFVdpFVFQkc/E9
GlLSs97H358f0HtxYWCNXPSX5arSaanUfS8XuAALFlsvnhPFqysE5jiIRGLw2ly+
HDTC3FUMD0mxxybiFbaRehNp33fa1dOaoNGoZx/cums95bdBTkDZxe64eARxzoMO
TXMiOvgjJH25v92Syu0iTs+F9NRsZTps3AmBEw842TZp8qXypk9UD/DMDoK94+5x
rfUTRzseKZbUshjggW6hD9Ah2jBUanwAr4kEfxni/f4WgoH6BR4mmv/u+VuqVAVr
C8ZOZvioGa8kO7obwyHwdKeVC/GLPOeJ0pdLMkrVp+JC4VKWDxjBrCriZ4hZrtPa
c6fWnfJGEjR8B/i1ag7+3gs95QzMMZKbnc0xuHuKcAKr1KhC20iaI3dwRMee/99p
oqjU19V1h1Vw/p7cSjR0PreuMssm0rjPQ/CxK8Zd4at3vIx84P90qiSgGe67ucaI
BQsEwuf4JWKMb3mURzVtNFlmoiQwD728mDtF9g5ngAFIS+emVl1GbWFVS524kq7L
lXHPrzK715RCLiwHMKaVwxo+H9S++gt8NPrwq7Zat2ZWzqkjpuUw4He4admfchaE
Jc9IwrPDSYF6mC4HTwJNjlV0cC9jKTGL3LNOAG0Y+8qfxrrKegMMRPVQBkAyQTay
X3+t57r7aFdVfMcIoBrPOZjX4XixMaBI+TFAiYhsDVwPtoY6RZvjnyxThLFpEqPv
/o4Wn7WjkGrjDmXiPc50VWJ0MxIDWRzzylnnEFYQQ1wK/6B63grPMXNWELtCAKt0
t2HTbhsk2D0Va8tVB5JNhN/8JR+yll3gUIuHYwcna6BJr6imYydNdhXgiuvxshY7
cYlcP002hf55w7Dwx0Qm9WakxIMZ11oh3xHs8R1kKtLGK+JPxGrOuYt8bMsceiAD
JZjPVi6AAHqFmBMmLhFAW8luGxgJg4hhkSLDOVoJqI/tXDBUZLuFOXokJltVX3bP
FenBc7Kng8G8vcLtD+RHp2bCQziaE1xkYtU5kiZIw7oU2TpTAgGHmKTSZdJ7thon
yVyCVrLO0MD/UWWejo/Nk69BLvNAzxDQjNkp99ld02weLpcs4ezwFGV8qsAXE5re
3mj+EHZOxrtg3GLbmMhEE1souUYeAt5bLa1gWv347+0EWAP/u6KFzHPjTMixV/It
6v7Xhx+Rw3z4wQmujaYwu5WTF+5joGNp3+/WoufAX3M7aDrUsiaV6664PwlxpE+y
RgxPo1OX/MdAgv3McmiEwI2KEbstTeK+eHQ/qSQ6lOWxfYFUHVbWrKRFOJ71tp+l
AKRELgNEhV4ioU4WOMyQ8zkTBM1EuuSHBti9voA4itNoNV23Yly65xAvjGGSik6y
R9sQlWMl8612lrbKS+ok3GlM/ePSxzVEruwOGv7cLLb2AWXoeXF6q+VG/jn0jZpv
M3j2m7A6UpXC02khOpXXYLfAu0fsGK/WZGW18swA2snoJSwr12+zQPVc+IjcE/jz
91gkH4h2YDeIpNGl625iWrooqzz3scYJuDD/tXnM8z2b3wTyTZJZiDDS9g8MGUvE
gspc0uW7gpmHH1QeGdklaAVvkFuadf9vmPxJhljuTqftnZ5AWNxLbQa/jrb+n6yA
gybKSw1YWThQTG09166TDhNWJK8IGy7hn7dVAAsa36ZSAFgzNu/1zudo3FIdYHD3
tX9UjOI2ArNQ9tvh52CUSjEQ/+tMepO75f4VyaBB5oUWbG5o7mrdBY9SbYf3o32R
bgO7Rnbrn5ud1/1a2i8VU0/tJEbnwZ7Y8/Of6yCOdwZgifb3rO+53EOCUtCd96Nc
bqDOCjTyZcA86ma56msuhyY69loiN+6qpxrUiPDIMQ/37P/HuVw4mdZp/UMVzpoW
iqlvYg0CGzo8rfaiphoSkx85S/lchrtazToZLkyxaappso1sLGtQJthRLWJxHwJz
tg59EwB3VcaIv95OdUOZ8aST5mNQ2BPVGaLm3AkuSCQU3Yclqys5EqZEqxIK+Atm
TBEyJEg23YUbM3R7FwG0yNTEO7rftLvigeCcPC/CBvtbzR7RiI7Anu6xxtBdnP8j
2pKlhhwU9N3in6AqtV51ykW1oKHIqDYfykoLcxd43HK0eOvRJ/JSg7D2Z/YCFdkx
NDYksBEmCtOGQwNmt2NGgSgpG1P1P/pBo1ClaImo1xdIEWjxUUMXzTZET1cXr/KT
6iGdk1qT7fLnr0Ec0rXQAbLzoSexslmzwLqMDOn/vmAGkhoT1HHIeTsqX5ncch3t
0y7qtyJox/+fW5JW7Ypb7YDFTFM+h0HI6dNv9Z7+2RrN1aRgfpf7t5NUF34mVlg/
3TaRUBVqQH2JkhX7+avU/O/fstfOLrf8fPx+MXUIqSs0OioIWTc/4tg+NmRvymN6
9O7pi3hrfVqGMQvmWPQ2A1Y4Pw79pEncHwAFwKR50I69GVHgeWnEIaLOxhxTI9sf
KfiznvMEzcYem9rX5QedlC1o094fCX3oRsOCvUFjnEtqynvSRSxkjoM8pychEXYs
PTY7yh6yYRr8Ib//74qnqP03Q4+r4SBpl8I8QoHh2+9t5Dh1Od9D6/u1CGj0LuB7
pJBR7F9pp8RQprQVfzwJAZ2oycWgtGtpua70mWzXBRRDPMhTrrOtrvt69XzplXx/
k9t/MDrce68rqXCTwtH6rNi/CXS9HmKASf/ikBgWyyVVMCXiI/rrUcYjebWf8oXi
uCuIU5gHNQ+vLgiazCA9JtTIbFUbXOYG/SAeBIcyi/G71EmK7MwBSG6BfUdRAF6F
LbR8ybPnQ/+gQISn+0QseDjKAm2RlgAJpapX38Go/HoJWTuAZ1FQ6xhU4Fn7h4Ai
oL6MTBSPBio6os06ny+XFR+mCzKEWsslSPiShcDNwG29qZgzK/v04NUkRvuGT24t
/hyYdqgdUxKaZriXQf4U0aPRg91b1PB2sBfex2pPc4FV+1bosPLcjOK/0eBrhO+M
j3virZSGTiB8UsMfOxMCiG5VtSdLAa/G5e8HQs9lfPZmp2RO22f+ZDK3/Xl1tJjv
cNHdPGcGExwDOT5trjnyXLnZsoppOpcmhrFgOP7DTLpHxK3e/n0xFHitkRnF5JrV
C3q7hDKqR9s2CUYXfh44xLcbgS18d8IeDVGKaXOuGhhQdy2s6Pcdermo3X1O6eS2
ULk2FxaCAS/zbvDaFeePrnHleyIl0MdPgGzFmlW8p5fFYkxAFrRFYs3JFD+eW/xX
27MtoImi48/ir+Em1sMK1y0i2AXo46B/9S5HBRe6ujC+YLyYB/osY0pw8tJ/ufu1
AtDv2SltQSqHCJ/kd/+GG8MkMgh33zg9a/KNpLf0ybSd+R8T5lODNfknpG4E3ooG
90vppfwKAFqn42yVwR7bOakF+TJlM1r+vV/UsNYMVdXorSIk/1/QOY2I3rgXI4Pu
qUB5KO0Prh5aCtKlFuNQUcL7b8N4IOSFySDUYPH+kG0YXMmLTr5qILEdZPvjE8uY
JA+S0m7Ej+5T1JsNlGx0ZX1Rlcblf2m8gD4X34ecU+ujbaq0O9slR/3iwL8T2EoM
g4X3Dr82SY+4g5EJZ6VTuTYgV82Lg8bZYFZJyNJ8E7pv6dYpF/R+lQLohtXxfLY7
P+ZwY1Od6AKAp2gECfM05J2Vu/9e7JxYzsAb5PhCRu/x2NuoepL3lezBiKwBCfXo
pXCuCv25gUchvyjqCLpwlWI2fT+ozD//nr4W47dM3uDBUCt/j7LNbFUk4R8HuQ8i
8ebbVwzer5Kzb1gqoYzrTo/4LyPvVpV37e0nPsacHz4=
`protect end_protected