`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 28208 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/9huKRhRMtvnNqb3Z+UU7TahEoHV+T8U3P3ufru7l1O
3DlgtZzb9QxCbOjthp9+wDkjygH0eUfDrEl1ovhZG62OOZhknDkJk9tIemCMa1m/
wOxOFzXmBef318pKGFQPAjUkMBM/bBSe5ecPJSavpyJsHVHykIiWdZBBCiu/0qxg
mgdCkl/F06jeoXMnh3IRur/ss76/GO1V6P2zxI21h5W4OjcacaqYbypc0lFiMuMs
Rog9ho8EpVv1P6Et/eAO+cwCWH62GsVGKypmEfaWWUURQ+Ovw8s4HghL/FoX+tLS
u2XnY86f3c5IhYebxZzIw3yooGCIBeQyyeSM7MRmk5uPISKLJJwKhWNlHOVcz/e0
0JtJ5PZQDe0TChqqotcZLGtD60iN5niDE+O853aNP9Oa7ea9Wp/cj22aa3y1Q40Z
n/lhPoU4O+yfvwsPMI2MUs9E13K6MBv4m48mjpN7//i4lnwc7W3S1FGP2qR8KXy4
NeBdTGkpagidarhg7CjmKiAJlYyBMK01gH1wP/JxAwcNMtfMP8p0349AT28AxLym
bBPCiinH5k2+GsFf3IxKvQOTdZPFsIkfWBksmxEtnzWTlfD/ySYZkiWWkcVFPCpp
LyD1aSJASQegFWh0PijXLEDR85+/9foyp+kGrwfcR6QV8bW7dYeFa9zZS644XLAy
vKincvHhD9bheiCU4kpy3PawAONFoGzk8Vycda1Md+GPWhOuIgMqkX0r1DyZJj8w
ZNMHsLJEDYb6bP9AeZBFSEzPSxPM3t9mHeNqSytjBoedu4MgA6dvImPQUIqlvyqI
O3mAy82R2VaCQ6k/EesKE2Q+jXz7R0zmVoTMGrMqzst4XwxRu0sSZOcYycG5TV0c
si513BON5bGheYL+KuBrcT9WoSYJloSiJJZV8ex9R4Z8y6X+G04j0Ap7Q74vmkgw
OW6OhWBorw8n8HW54g0fC5E5NIp2QsPlbYmBTy6wXzg350oeQSaWd8+lXLcv6Uxd
vrRs+ROdylucu/676ibUVUcgrkdJ6NEwh2VIQbxJT3mGYnRUkWGgGmRUtD/Hweop
UnNzpRBTs0aNl6AuOOWqKtbxvMid9vq+pHwrooR5Lh4u+vYjwkjOWB3oQNlWYCMO
r4KQhVn2lSDD451D661j5Y8vIPAnj5G9nPRU32R5TOggLINv8J51vBP9Fy2bm4XH
t7k8NzDX8m8mqtv949op0V9pLBEvvUrQthpq3PHdzfMF+1HJ3Zzliy8g69dXrqN3
W+YMMq5/RCwRmwA0GVq9updPHIyC/hP9UKuZEUG9LpsFeqmw8tDHHkka3mgiPK21
qKegfZzMKirl/AMukpJyK7cyiaxdrIykwqNCpSKjYeyZOx9Uj/j/ZrzAT7Iur1MY
mi6kmFqMsO9Hl9OZemv+Iqnn6iD1WQZxiskXXSm/vWsDLYd+VZlQcK0K8HQ9CZU/
OPS/5cizzO6cqFk4STcW9ypTlft2uDCxs1TGszsWKAjy/DfU1Cvv1briy37/X5TI
lE+Hd6iHj09S27nQMuTXOFUgggfKjVaiwqW+PfelZz9IqzUfF2XHkcbLm3ZrXNgn
240TwWIb29xkAgga0dfyxmWndtdhE5tGst9ulb1V/glihYPDuP/NdOKfwNRr+ZMP
HiiLduh47eupJV9Brpobx+p52iZ5F2JNzA9hk8L5pP61c6y66T/UXzQnv3GMoNMH
ByA7bX4X+2S9m52EoLDZMLKI3kT31pL1tW5ty2IZP5IHn58TSvi0KPgLztxEwzmn
vKnGIywhuYamo+uHVQKZ29pTRQ5BIBPfwWTkNMotB7VMCwW+/wpzdRHWw4tlNRgK
nQfpKjvRZBPPj3LSFATF+NS7lYHPkgDKavmsZrI12G0xTciE00OVagNRwZloocyu
66trL77cYayBQ1PI+vdrBB8VYNOXwQLgQaTu5/rEHwULxzoAVZkdxcuuWKYVBrI/
7o+oGjwO67oNgksq+6aZDK2IZ+7aAznObNgDvKnKfdbOunp8U4zFde1BABYWk828
ZX9ylT+LlVeRQppZ8KWkL0rXXTSsspg2lUgH9PINy3tjUIcY6QfoahD+B9MZPf0d
B7RCLvzY9BoWpzguqG4CwIrgc6/hKTfuvMKa2xuWTs52pnelMbRyFWehq0Z397um
G1LoCY3ITqmu8TUvPKUkWGNIqfSIoUreDE/ZXCfQFG9jsoPO8Sza0fs3xbf+XYFv
0lqBrzYY2+3dnzSmsaFF4XhK5PnDB4nSBdz/7Rsd7diBkgTg5cT9l8igOALr/aax
JDPtELmQflDHm6u12Z2CCA8gM2xIS/E4hrdnVi1Fu5swt4dsrACkfCL6JOxS78pG
rgQxHnmxYU0M0PoAo0AQ/oXMlzxX9mGe8YcEZWPyKIIakbOEvfrsJkyrMU3/d5HP
84hBJMN0GASusX0UKASqfPRsoD4NfepkR39ILqTCluq4bbPSZ1WEut67xVUxghKx
JXUUCd11r0PPxrsnQ1sV3H3ciQ98UCl43vXO/pnM6+TeTUYSr8vW4cljyJBz7eHu
vXMmXbl72gqyzwzlbpCKlJ0yGKAAaYOT230Ade50MtR62BIaCEviyjiHEX31C7+l
l8ITzGwtnVL9INNgJIL14eIZ+RkusMBihGVtnrEH90xd51ya0deZtLRHRedHovmf
pcPhfjl4qb+d2BoHwQFbugEiKfRdT7ltpO8fZQWwGZu+U1Oc/XAeHMIrrTDT7adq
Iml1oTHyn9vmk3dS7ndOmuw6JixeQCY7Vf+oZixDmH8S5edB7NeRa/blRbWazNJ+
UEfVQhNA2GjIpfggmwck8oaSiF8P018R0DZlGkIFS/vUDSYLFipj+wMQLSA3tvrZ
Obtgs3KYz5gHkWOhBffhJeokdQJsTVeVIgj7oP4a2doZemQr5cfoTE8PnTVYuBJz
VcT/l/Qz+KfODyt/yyUULuWrhCqYaDYeChmY04FHnVZz3KoUl5ClIVE7ZvPuzpTN
gjmRZfX6FhpbsbqKgq/koys4ld45lLlRR6Ox319ADV9Ynh440HoPn90HYO5NvMZk
6Fn3eD0Lq+zzDf0p9u/Xa/pcI4R9pxe30lx5nuh0eYFxV/5GBaAs5h8JXYWGwyq2
lRtQpUMoIvAqhK6kaleW/+DqF7NcOYgvjRTq6PMwov38oH76Nma05RyL6fYXmMo9
Q/XpMh6yLMTi2oOhDhZQ87/vmNERYoAsX81XEf/3WTL+QdZ9LmCoIMYzcBeAxTxM
HtS8pgyDE9CQs0NBAu1ruAtOtXOvByRj5gsaqoC5lOTav+CtIGR3knDjg7q9SixH
a5T9MeGSV64cLjCbsY0aIVQDAH5e+3Jt6y9SXP+p/WF7PRD70BwzgeSOoztMH0ki
7HswAp+YV3rZ0bfW4MVLHG0krnaxW2G8OGAGUEY7HlHak77VbYKHY5sP+hUdADtB
gGw19wGj3WAqQmMkl8Bz/QCrKDxShsXpHIp/lHEn15RZcQGN+h5B4/mVWg118C47
LNXTQlO84l9XptIDm/8/jsFtYxS++DzdosClaAYvtMpl1uNNzFZJ+1AiE0DVyRuo
TgETxY/pnz49XjQeQnPJ7D2SDa8Api5LiXSjDi3nY3lUKEVgYCX1b7i6/Ud4W4S2
1Ofa0LLn5OodykoUyc2d4kq2Xk3AdQoUl05opWBKLYxGasU4883d7ssZ9S4RDmm0
Vbc4ded4RsZKQdPwrPVscERdY9JnR1eYbFSQpheyPCcUxFueGA9CflYeJGHxU9G8
OP7WVqeuoNnwUXNZ4aD39cCBwZjV2fa9HscUBUHgx7OqdeR+l6kbms5KfDn7xVMb
I8HG0faIqY3d2aJ+NzOA2XnoF2mmzBauBcBK601yM1pODpIUuzd/CyRzrADCC1ZC
A5nfy8g6qMJID/tfUx4YTSWz1ZuEbMWZCNbt6hp2EEQ+OVcSpmmKh7Yp+Gu/iFO2
ngr6HhKNYz52KO5v38Mv0eOLnIce0fN5h5KvVcCbvDQeCo4JRxcZqX6pPpd3IIVa
NzS5og4QzPprNKPo0slkor7cTkrXmg7ixDyZTdId0yTMyDg0zs4Qq2b7O4pgRimR
VvocPXpPWopnP6CEPdBENKucd0VC1sSWq4GcaHHFc2sgQnE3kxE7ofxg+zSg52bM
MTuzQeX0AkVeEJ+YT2fKSVbmQpPCP6631NEwlZSv5de2N/yo58KDzRCnDkXtOqdF
M120ePMPH4atVy0DbBSWLt5wP3V5hvkJxjdqND34RMXm/p+lU2foiCaAmR/wzFLz
Cee/glajTrOeH2K5KYxaNNeAHlg0Br/mmcRXpU6RzjYtNlaj4+uhYI6cNGRV3AO5
FWWgrogaQi7KDXqOC4LtI3am0ktIwgE+FJod2KBGWNNalAP0Hjl+OIpRXIpsXnRb
eVjniQsuKdPgeWS/FWIBZIyyDOdaR5zvIbVP4INGJF3Cm8Y2XaQe60pElhgnDMJi
I5Tz6tOy0e10JgjcEqnpoihfzpmffrvBU/p6eaWthEum1FuVT0PfXfD8vD71/mtB
6Kj7+dYa9s4r3iCLDuOMURqXgk9juptIkPiJU//8O2o4mlnppo/X6eyWavRge4pw
zqx5XreijdUt8gpS39JJJ8Kg7vetN4q37M+qWGyAFojfxY2MOtfpqJNZV2594teS
tUy+VGyKFf+ZaXkSgGgsQlS4n1tePTFaup3+ykJkOtPPxfADjha2/XLVhPlCB1K2
V2HF9IfBUd+30AkbrAKCLcibkAQZa1A6BZCf4eJT+z2js/MG9f3WXb/eOz5U9wTj
CRch/Q7bHnsEC1p2BA1dUd38/Dp/2iuf0sQw41nIL6sAzqHM7kLFRiwIB+FyjXNd
0GQk3iAkEPjRqfIadjX2ubHdTyoL9NRfYQtwJzcHioHtTowH+NMdztzwnx3I/IjL
Auw4Bu0gX0YFRq101u3ySlpvNzXlKdgp0mtcxxR5vKTLWexPHPWwZuXtxRC6GLAK
ktrXNBcV5ctnqDazhMauEabQOq1RBAG085xsOtBmFeKdqgHnClnfDDgLedN8oz5c
11CNZaK2NIXlMJqfydabD4FRx1DFyZrQQXJqc+uRY+k8GETGjYplKk6CXkVwlHo4
iIh36fcdbi6hbWEUxZ3CM09QphafvFWci/paTtN2R3Mw+aEfzHyh2ScH6R4il7tw
g9GXSSQO0lr7gPlb8aJeMBVGHcWSwpn9/8lVeFz90UqFrmEscQIDnyjB0IOgiqCw
B3rVANVKz8mjdU/cmPbcFVu/bTtJQNpd9r497VY7dFPqNtzLzAf2wVJwnXG5rePy
aBZlW6+02fL991CX3gK8Lp58lcplOYrJxB8+dJxZZdm64TAsJFfwnF9hccW8Gvfp
4GpBy8a9pDhcwquhobLUwQcSQuW+qDPOno2qVAKu8GCqKfhHzhGeQjAtbv4iJ9/w
hMCuInkVcB1KYRytH7Itupjbf1lp2/xyXqub6L7YqPHFgjy1aibEYh4W/5xGwbIS
MEH+d7Uz1pU1OjbXvKYSmW94cT0h4IjHmfGdDYOg31txFomrv7QYkRw2J0U5QMhp
LcZRW0vUlFI+X5/vL9wR6svMbzd2A4heOEB8782M25rI47EHc3hqzzdB3fLUqm81
mNeeVxR5yGdqqUknP82/3KN0ymZXk7E+XUpc0O+Z2NSSls4a+RPHdO4ljh2ftt02
dVJ75OmBlVrsyqONpvkob5yv3g3c0ojClipVsdCCvUpx8XXmR3ghW0jg1xFAHX2s
lz5mHvrlpS2jGOD4NnLHm6DCOQ9447gklRqJVJBwwlOGsMssTIZDlEtKWELv6dNd
uxdf0CxApMsDfZO+W/QCacmo6RsFLflNDUWpzG9cQyCt4kmNGaFQqBxkQfGGI9dZ
WTfb8QPHShRs5NwFVaT3kyRDc/pAobS8gTyTKNU/hSWUZVwJPj3BoYpGX2/m/9LL
KsVdsrlc6tsLVGj0lz3cj6olDwTTjDkGsTUmc10dpIRLBnpZmKPIM/Vw2Y3JxRCr
lkhEgpPGfwgc3fpj8ym1f21u/DhTUWSDkhisL4J9beSnY8rUvyeLrcn72dFJdk6k
XS6gPjPGFdGIltYvG43Ut/dzGD5kKEiQsvffQq3jSyiflbCgonZuZi0nNsHFrBqZ
DQXFKpdVofZB6yKJURImSGgJfa1F1wi/F+5K89UjC0DIHTeov1nSqZEo1RkqDygy
0t4TLMZEzc25100jmwArrp0gA1k01gVGCKOnorPGs/NSoshQlMNM95K85urFlyoD
nfRuHhDrTmS7luXWst+d+jjvtF0HEMhrhCgt2u3YgTxuTxL98+L3ySTrkX8WF88S
bcfVvQ2NKpMJMxQnfoRgcHGwSuq2FUo6iVFEcHWslBRHBBNmqUwU27/Gw6A0xH4B
+VV95DTRPta2M1hzGui6AR04hsvE9khlehAMJCymjzOr1wW6ZSTUHf1p3wMEhfcC
nzKQIz3v7pkVCZmPuHTIJQ2bRunRMBenahduE9Rki6n6gS1gnXK/dpKSA82Paze+
08LyOme2pKXSKRDKgMpqFV2dgXY0Mo1NXzOGkSAhWnXg4hitiyle9DKKYuJwyJZU
/dPt9q4vGhoT6HU0hxnmF50S8iKAdXm2h1UEVScabUEmurbMPJZjlpQfLciy6sWG
dA3wl527+srZxOf9vL/ZHEPflIt+E/UKsPwAkW4FxMPXpgnXz32CAyFguxayW3vG
gj8aHa6zw5wel4+qEKoe58Prwd6fXYpRH81LGH0qKG5gAugHyRNlujfL4AThr458
AzfFLMJwZd/OU94cv65vMtnwRlkfWFf3Z8QV4iL4/SEWIwmVV6Ye6ibHpd9FcFxX
+CmigscpGGhfVaxPOWGRlbDanQtTE1PwlfrLADMqpZXSqrsmrLv13X2FT9b85wjh
ZuvVk+VVmGpgNoup63IHo/YmPS6Q/o0o5/sSsLRpPC8+iAVc9umilm4qRtdIygmH
jed8XyzHSrq2VPtstg0BoDw8DmwLY/qhNFXjNO/16/KINYwAqwrctVMLBF2LL+fY
d6vf/6N/WzW38EUBN8N6m76zAyUDDYBpjX8tsOZPLjLsK14AxBoPRVJzLOQmbUkO
rsNEGlJUOaL6ojDPy94VGLmQ0eZdRIU7WBx0UKTECMSVUeWo+oXikyPXFB2xrFO6
N2DKqcFKqYpbgUd9CwjXqf77ID8fml4ZrYlV/Bh1FtX1MWgapCNoZCkO/Z12KxaW
a4WxR2In7x9TYwLDUV5RnYe2iuJ9JWc4hZmmzwfcwcn/Qyl+QtcLlG6vUYTGCnfB
TCPOKgesGRafd1u4+srSDQsNRLasVwh7+Dq5AUwsME42fePC/yU7DIxAXCWuOojq
edMLFIjhhDkBaoc11mp4b/U1O3ePJ7YXAON5HfWDdNobZYG8WVeaMPHCleNr2D0K
ug3ufnjd2zGunjY45+Oa4oSbtKCR2wrCq2Y5KbnQhWOC2bG2xisyp6fafYTZVOzo
QIanbCdujjwKxtJ/54ueoZTS7ZJzxSj2w+uPBztGjtYfhz3bJkcRC1W69HO5jxdv
s/NEakDTY6IJP45xvRlsDg1cB034vJE9C7AMqECkFGic2r9wtYzMntnwK0CghFGJ
oeKQH1PWTtX6tp7xzmeYfpI1rZCtkuZW8VKTDQmN4Qct7AUAk1SH+z52PDFb1n5+
3PBJTuO1/bzJJI93+lVa4PTUhLmeM2MhoA9LDEppATRqf02pqnxCeWm6vU9PeIth
fhBnsh4FBlG5wXNIeBW2UPQdUxH4slXq5SBhxcpj5o0DekiGlJbzLDDv1xRV+dlE
Uih/FPE4CxWWwBtc2C8TuP+HqtnhhbHz0GDuLiuFqoWLfgLThGY4Ig/EZ7aw/niQ
dc1SBrm3zR3wOVVi6t9PrNA9paoRBAqlbZkKmQM1Xzz3bN728T0+CA7NrdTNOW/u
gB6cyRv23/ltYhd0S8JONOhuOLYyQ1gadZQ7MkdSkH9lXxGGrXvsW6U3JVnh1TAD
6Ul4HVef1WtrZFGQXZxgbST9eG46zYRXtAt4ohZbBOD/0TYCVdFf9xL7dsejkzfq
1VjTY8JQDcWJ/CtgKP/bzr82EQh3C+nPcXUZuxxz924Uwhah84rLUMjKDH0eDZ0T
HNBlvOg/vhZL0bZWLKI5Fwm5+WpbEAOINjAolpzP3ZJhNiMoJ2XRD2r/68PqHYev
yqZJnJhOqj5t4ZLF90bKUE9coi86tNg1mWEpNZ1Fxb4AGQDLEIdsQymOjaXRirMV
DLwAmBQFRjV/R2d6wLC2w59TGgfbuxsbruHodEsTOZc1SSkz1ueNDXG4bK8K/NR+
kDOoG5WZPuYDrEWAunk6rRYrjQrvpP1JhlOimQyUbNfiPh3BnhgvVSCxepLrdspY
PMcPfFOordH93yK9yNIXlNAKfRgOrL3DpphgClaQYjBe8GJco/4YML/Yn1Mz39I4
/AHvZTpClEGMoH4krYBSwtN2HMBNq4bRhpuPakcpOMeptgByuV51L4VhuwpFzl1q
j+33uWTU1SMbhjHtLFgbgpruXMC6YJEy4fOD/0E+N+SbMLypIMcSWSfHVRfjB79H
gkMCdoPL+AV4qHoVl+ju/Su5LI6yLmA7BoDbEFypc/BinyipdPjE/J3+eahb7g/q
WgMs0UbVZ1VisrGnQbE3uwHlQPj5XjOOuG0R+Q60zkAxhqhC76BHLTrb+PhldBDE
IEXkxJpU08rhUslUU9c00Eon4ioRTfK12XSdqFRp9wi2KyC9VxkYfyU/Lz8sMpb1
gmCF/dYx4Q08bORzAY9zB94VnRGksj7Cf7z041cwj6fHn0cszTxBi2p09C47u7oC
TWvHtMqZRvM7LwFy5amIoY0rRpZ1+1CZ1b9+tsP0MDQCLrKGw5QsIA58AqVDQ68c
BqISzNpitk1BQLdj2VPTdNKBgcDRoH5wG35li+EFG+6oT//w98Ls+6KE3+FGuu8x
d0/l3KUcTI4ifV/tuVl3pEkKWwpPMYkHNI6P1uSBN5oNWORDfbVSI63RM/NSe6EQ
XeHrqsjrlWADREayc+b3CRiiIko5v5BE0hnWhokFxYQ+ZdTXBfxmlICz17HsJyVC
/8EOerq3A41NKHue+WCpA9vsLnllKo423nGfbjmKK2iAZbTwiMuUA374z+J7M3pC
pEzMej+wbP7bb4lI6eRXHjqvrMoloG6nsIRSwX0/hIgf6D3dMAiMYMG/rDJQSeAu
MOEETyOHUZvAGCZVp2oWdO+gU6LQ/jMDP3uGz66DSeES8zOZ+0NA19/vVw8Nj27u
BUPaf76PiNJunStrKSaO3F48gXe+Ggje4ceTTEKcnzUIDQS1NG/iIah4xEipb/N9
H6OFE6jknka+XSbIdpoGoc4aAT+vel18bNMsQ94a0gorOh6yMaSUFSehOClU5zlc
RKrsCuWuPZT4IH5Yq3aIA0tnrcV50K3w/mJHjdT0WeTatbi6JVpMuXF7NKEQ2zE9
E5S7qclmuEF1jWSyCLA/Led8p4j7Saat+M71UZIFzvWFnLqSQYUg9elUVhxZhK8v
Q4JmINohjnkm/SfcGmskUZFpmtkGxJoJaRCSAYJwZzzUldrt3zNH0eYDak3DtRHs
HSyFQcvtMRBeu1jDVWAmH1KE+FajmC3N1Ak8JC3dOsPtrTwhdiIBkfBgIJcV2Jmv
mLsRXYDlGU5IExUlJ6lTAkcGPOLhsHcwqrVEeOcTvvdtPq8P05xG1RwPQG+iJ2V8
MKIxhJ6oiT2vh0gh/vlyYSyJqY3BFtJxD4X7QA91/GEKTQfY57T5U+lEulEuyJyR
VvzNTkrQ2+Y2kjDOIh9Z/k0njWT0CjkXtExAclt5geSmDaL/HEtnYn0BHTwLA8Fm
k+UKRYSMD3CjB2VJwGuooUo3aINvUkxswOzmpORnTNnHI48gkI6NShG4HoU4oCNw
ujncKrLXB2eA0WXZYx/T0OvUFN1ZtOOc832mDQeSJBZGEuP9QW9jO731P692AA+6
5xjR/ygVVLjsuLE3Xuggbs02iEKrdsFcemqYoedimPYK5FguJcwR3qJLwShdfXbk
n7petsoqJBcD+O6/7fbjP7h9KcljQXTN+69IvCvC3b2ctTc8iJz0G+jhQ/Re6D+q
ctlJnNBvgOhkqmowqCLb8gsplp1/M6Q7JrzlnnKMsGMbl6qTVfQKKe38KdpRHuMW
jduxK8svmuRP0XyefPUY0k0UgPBrBdwLXbOV8/Juwj2WOCAaKVMwNaAT+uUJiQP1
KUsu/t6UBBmCEvmMvMDlcoJ3LXI9AK3eMN/eGFsoO0cAu6vBGaSvgt8lgtL8rcR0
Dl8ya8/2/uOGM3DX95/3TDmsKBRMqWOI5iGTfkrLN2EfQUs0YvkFcUvSquvy4Gpe
F/5y316tHP/7mfFeXsuNW3eIhc14V0Csyviex1XaB3n9ZR3uRgOT2aI8BlWaQ7/l
cBQQzWeWLsItZQa8KYa0w7YV4jipcdpC/nNXR4GAdJCy+apAjda7ZzEXGKfhzuPf
DniunLqRWyASywUPM/klm+Ra527wc/4a0y5OsPl6hBdZqPpmr1TYYGlcIG0X4pw/
V0M7n1Ffr3+k31sjppY3diHMvGbVkd1eLUTrat2M6E6mLnua54tOvOBJcwQXxRih
VlinZf+bo7Q2oIpxEvPcoFP5JfTEfM70IIyHmlnUX8KJ0lf8zokWKrCGMbOBHTpa
79Gxzs4tFg6hx3IpL7ENaEyui3GsLNtjHJy0aVaNMYy2Ag+pJTqMmjuXpxYy+Agz
QiUKyndhlSK/sLgfmRGIkPwvv/6WCq/blNi9tqaIwiVErrKwYDmKfosW8lwh/PQg
wq8OkyXUQCms2XXa04BnNqroZ0zsaC6lvUrmN11tmm6OFmh6iC17NhQspMMCPin5
oJRJNpj4T3/aWebzhYCx5Boze9ExMnFKZJP7x4E2b49X2MuMmsGyjJY7T5iTZcpN
Y8y/H0vwsxWosLGDjV1rVKDoYVHJAfQWR+53EZViqXbZLEzvyc8bkH58IpDPkzsp
MPEss2z5JKIaJWQn6jF6vov9pWA8UJ8t4Ee/xQLOs0lxRJ/qKuV1ClGHWg0wjn1N
ZgXR6FgAMAQ9gJg+YMphx4Nr+n5cdK7PcsaD2FJwemkL24MInWuFgAAl+mPA9lgc
PfxZFvpVyNh+JZX3Tj+KLWoDOf3ZcZVuFzOhUFY+rssGtx1MIMeXIfPohT/nYQaA
9MvzTQTYSOYymPoGVOe0eBFqIsrnL5HF8YxLmUglq5KmBEwdFxPpl+ECYMqyUy4U
hp45IzueAjxAVw/O/sYTbs+nH9W/YU0jyFLIWSjd0mVWhVCm3yh3zXug8SxS1rtp
zICaWu227YBdn8Tw/ZzBx5U7ymJf+SrH2gWWWYEenyHuM2UHULPHkhHj+t95APuL
zbJIV3BFH8cS3edi3t2gYXQfRlyFKQZOf8Np4+nkISu5ZJzQNi5fLcLUIm7kYxZQ
5db07QSW4FNW4uxKYVWPFgAz8h0oRuV1IZvZJ9nfQOTLrAZbIGUKmrjGd9h1euS8
LjpM61noBszdcfC53Fa8RgXAoRaasBOmg571/mPpiZAbjPgT322I5TKTBPYHP1OR
yCEBkWxicy6oJBTKnyWPgETS59CkysK7yMmL5snJZXYYmzitJyRfzUC7XK6/eu4M
IXoId67fvr1by7GofDTtbXuLTylbZS0ssR/qnT4p5v/BQG9M0+TYbLJ8fEEuzYbw
gdmAc4DzUzYvHOKIYngVU5GQAkaPQ/cXRE0nO0nD2JFYDCi4X6F8WtzMcyrZymor
CSt/2gGo4cikHuUDzrhY2oL2UqlDSGkGijrsJjckbWqOMS+YhVGA3w1HVqlDsmck
KTyMNuISx3XmmSr7wU0bhCVxXwbI6/j9HbRAWA+WKQB+LG5tXekfMABqiXFpjSbN
COfnz22sJBVr2rMRycywELFn07uOoclBgm04uY/ZqkTZGOaRSGWO2QMG7DrZx6jm
6TUJSmN6alXetUhGXEdRGZ10yYrcNN/Z3sO4U3vxMCElHEqfHj9Z53G0rJui1l0y
3CDpLZCGGrEcC2vixgCCKIyHOrF5W3ZAeUNNv5uRlAe+3KkYMSR4x8Tz5UlKB6B1
KWpKsVYMdU0ciqWEIn5FlM7AVzGIMwGY5MgUDTVe1dKTwqPiEQhNNhTon55L4UHP
OLVilN5MvmFnWNJVn02fLD0wHogDNER8KUlXPIYKcbiH3AenG3phlzS9FXayUJfr
rAyR1ZSDdIueje7NlWiUTbO14gY28hG1F3bYH13rs9KyHi0AHePNUMmpHVAhliP0
4dj+lIA9mbNWl1YsQLFkArRRmMyI/2HwzJER7DmHt1imzlFLy01cieH7wVIa5vrQ
3mFwjJbOPzhkFRi95TomKAd7kvT3QlN/Mi7Tyf9sYKH0wTihwpAjLmUcnDRlkAOm
G6CSnyPjZVwo0SxvJGsXyEmrc5SG6bJIhfFudPOxTiMkC8EwyRsDIydLKDghUsk5
ZYXhP01iGpz7gF69BJlZwzitSkQqVfXMNwEUq0NouUJhnj1m4vQ+h8FaNY6NEltZ
vSOiMpR95dprj/eq+woPcF3ZiCSHEYMi3+tcYO6UC5z9sOcN2xJnhwgJA6rcaz1E
EUSO36AzJqdxnKsUI/nK8Nno00YDSjJEl4MRCPuiHCguWT1f/LKDfP3wDao2dBVq
clyR7zVEvbBxaeymFr0/30ECgJ3k8H4Ac25Z0y6PC7etOpK1uG0/LRkOIJ42rB//
G3iyhg9eM9BECio+Xz+ACx/wIZvL7lF0COt8u+9wQ15t03IHHNa2lP2uwyccYqmv
oO5uMsdOcIf/E+BvsTDGVqJSpCbvBAANfS+KAiQn55qObRXpdyGh3JcpizwV0qrR
b+Wn2fn759CBp8yHeqeCnpJMSMlpOyn1zNYzjbhQUrjZub6GUku/hDY1NSP0M6or
80K2qR8YA4XOfk91IsUBvC8t4m83uJZSznauR0nWHMcSLdHVjHgQpiLVKtPxsnWz
rJNu8f73spZdtWJyXvpE9eOTN5gzS/9DG3o935dUq/vlSW3x2XdDUrDW1yFN4dLR
xeYx4TWHt2Qx5RWUzgwb0GguxYuRy6nmMs8svdyOKIS0XU9+eWKMZ0N/IOnT0eav
reWFvo8lIZr9WHFBlUnXt0xN9Z2g7CzvbPttycnBc07qeZHO3SZhE+5NQfXR8YDn
2ovmr/8gr/U2ZbfRaB5LFVcN9QwNcC79SsDDZF49TcECyCZ3obqAZ/i1WqUL3Grl
6VxGcmzNCTI5jOnszxzbI1AjPBnblcdGd/7IQqDoKmKbxe5yFKJnpa5Z1AdjlfiL
7LAzvC5fkLFw6nQ6+MlrdH8xV2IYDxvodeweztThuZNxzCo/GiOQWyd70LlTh/mZ
nB2HUpkZ12QObdvm8IYbRSeBnPvfF/OPBMF3QcYOqkA9g3vvFGQo+BPKoZh9PIlc
ybMd6a3qmvubCS9Bz1Qn9/1qfHj2/0mYziN8T+3EGKhKrLBqh76fgPonng/RXfvm
e0Yc9+kahgem/w0Cpc2Jcph4ZYJETpbQSDY813xWh0vmnCGjl57JUvm4jBtfJdrd
HczlpdE4j4Ph0FFSoNRmkTTE296IRWQEBjCaUfBkDNqc1QSiRItrCRh0BlisH4Qa
UbMsTCmLrc1oIQCK/wyrZx/PjYvsicqd98A9BLqOa1p+E/uqdjm3cXlVyXKVoWy0
bd0/9sZE849e77YOOF8kMxA04ngHGV1bZM+Qb18HaV3bAPPR1OPlA0okCzIK3Sdk
7tIHWRqAD0JILhcXNQ/RJK+mOwOSII7pLImx55HzPCySdOllsUPqpav3XTkj2jk9
D/XlOr0Am/lAnkU210j2lYUAKQkbJCk4J3NWRuoJaVLsZLVCTzMGkp2mqx1EuzZW
JQz9LKMSR9A8StFY+PqGMRKnPGdTthIoAiDgoBfOSn4uTHJnCXwl8efAq6dN1hPJ
83mdIVGH1t/podMv/X7/3YBoVNY5VbXtYjp/NXo9aH9yGj3W/kYWGCX5QefXaDcU
/aL3u3eTyR+1z2/MGZ10iVv0qc8JJB4NlOfJRKuFaP7xCbvIwFvOiGmBzrjOwIRc
asMn65kIC/Z5z7FVJqUbASwmSzY9dObmCyRrGn4Yj7HAeyYDnMFFpd1RzS33n/M6
QO4Ww6Ehk/sJHjTwqzD0+tWRZu26LnreG1ZyWAMywKnqhWs8ktxOT6XCjKXOVuyL
NcYlnGaMO9ynhSP7RNznGIFLlhVVkxnl891UaKKI1fvMPTdblB9RHEinKVQZDrYc
ld5tpsnqmMJXEhhP2bbmyruStf+BYnvE5a8Tsfrl5baxH5uKprudi268yTp/VPKb
BY/08BHybgMFi+e6LS/rVSIARbxTBJm8RmS/x6Bl1eD8+uniuyvC4rgEbjRPIbuo
pYkZSLzFG8IFzk6CI9FyAc1rl/lnhIGS8caj4Oe85RkQcDEzsY4uEJgK0EpntNUY
NtCjfFxsfrOGj1xXlRkILYaRu5Z+HDS9C5AH9C2sLzTipRHsgOeC6Xf+Sxr4sjxZ
+PSi6rQHVlZYlaheFIWIzYdhspzgZk7gJ4h2HIxasQT7VCwahByUjo5KKmYanykQ
tKjx2d2MvLInzVXfDkuyqyA0PllG5uUxa2J0s8vC2qioy0ZAseHcT6/5V8iAebQ8
wZ8SuNBQY8ONk/LUwOwo9s1A8fiYeoVL9VCrRDACsrAtMN1wWhDxCD8cRF7+IWVC
zLsxQPYDAEqWFPoupuH1cxOt1YxS6u0pvLxlwdXbWR7akKPGOWw9NE+AWMrx7Euh
iNiDbp9eP/8fSA5RpdavkyRnGW/D8087uHsvYVXnFtTONdoX5Sxw4XMn8DBX0/LD
8qFz53sJ8dwCxzxWuLK4jIqs8+B9rWOlUqtRoK7v0UpprlZiXtcZPC3KKTNhYSZV
FLSSS++uH5S06bbl89yWzit0OvsNtbd/R0U4V6N4Cxxb520uNTZSoBdVg4zX3+24
PRHW/8NX5by/mXeF0SOEUUDxDH2yEw7Fl/hNuv85GLBvLL0VQkpy9Mva8LW/wmRf
LCBQ7xS3dZrfeUpY+Qgm1OogFKdY9zVj28N0osc0xSB7h+kw/354IGF0IfVg1nb+
ZGmL6KWYg+R0eBYj78MHIpMD8ymNF9W2n7x6qanMv23+I600ZKmMH9Ifgnj57Cns
b7JOz4iepNvjjCLKVaO4qUtOe2Bg7hd+EgJhJOxENpdQFvx/dD6dQkdxLR02QaDX
5LcY+Q+nZ0gjEXOwvfQIp+gYypnTWGsTliUA812e/1rinQMQ5/PRcMm1LMaU7DX7
EJE1M7lW0rSs/NBOCJ0/hzhUHn0hG70gyLfyhLNbYnr6EnHlFBmQnXsnkMZJQoEH
/OkdTXKyiNIj/iNHSO1Mh6KnTQCNCvzC+oWKfCC+4pFlEw9ZspltOt9Q5r4/KOe/
po4aQm+xhzIZ9mBeZ9PITJjk/fccq08RJx503ncE1UiPsCucTzM/KE/pY+39gWg4
yg8ymXw0hnF/7MfY3RL4XJsXV7hD4YNbQhHt7FGLl4OTk69+3jQK0VFHSc+Ps54D
9Xq6ex48yuf4qwZ//4b0YF2Ywa8wj597pcgG/S54tiw52njQpnLonhh/8+ovgEzI
Kh8l0C3f2vUDMSffHNvrB3txs0C46phoe36wzvpyIpKI1AnnX7Sy5SJUtAcx9DWK
q0U1QkCdm3odWHMFZHZxduyuiTxwEo7XGjPGRpEWhDS2IZ/rBnnOoaS3kA/v3JzR
DzkoeisjFGtKpkBRoJB/L8BkHi8UVWbVKI2dH5xwdAFu8i6Gus1cB9pfYG6c7kFT
SpyZoQBk5q1Yt9+yHq72kT19pdX0QmOiDXTYBZlfmoZq7cNic0Obq0gSiPB3p9ts
Iv+Xdaz9w31oy+2LXHZryA+Hu92j6R6xXC2aw+SaqELbKONbwmWJuIFATT51iF7h
8LQFMEWFsx54rQr55xwVlX+gzyNQG4rV/tbRxM549OaFUJSTkCSYnhMzsNaE7swg
VkLOXa4Z90sJrKDv1JBfuHauvQbVjY8xr3LER0wypeuhbgQTGUs9kO2i/JgQorE6
T7MT53zY1x+wcfRVnt4l4H/7l23mQSov8g9Tub0DagFbYTzLPf3z3amtBfjl7RCp
LLQ2qeYQ8IBC6xWxSGKb4z24kBtGTDQBJaifoBu44AmuEJXRYii62uNt+a9Fej3m
Cx49qU3Kq3FkkwiwArY7QbAFG3tTGfHk+LZO7t+NN70+tqqRfn0ioT20KhTWZa25
deQg8xUGHYXkVU/fjEVeHtgHlZN709sft0Pe2k/fNxT+qBKkd+J2G4fci+4WYLv2
9HYifhuEmex+GeNl6U5BbXB4HShPRDSSgXWD4tT/q2RS8XxM33DTXSP5stggAKAO
Mn0ZYA3j6vmYm1Bphva+XOM/iRZ6+q+PLqwds1hwTsLNTgnZNJlpvPlDq7E8CEs/
WGbbY2mUhjRHtuBcqZwzuZTlGyvVkFCp6NKCKC/dJD5trPuHbVxtf2VxIwYhs6mT
UY8bR9uSZjcop1s9ScQ9HrmR0KETpVwAuln0iQGx9LpQFcw9wFTsjE2k5KlWzJe/
jgDYK0neF4KH3dfTM04HQY4lySb3kZogKzz/bjvuVawE3rSkpucCL/GtDuatvmhf
5ZtSnpphqOc3UOy32SwIRKgExzqo0B1WX7gD8voisC+wASPB3TaWPh3+yHmzzvS8
oBuSnEpuBpecCUSrROLPLjY1m99aMIehj1fmR8XneUXDebQpaPnp65iHrwVfyeQw
mlGqYpCfML1nYRO+wrkk1H7DHNSVAjJNl2w2Cv9yOe/E8l8inVZc/IStnp43U+ra
H8Tom0U6iSJduFNiVQW9dKwF0kVlYroyObJx3EFcAo7pI2/vKB7CVyZv8C5E3kvS
cc6638GLCqxGCULS4FQXRc4f6kMOO7Cvi40e3fzm9lLSYUj6Fw19asgEmH735P7d
Ekvmkaip8GFWBoYi4SjHfVGdoCjXyLrzOhZh5kZU2UrqTC6YfqsMLVNj/Jp6qzRq
1j8E8TA52xeMrRhIuSu8IFtAPtXeUczKEaf2sdufN4eOmmth5ZLFm+HBPXGtsnJ/
hcIquOmH84mBVxhyWJKTB0kAhLJJ45dL6KubJIxAS9ufCCqRqOBPrp3b4vERwOak
azXGzy98DLEtwKhF0IgHUZUpqBczbLbsim4Bybb97WN24Y4Z9Ubp0vxc/GVTXFqw
5BjMikJ3ISxUp6Wg4IIh/hMsgx3vRd4JGIIQAjtb5UQ8bbv4qR044roMIb7qBL/K
MPIRxMlaNCNMaevR9uu/U0vsva2D9usfEjVjXUtM1WTMnf9qxZwGdppd76Xy/zUx
1WzmsMiakhE4hdvDDZGS9IPqxv5ygv2fwpF34qH+QPHFxySZX5YueHg1T8mUun4Y
AhDd3UC25od8aI/3P1+SrwyUl5Vs+P3JCXQntc6QV23swcE6yiMNYo50+z8J2kLH
snMrkie6rhD9cKsfEvTpVOa9LUb1Pwp39WYkjWORs8nErVFLvXiN3wD++wSm0wBb
aM4ygXW3os9+WZ35oJE9xlbT45yjXDSVHWeZW+PLVdFWIrkzOz1ftQ1OykWtsMb5
wNl0Q3Y/2TgpMWiSljKYeVarZsaj4GG3AWWN1hFUSCIDSxRbUbj8egZntg+YlrI4
8jfzGenltJB+sA4QHdIS5Kt7nRHj3OFj76uJgvfXVAXIQXJZkEicICGP2M09Ww7N
byJK/viQDfgT3Io0Po1/5k/pnvB9+m+5gy5nO477MGt8682vC9Q6AKA88xJxwG+f
xr044BFShVb9AQhsmEg58kXeb9bQSndNzqZfJs4SLX01qGSjHSoePLgQoQjADwoz
iy3Uv/CO/hkQYq5hgVqroF1ZBhBQRyZwWXD4dA0HRj2xw9M3fr8ssPa2O/vsEiPa
VLNw3NF0Ut4lxTEEgnXZuIQ+IQBaOSqey89MNG6kzRwg5skmZO6SCY35t8uCsj/Q
o4GWAK03SgWcyV4vu/QiIVJbSfdQjPhS6eqbD2mKOesAMvB9glAq9BUtu7zycHFQ
jvq2cwP+f8gNBek6wQIdMiRtp1FyvGfkEJ4WriNtvLkcZDHAk58X79Sh5WN3xPqd
ItPuEKljnmR0FBE7AkB4LpDVMVKy8IOBmWsHUEHGxfuLtDbn3k762Un8YxpP2tWC
1SyrJq5fyrIX5FgM//lKNc6RKaIS0Lzz9DdMft8sxEk5n7vZxN/PG7Npkp7+429d
GOydK9wBac3kjcEuqBtRr0BYDc37EA2CxID6ndgJ8kFVHrv3zECzeRQ7j+pgUTCo
lCofLfdaybA6BdUAW7PbwI5G2dluM2eIndVXvnE8I47YJl8RnnAJVJoub5WMxT0+
t9w46tNElA/Tio0AaXwYPqB02yzYmlYLmYYXXm3WjSCdm+1MTh5K2I96z5EIC5sh
GhBQrLFNuBdnOc8mt/esKql+s33PtI9Z36O5yJ9Wzrnot/zlJWBQgIaZq29n6W5G
j4LnAiY8YeZU+rgqZ9kB7YXD1GlTQumJsEIdKTNDNFpvaU1q91LMcG39lGvydRE1
oR1bVsyONzryeaFtYu5i4pOi657w+KThZQ3XNUFkYNC8J7c0e9Z4VJYp94bR+hWU
9Dj7vdXKbwixpDuy1CyUzgD3x4imse2no7fmakTA2W9w/V8iZV5/cq0p/2UeCt60
U5f33lKm9c9Y4OXWGgVray/S71M4lhRPGaqvoNcCjiJ9mw+E/qrnAbm7OtC6PXLJ
Q9N+s51ACw03IE9UKhG49eGPS4D++ISqxzJ2XnNuh4Q/Rn9OFaqwf7iNEsYC7W1L
/EMss2WOo5JumTNdDtKH+CbvNEOmqjrxXhfLV0jz7uSoGXhWT7eHa30xgz71TS6N
F2eVBtLogYGx/qp6qg4BFsHrO/aB7V+4mctuufufmV6r7iUC86XUx6YA3Kw0+2AN
uaVk9wRJYVstw068GRAuJM2KQkyFiseT7OBnn04jXbbr3mF74ux/GSoglMVnWW8E
E2Ao9l4ym/RBDwBiJP1Kj0tKR7B3F3YL39b1n14pDcZF3ee7b+OBXPdHa6UHcqHA
GY5D1Y7BT2XQ2PVLBRXXsTV+vn9QMhwFhYiRZPDwNTAh+LkZW8xT8ISdXPvaAqoF
cgP8sTuggNxCI3nulcRX3VbBodJB86CD+obJ6//XE5+bqtKXwiqqAzuz2c9aX+Bp
LeHU6bQN1cFUR8sqljiYpT6a2qlqYmLiR17whLrbnFdYpU1FVf8uscjW463T3sD0
p1SyKH3IYOIGpXIrGuBQQ+PaSWjCBVqgzmzJu6f+yNjaVerM837p+hzKz40n1LLv
zxOK9evh9d1kqwKDMJ35oV8qzMeourggl2A3ERPuBObBoKlrrNHI2FGmmDJCZZy6
w9+Cz5TdV6SyM2axCjqLd70wtcs7Bhi4fr95YNL5kXE0cQ5P8sooceqGjiiiqDLB
blGke9FDvzXQjyJ/azFwkHEYNqi1usT2GMSKxxtpBu2E4OA4Ag4DyJnunGMAlqY6
5pF3AXwFarZhfkq7Vv3HhufnmGIZSHZTbxe9CLyNgBqECePTGg57enLBD3bu8upg
jJTXwKNfwHaPhQSS68STW5ikIYXP28wCOQ9vcmgHIpvIm0XJCa3/A0pA5h5BUr73
HQf4Pz1kdHpGoP9N3eg3pXwVhYXO4cBOH96bODE/+DS8VVYJG2BmEa/Po+XttaLf
8j/oGZ7weYRazK1fWECnjCAhlfwS6nBATVpQv1phBttWPvVwioVhurHrjXIS3NeM
UXwK6i4guZ+iA2Waix270noW0R6VKYS/CBxLK440YwvXSEDio3m9d2wFWkRZbLWJ
WGgJDuRXrHTwXazVV6mJaKng/NT/QxWeWoynBCtfMZok3GAD2z5ywuilOSXPXRnq
iVfGZ1iUyTaEwSt4nblwi/viRwT7GRz6iH45dMLEKXtQ+NYtKZDc5RcuG9OpbDt2
rDAjhjvReHoJaUkAzmzcaUAxPlsXxeOiev8S0JkT4yep0Yk0uL6qJhrVCAhw4t1C
T6VjuMwOynJIfyGqW0HLLr5Ey7RA1kUKX7YLNvVA8xlaMl/O+hRCQiN2tSsgHR/5
OPzroa1IK22tFkiVVQa5WItBHzwpnF8iym6UHdVdMSLM7cfE1bFk6YbNgBQDoGOf
3KK0qI8HHqNoXhTDCGsK9Splxq3sjIR/o+O+QuKrFJ8RdJNISk8ZGbQbfe+crrrK
9syzM3G4lMuqohb0Ii26GlOOSid6UfUZQmtAtmiX9s4gTwl8rUHL+hcffnoJzEXi
bVUxCaEWC4NnEHRuKSBaskCmfnXGTaje8vryqJi/BkafxPpHcUqcrolxbRKSaYfR
BBGNcjPzNJVnq8qE0057Vm+eWaOVZ0qmfFkrAYsIfUpmX90vxzw7ZJJ0jt8wpuDY
E1W6Y/qX/4GLOr1WjDL6wFqDIFnmHrT94ALiHNgaj7u5VJ+2bODed/wViR6UDUD3
29Sw9Xd3rY4cWZcjYbm6CJuBo/VvuJVfV8IMnF6MdH4YucEwh8LRDa6LpYHLaWY1
4Jdv7gNxQaZK6qGSvrTqqWB39GMbBKAbQIb0AvHNCgDsyeRZ+hD9bL0n71Sc0mug
+Bxu3xT+/7uh9SxRCwjZIjvF2F9110n0IaIlCttdX7uAveXwC6RrQYjTvNfZwwhv
YKfieK5JCGbf4ITi+y63LsJMlbMi0rrUiFmid4JzdRMxJruAFVDSJymMmGf/dL4p
jHqo0lDvdVJ7zTZ2JQcvxqru4v+wUsyAPxKqgAwLnJ1YcOqKz8fpGfdcouQigj0B
IxxtbgkyKqUnaH9cljInzpeIO9k/g3M55YhrHZNaIaXuneV6oWhFE5zhkXVeuT8L
cusn2vokh1noyHY7LRFPVinTocJqALigdsk08v+6VXe6c3iWUOXR97eGmRQ167iG
CL/Wq5tl1rM4liyf63MiTt2cXb7bFKQwGKkdhtvmP7+ro64HiPl7ACWBhP54eAmi
UluI5f6fKZrxbtWNENHiaAG4UV1WsLEXmPfLpmdv/TM/b2Ioo4nxe1SHWateTcsA
QvCpTUtCCR72f0ZlIOS9eKb4VMYoeeyXNlSUP+iuQ2ackDAqn1Y6gcS3NucKRBzP
kTQ9em/s42HHHfrBhmphmlqFc/JJPr/sD2kEqet60bL8VERpOSqeX9km0fg3Ze4i
EdWl3V8HGGbElKBY5ztaMdiLKGDF5ZXFh/F43b9A97m0vwCmfl637I6nx/uWJN92
teXIdqEAQmF/fjuQiOeWw/jA3/ZtHGSxPK5i+FCQv2hRwN0CVNxJGmdZ6SUT8bF0
zEv4KiNr9+/2eqlYlgeNYIDPGMH+33JWldvHOHj7ENNqlfICTeRNpMYAYd4ddBPF
HFz0LjB1xJQJBTPPhM2eZF0F4EQyBUtalrrU1cmnGHBa2xGj3zkrxGdig7lRHvSZ
0IJpVALkZq9I8mjQnWvWZ6SUB6nuxaT2dzr+yK/8cQTCZbBmgi7UTLPtBO+kZ8nD
t8jj2Dwig/uHZWheMgK21zz75pb+3PsPP7eN1yTR7GrtIdJKaIYOHEKTRGP53MZ2
EbK1VHMAcewHn1/UxRPnjbBH3AAkFZUQ+8HjnOnufTieN0e1cW3zA005q6htwKHG
6M4yMcxk9uAJVRDRkw8yw7oBcTxdLz/0OPFGkcObYsOJpzlBmt3BLnMgGKCZzgUD
owrtjnJ7SXJTX95wi33fClLx1u80ahjLQui8T6EbyXclxZe7/mu5F95lq5hl+qPY
5+RWuvEk85s5xotju/j1u6BhHvJOc8N88tYNM2aEOX9uxl7itoQ2p5HeJ/cd4pux
oeQTbxB2jhCXXoVxTcpCODawV3nBiPTkOkVNgGqex0jkPTOLgvqcr/7dTbywpqaf
nKm2ScrsHk+++iQa8w9KDYNeMvLKt7meItd7zjK5bk9YQv2I9gb6lKoro6MK74Dn
sZeOOaVNqF21cA1g+BZGzK2SloNfsIr1GhajB5Pbbt5TK0lY6KM4z79+vnRNmF4T
a1vkvB/7NadGBf8yB+JWK5NwD2w0ubLR1PoYJpbl15GyDNJbzy3vjGICEpNQz7c9
Z1zVuqE4kYm5pFB3D6+FDDH8pbn9pv72Q0cG54ft8IqZegZFuIeVNbN55Dlb4MT/
6MX+XfMEdFbHXWH0lBB1duQN9neoxrvg9Hv+JLkhjTremhWCPtUR44VVqM8vbRnz
Ou2fSzQdMf70kpz1FoQulIXZpN5ix8hN3xMyRvC20K78377IZFAfSj8qkTcQgM0b
3SIfniUi31301DZNBh3TTxCBPc6XmooYpdUe3UGT+FEUt+qonxTrlju2maMN6GAD
ms1U+Jlq4wFgeRcc6FPV/EzG6drWXZeAZX3iyJlUHsfvcrWpCcV69jCqtWkxs7pb
n+djUttj9FCHRJr04TrEcUSRQCPFUpkeopnPEZW6+EZ/HUept+ZgB/L6OcaYlC60
vzw4VBNRy+g6f8ur4eETes+WuNGh+3h+JZA9Y/Ja84O02g5oqK4E7Y/9k6rE/06I
ihYqtUGic6fWxkNjEW4gXVAM5zAbs+BfX1tx3mQJK0M6dOBkfu7bzhwPjxvKcWtW
k5mSdQMqWh85+U0HEKEdtvRXcNk2qKUZVieTyZAARO577Pu2KdGrYtEPxUuPEQnz
QxthTpGt9TyC0o1A2pr8P1UVgsQgOgAiQP+qYrA43IHx6go2VDcI8ggydpa66O5D
aUhLLB3dS94AmPAgaGWPUnSh4A3b4uDhBaGXVQaOTjQf/ojmzHfxtmsyjQ6Bj3x0
gKz8rNErgs2mPRUBJQVTKoD9OctNyeBw9le0e+LXs9LbflvQA/zCc5uSs4/7Fsdc
TL4T84Kp3bI4K0fEeyQHfR2DLyKKTBQnidH7XSPuJwl8d80S/jWe/tfvGLcDby/8
QBtKbOfkfrEm49cTZ5KH8Vu3EhlE1MnOq9XX2QVbJy4ST8l/6cC+/uKqBiLPMpQq
Jd3id/yfBvXMqu32N63ddXu3meev8GZTemDmf9piQOCvHgRco3cPN2OD1f5t3UKD
dezv+ccThfXcC6IZ8ldnq+92do+A6v1OT3c0SG8hDz2yALtHYSbxn9BX7J/vJ//C
Tsa5jK+/2seUQFjb76VmgwaZhghQghFtP6s5kBCWnF3vJQ7CJpy9DAI4xQDnsYnS
As6ITSqVKrcCxIwCCPEa/6dy9R7PYNxyzPVHpLY2pUAzP4n0TjrJDh1qOqGZNsHH
osKCs1QUSDtQnl+c/IJkW1sEr1Crbb3orblcxeJJ/Gpx30bRv43twag5ox2DCCSQ
1gKDz9xVyKI/kdQNlQJ/XHP+GotYhLpsWb+g6SGVOV801F7Qye0f4g0M/rLX2L8t
lfPbAIs3WmW3fHXyB45A9ukr63BGgVODeHOTrnAXHP6PTQk47OlxBgKMRFmb+Xmc
PBfZBsjDCQwyNtzdqhQHwb8i5VDa9+ktWkRV66c00s3dtDURLXcR/HkZbEe+8Kl0
49JtkEdqczRdU7aqvLpn9PBELkddJhobcVw2C/EoGQlKfoTo1k+LYGxq4EYkaaOi
i2ZwmLaNEQNM334vbMa0nMc1/IYcJ8jLap4Lu8edQvgsHNjNXvfb7UFY/sXwj5jS
aUE2x3yyJZeQhhedpRcTWXVX4oOJKYrE6X71skw/BBFQcpPF6cdx2617Wd9TCItN
VxanQdQlOU4P5hDHeUqX2YD/X3hYymO+xq0NO4MJ8WfWIc7socc6BzPllm2rZWFm
ulynTzOmYbfUOMZHwyzCeq6NiJ/Uu6B1rB3l7XZrxb+JWOrwgVnHOL9dgksB51N2
d00UcBdmCWLMkquOv28Vf547BNmltmE+kH5kMPMtCQ80IJwoobjIb2iVglLRHoMS
SYPEjHoJG+mjrKE+lDBukSgJFRfoZSfyP4NFf1/kzREjbiSmlH1iWUmPylruNuzO
dbi2Pg1u+dAaR4o5ydg876lzxbl26oXwnYF+dQOqh7rzYCppkLkMcrzv85JmJkPy
ueq2ubmn+Z+Zbhy9+USZLvG3tzSAhftRrQGjNU7vM6vnPMNI2ixTq5PE6exi3D1i
6Gq7mwjrpzfrNQu9lVKtGiLGWR6aQCCKBtBYoxaIyLBwKgc6Btf2QZuIni/2h38S
3pm8RX1Ol3DcHKaoG1lfeuj5CiHOH6Bc2XZ/TqMI+IglvaJQz3qEmbezJhkMV70c
pPzvxWAcHPCMF8/Ko1wO/wUfzzP4UUeCPj8ja3DMr/Tj3FN9RmhEQ5TIpshJA1mD
VPIj7qXTxXvEolYYsuRDRJvSWp2ZbRWbRlEb9RWbzVCpFudM7HoV4NGi6P+mOpUw
wBkfi6974hd9Jl/JbO8LuscWdVGJl6PC9YCtRb83GVlHNmqY2tIS/P8YLAATkm+m
ogE5SaKjVsF9/Im9X+uIDr8s66bj//UXa68eYH0PwwCHQE2eVrrp69ZaHVLcS2Tl
gdd2NJN/GxKaJT3H0CpIBnOv+vn24XkNHR+iOWYBF2mIrNNPi0Bktwb87NbwPOvd
sQ1lCl1eRFQ/Qgkw3qo0rCshr5lgrqTxmVhYTAYxOlIlVpQ4rTvBeWk/PJ6remUk
0uGyKpM0CqIzExMHRPxsVmBjyzFX+MS/TLIbPNEY85JO6XqBBSHMILlnvlcuuJvT
w3n51Nw+x5apfcZ0mzrukAaSClKpii5ErhdYpywGUC5LWQFjHmun+PlKlbqA+8S9
BfM4YoNt7jpW1XrfHU4IyXuSyYT5wqWNCGbgAMthN3+k64Jpk2AY0wY09UrG78gE
tK+i1e0shqPxFl1VGsb0kYWsdHAscBARqTgn6jKocMJmrt/lUdUCicsHdhs140Tx
0/ZZ5l1TEPCEsayQfVT6FmTA8KsVczA9A0H/2x3vSjpzFFoQveUZjEGfyxfHfWS+
MIUdf4HzADOKchQ+C39FYobHqP+uQMEzB4H1LmjOfoCPrdb88MCyFBOpvZOq4ldE
yKR/TfF3OgkKKNywfX3h33ukT3saujQAcuqcUDp0xRhbM8sIqmzlSj0krNRj0F1Y
JjwdOFFOJv11KphnpnRMOSytqmfOjWGW0wl7aGxa5aZCTTlAvnUFWuzQ8KELhxX/
VFmjg6Hz5/R/VY1suOiqa+8N4YPBpMRgvDQRhco0CmlNDI8ysAzkM0P0z0IYrBsj
q/TAsJkmHBkRvuwRdzWhELaPOeGT9jDqeDskV5L8iUKEgkfCvDE0hO/B5hLusmCz
GjGgdz+joz4hR0FeaZ3X1ZuSkjorewRG498PpYICsX6Btm2KTvYVaj08NUf5sCww
ekhx38k7Q8ac2keLfUcwve1X368yU7PjK6IX6tIzK4sVLYp8oWNraiq4DL9IoAQf
/Eu1kSpB/MMkdGZcRMG06BeE2u1hI2q+xSz/W1bTxnya/G6VWtFsnVV+Rc0C43zk
5qJUL1UmJuNRfSHLTMteWvYBJw32aizCx0npTYg4H5u8K88tlYwkL00PEdWkkGhe
0i7abiaX5HyzqNbl4PvliWnXdPNEVVG9AEhZL5OnmDRraZi2ZFsqVibKId8dA+RC
65Xiv/mwGokW/+4sWRXWxQhyj0S34fcT04rX8Jzdfs3/l72tJi7OslCcUZPMQDn7
0SxQx/qoKnXxVyZoQ/QVHG+WR76+DzRP4xIk+LKa4gFdXFs77dPuz69BzSCJEZm9
wwkeKJjJYc8PkQbBK5NPkWf73oARr4hag4IX2LxOQMqfJp0wP3VD7ZPU6J26skYs
xydvIqSuRhaWefTWxCs2J9Ni99RiamkFL9mPj4SE/4291EtBRPuPw22uyY7qSO6Q
k8NaE3/SFtN0oDsBUwa45ON2KIlKOEJLZipybjdq4hwkFloyRuj9sukwcgaYAABN
wqAO7iOC54rJ1CdJNC9DlX9jxMq/HJiP0kel0iAWTTWZwnKY/y/6+Bhd46Ck5pEE
01hOk0tcF3u88MKTdtIqvbgpew2Ve4lhXI/jbmRaXc4GUvzprVuAbShto5fs7TR0
hJpfeUAMS5+i9d/GnnHgaTHxhyYrdwkn7gTlVJhh4CFST/bfzu14gWoW5PWzpprK
Vnwlks8zMUHtdxjq9ABSzQoYfq/t5C4JYfAxfNVpOSoMjb4itvFxoNtbleOV0JKE
PVsu5aEmdrBhUmIPHSiXCLegsyQHp8UJ8RDJQjrko1d7CWMrA3LYAW+YIs6sSc2M
Fneu4xFnlGl6qonVujwxk+l/FrEkZuZTtvs4faWkXncJYlBYnnDpM2SOTjsc68jU
Pn1MeYDBdqjG0Uz2Fh46d6XKEjh0jVrWKMpXYBt08zDpRaJ+Bg3D+kDGR/Vyepwm
UCyCOhX8YD3e+RQMMgKnA6mrni8DAwuI0XSXYa9TalghDq48SJX7uyUX/+jnL/3Q
C/LWa3kqNfQtVxOooOn9RTz6SDOhSpUaRIwSGB3q0208ctldCsZTa5OLXiYuMoCU
626DnRRdQ62vKeY8QfuB/k2Ue1qFswyLH09f9WIWHNi0/SJdEO5MUK5P5KpTK6qI
xcqCMSRgGth0YEYhLznwj2Py8hRQ75nsOHPJK7FZ+77Z2OULguxOY8cWmGEo/4b5
2OTdBo9lW0WPp3C5Jamq8UXSh6yp262nmgvchrNLbOS7Nifggx5DPbeF6/ULx9um
m/ns0VyZ5QvR0XKVK6Be9hXh0lQecLpirHSWoZd63wkufTxSVx3wxLf8o7mbF4aJ
d1rdHNDhP4bxoGbWrlfGnE0pxw3gVXbJc3wl9RxGFGigFDJ/c+dYGi6Ob9b7CAEP
ff1feo0Jl0JdgTjOBWo71LINCRhibr4Qqn2teBslzvADqoJ5rNzwfTDLgbSox1PN
fgpgqsVnlRqPv0zUZRE7l+GzCvhWhJ3710kxuV8wbYALjXisFdaK9/k2kl4ahB+h
QWpSOIy435L52V664gTJ+IbatNqwIeJQXKw3RhrNvYnVQEzL7Yk7H5WGGQLZNePT
BQs5jeMpss31sHYJwK/eiX4mK83Lj+EP/koganP9o4GYIX2OH6RF5tBe3mEjjvbW
nviFG12SLJsDD8zlhgJQFd4y1aSd0tJyHdEHselWJv0b2XysmfMUe15m24yOjykw
eNG3e2dqJw5OauCYIWw9/9mCFGNqq6r3od+bydN9Ca2tEpDLaQCwK3unpjkOYdeF
UokSFCe7XaUaenpOsgsbUOfiwlixUZ7sYeEX+JwmoLDpF86tKIIyjEDslLFHbpzN
lsFYopSWYh3l011Y8Sj1/6ViibdZvwYDvzI0ymf5dEloQUb03dI6Ynal7Nqzj5v6
B08xO21FqM9dMaGUKZc8GpIFd7+mxnzCFaOGj9WMuAfWKmM6gYZ4FKUvIkwOICHF
Ssf7zD++odA8cYUY9Wx+AaSnVkyBJfXkbf2UuHvF2dX10LbSOwIkO6I7VdTiRKTe
WuBIFbpYNWpZfPdhI52BKybhF3ZYtb18n7wRJZhX5kP9Wt8LDGbKG3M80QptJ1fh
3Ppt76o7G95X+/AYmbEhG5j98WRL745B5V4fE99Qj1P0EsUcDG+tNCLYPFEtY9DP
eYdo52sAbD1+g1aXvAWamRJkwSLPL81jh5UEl+N1Z2UxykEqB/JfARxDvanTvAlX
bZ94BsQGos708VmeU95wmTIs/JMK265tAVC0MxxCpREse8PaoB5Ek6/FWjULZsp6
ZQROWVGIU46IXuZqNCKrIXMljMX4ZZJZV/wVpx78N/1iS4KP5tcfK1pzsWogrBP1
iIu77MUJ06i0OrSSanuecIAyPkXrzwvlOOoJYFLf2C6lmd/HJdIN3bWPTyzxqpM8
QYjd8FIMgLgQ/n7KgEJdWnVn5n8Yq71yz9z8qBSy0HkREAeO8M9dP1WTciOWq3Cc
hrzuy+VdBcjpLGTxSvpPydc3+NTrSs+sOHy2LuT0fuCnG4dFLzCj9FXFVq1FB0YB
mCG7RnT11YZsSCDpzgx38qmspAIaVVjLA2YpHhhPNIHpYGUt42mQc2dBoRYIS7Vw
LosclEXHvSZU6vzOpu/lOrtaErSAYkWoG2kO/UYdIZ/CC1PWzznIphIdNvjzQV1H
Jp/Q3cPx8xm/+JiS0XFxJVf5ibTkpHM+HqZX5xUDcj7xUFkMVp6mr64Bivf+VEEM
23NCa4HaBo8rn1qbOG0jXzBaAx2vRi/TEgalZo/QmYuaxMD/Mujs03RkIkpIvDrS
WIktV+F45E6gxZLx2DxAE/78KzHV0pzvWsRDizbzWgrSFJz452SKLl8ai8/Vddo9
GMyMoRe9sz/swUArz8uAHKiGkU8tAp1yHCY2ZkDbRi10+S5Ffp7RGDFEdM5Z7ya8
ZidK7UASr4p7DQ0whEmw6RXDYna+zTyZ9pYsmTD5IJ9do5bdfLb9tSSEB7PuEsXV
SQTeT4Mt6SjfFzk2bE2ry3EYdskR47HTWZLznBz5QybFssifvXGLZOmu/12vSRXQ
v1+6G+6HLGyuhB64hXYvie79h+0lRanO0RjBol0PQa95pVWdCL0ve1f/BkSgcF2J
IKsr7LYBBT7771LLbHmEfMrBRHyhJnyax9Dsdb/hkgI/MioWSd/F/5fVppseJkm8
yZNEJb6fcjxSG232a9PJfnWHbxBqVJV1aChnqkkEl/pjwvfupPg7fXbikmUm/vxL
cX84ScSHRKWETpNloe8tvcSyuAMqh+qe5sbw8xmmQMGl4hh+nPZdrSUzgq1oR0Qd
vqfJNbbtVwa8kmJAO+bXFOztG2ca8KWjzFIK5F1p1vuuyWcPGamIrfm2uIk6RpSG
DpaWNjKkCF3O33cV4R4JDBzhVwTYOvYBMBl9BWKfvSW3prdF2Hq3uQphimY3J35b
10m8CHPQWACzAZkg99P23Cp7nl90DE+36BIvAC4EmBEACO4yfWYRJfnodVUwcPhB
mAgmALiiODu+nRlvkPdaHrdQrKlWHdI/WyDjxqG2raGryRF1k9Pq8m4q/CfI205x
s6pgwJoEWjkRneqt/WJnDQuZtt7niaCJdHZVxTANhm8ljFQkMM2a8HjNV6usfz/N
iJNawP4N+FAoP7gJ2nNx+TFVWo3cYqqJUIJ+bA0y3mFSRhjxRomsaa7hEAhsCWww
6Nm+FMDb0OdyTzbgPW1xwsbvk0jFJQRDbNb3NetbySY6bJvODDh59NwSmgL5p1P2
ZuuFQo9TXevBJEZrUhNqR5cFy/uiqQbdvSdtMV0nwx7qyrjmGttT+Oq8jWQ2lF6Z
lMA6UZrsiK4psP5EPfPJptctXZUMnIshya0HJNs0BxFuBL1V/o4bc5YbsuGNdS9L
yL4wZKp9HlworiQVM0aox1uJV5a+CxJEQuCxDWhi4s/7xqEHtTkQ6Wr3P3SGHvge
0DU5Yfgox6eB2seVJT9feMceHpMO0+nCNcKYvpci/QA1/REXnr17bCaKV0bsi8Xr
PP1qDGfiL4CFFUf1GWe8zCo6RKHo6v9UDnub3OVOeNae5BsbzAn46MZq2/gTa2pA
g5WtGXCa1Nu7h15rhYrN9loCpsZsg3RyXYT8H5GMz7sio6UlleRfnS1LwKE0nLmN
LHlRc69fmxEsAs/6y4ihnBGjbXLjtLgtEHCGOkXbLFYDJ8hdVdQfgRH+yEsyK1X1
OPv1nWFck6eyf4iA1ip+LO/8HSbNaCx07sPhLsRlJlF7gwm+EHWCLsU1U851AjPo
tpPbwyuUVlzfJn/NeUVf7WgtQxqnPwiIU2OghWHrcGxSr0ZOX8+EZBEzKvpylvE4
VovW+8e8/UL+ImRDEa10+XWrZy/hc0AbbiVrFr2PqOASoTjI2hOsXlW+YYAPr/G0
gFVt4WcX6I4SREFccp6y/56tMDmVlKclTk/BU4F51krOwvtzzaBZLPOYF/NMI0Ct
qOjx9RYw4NU14/MlTz3NovE0wpZeny6XNxwvdeOjzXNCMT5xOvju7jWyHJBVqL70
oCfZAGAWUDFoTOmYwV0wke90a6mYTimiSUhSIVl+PhYn3oegiigv490jQQGOG6lV
bxTzBsQkQ0XvmbNgKE3/OPVzAwgGFL4HuRiGcvlDG840TbejTzqz/mM2LKJGeBXk
qhETFasaxkj/nYB2ldvrN2V9tx0pNE2z2jKoOPfMptL+Hp40UiAB0FSXsY+r+ILX
wMloEkcjJnV2XwjBZjTzi5pVjFd7YItORSl9Ih9QgMSCN9dG7J3Xbp9bojEFP9eF
xe32eJ1R3EuEtO7d7auLXKrIH0LEBKwmJl/8zdBxhkv4dVaPhi1ivTG6EpbJIr6A
VcjXry8psg8eoZK44ORWnJYY+49pprr+8OiDrzvbFAyLcVAerSG5oNK4L4Wu8Q5a
cYIYCBorGIj+rd46zTSs4as4IYC+v23zser9JjMG8CQoxzIXcr7pdVO8zf1zqvWK
QXIUhkz/Zgwk27RHT9CQaef12MMofn085HS7oIb16RWKpl3mZMFnEjKCRZ4cyRkD
dcyRD5uoaTxuTsMXtseItF0VqCKqnQnmc1nJ6YizjRNbn7wMRUz48I0uzlJuBX4x
WYyb+Wq6M7HV9SfQ7iRp6E3tFO9n6jCylitP9KhpnJw01hxB/DWvDBCBPBZwOiVz
6H0Kn0gnC3E/os7g3AplNUeKYoVAc5+Vn7YIOMzz+ycCpnVa1ooBadG25SlwdETl
h0I1qFKUuRd4CstYGPiExtS3SG/UVk7tX86EFNkkp7t5/RT+DvUFcZHyhYdM6X0O
AGKh3wErJn6wLgq/IVbV7ZNveCyk0ihReGb6nPDrerSdZyvCSQIwbbEJyjhsc+QD
JtIBiGcUk+soaUYd8HO6Nkq/oa6uSPfa5omSvcd/jRYFosTkrIw8qSCr6QeDy7YM
k27l0wiAx/yy5TMjCWo6fEBBYr7Ihq+fyHGHpQ0G1UBa6hwfXVylE7TVqS3UyTG7
fWTGI0SLtyW6RyEfeaYufj3klL+04o9Q28fUVRcXPJ6RW/T6X1sD+DmeGpAJmc+c
yPqLYVgDsAUtkB+6Ie6bBVLWInHjMjcJakGCFjat6/OPkWGSAlbdRYaBugZ3gC4A
eXBPjg0RP6+eDlZISyyADYoe0x/flCojxOqPu9jmpx72FHKvaVGezSuMww8jy3mH
9BDyIYN6OVg5QkRNTo3twTutQFdJQMn12gHGNyenQRSZj0t3AgOuVM2o0thLIjA1
w0aHnZ02/UZ9ZjLg220qRxn4RZncQPeMkk3jQ+4o+vxHP2piym6BXF1rLIEW3COG
l64isZvnICRDxc+9Yrn5Ue1IIwRG/cdzgIER2wU1LOYaxuHqXQli+2DslMAHrrs2
DbtY3MjgsCC3cLvyOrdOuIYG9FH8KxJy2qbH8+0e4aUx//xJuAWfFQ/65JxW53xX
dauxbug16B15kTvbw9kuQ9jBvF0SnS4sZMdS7cjG02BdFBnhP0VFKWWnmFJgClia
t3qjwN7lqIsVJj1ZVENDA39SVBPOE4CYWM4kywfIG1TBBjQdEhTTgLEhU9iULlYk
nm5PtY7wK9UyiJYNJvy1hBsWceLcH3tytJprFle50UAZ25JwGL56RFrf1YoEw2wX
zagun7Y8xP8VWAx6eeUqvcD33AnKGX3q+dAma8i1jdrifojc6ty2fIV/Zhi0rgwI
CzzMMF0UsDYQXtEPKFIhvkuLl/uJPBGS3vnWYpiagKptkwsf8pDjMKVVaE41Gpnm
0LTS3Z4Z2IcoSZgREjIZuwn4N1T5jBhReB2hs5pppntMOGjMWhbYsE1ACtBKkSbF
Db33EqSKaGzPC14+cW8T8y3krNW+yqqXNMCknnxk7xbF5ncfj1S/GFAXSZzIqJCP
O9U17SVtlHpyPDW2ip2BURhOtMGimIZYX0r4OcePpggt/HwHfDjZTf6YffNL11/w
2OK9TIzWV3YKL4vrQWchhvG+2cW2f8QWuj9f+2PFDyGpOUBELL+V8VDSppDzucrc
JKMLmvBseEOkj0U2F61jlQfDxzK9j1zLu++07Vn7+tBCSS4+oNDmNRNpq0EFs6u7
t7iU4Aa6pPYiHjw6See8FqOg0JY+82f1aBMs9PrAX63NZyrgybP+w0/Da8dwGu/f
RusRnCmCJFWAfn35MdEkJpKExsX+EUWk8bWc3cpW33KKgjGoJAU7ppZqF9HHEaDd
t0+1v1oV49KeyFYso69O/CXAaSNZMCRZjTMxDO/YG6WmE1hC67kp90Kh1sEoYPgh
bQI9JD3UIpHJQks0Bu4z1/p5W2WxvUR9fwkSyvjcmgP9bsvdQXon1eBjSYEC52Qw
ptM8jkpzLuYq5MyM8+iuvsUUBEQbYvht0v06DvKAV6YU4ZkkqR6j7Lbx/vmo+nlV
83CCbo9E0eTlLtxVFW5XgSChqonzak4sxAnenCaJpCogW/aA9EEXUtgS81ZEja55
22q/nnGBUEPoDCVbB+tGqX2ncbEfIzHzEPrV3X3hcVXJvMqEI/O+k6eTIEeV4pN8
em6lTvtVnTXnZohYePrvFhCS5xFhgRDZBmSVNDE4sQr91jUpEDc0+ozU+1MsI2kR
PPmGj6wtExZsjeZq9546Szh66KAVVhag3Qt6VTGojLaYqbCjcd0XYf2J2X6SNfOd
QNBJiPIePHch+Llw9T66DZCPh0Lef1IfjciySdf7YeCqTAP8v+kx3RMxn1q+Wd7s
ion2y+5LkXtvN0WfYExL7PJcSbfx2HoyuSYZiJ1OOSdyXh4idBTMo4QTjRIF4D48
lPjdu6An439lnJ6x7hslIkxCmkQfvWdmPSVs5Cv420L83lRriS4/xz3+3rTPVrxk
/2rX0rTYoiwXpXso0RSaAk+KlLc33I0oWIrJzipwyvhgXyDvlX8j30bZmgOe3BUX
Jf9Yd2K12fbV4Gmxqvv+oWBhRZvD+Bg6JgZVjNS/+D9kRproJI0tJLx6rpZk1CNs
l0mDX3GBOHR6echOfAK6YR51tmxZwTiTB9DYA/BQ6LACFxsBQkp1RB1E7eHiNeWf
nQCP40bbxVQzLPqs07PZ5ZAPUQFMeGmcy94yc1ptKRJlnc7Cl2Hs2XqwSux6gGdx
zXmYIZEZXB4L965NSK2dy/51MRYmNYcfeuHej08uZ6mansWjLpdQnUarCW5VYmCl
PWMaWf96O215vPjaZ1bJWNEG25AdTvSyOhQrH3B3OAatelHKpXaEFS1EQTwa44p9
UhKEi/b6vmjBOCIcp866FNyswmdMsp464k3/pv9pOjba5f+iR6DC4Jye2AYxDvpU
WQN/E7ep8dNbFBUuAe3L8heCGUdYgQGh2Fkn6s75beQdBph/Im4aNBNh7KIEoQXk
o5TVVs5n5hvSbUuiR0LWMMlCsbJ3iBvbyPn1dM/Q3YjJBrere1eqPotypqETNTWr
tfmTNjFSXNn70xXex8Et0sbujgTeeczWw1xqwgH4bAO1l248bXbg1H+krGWbCxk8
JHMJshhn4qkiqAVzkaHOs6/G2RM7KFYmKCpeMhjQUz5nUncOJQom5m2kvc/Wsx1H
3UYRascExdM2oaOZF96VE1Qutp9Zpyt/sRhhr1b9sr00y6d0jdKlRY/iBhihE0sx
lyiAGjfLof47ozztoV5gY3eo8tmdrni/ccLf1NPVMjZCgs8FslsGXL45R2w8zJdt
/iYbiFKYIB4RXqvni1mQBYhPa/ehtRhMp3JBWCVr0EKyqY4UbV9JlY/myW+G2s57
3ZX2cOTyF+PMqIkDm8Py9Wxja8VKEqxJ9ZjZjzW1vhbCBQO7ygUGFeKl27x5diEn
2iorq0idGo+PtXyTPDHX1DgDr/235feSWaHjNA2LJyCCT4FO+/G9q6kJArICUaSH
yipCqor5zUz/FI44GrgjMbO5ljPQYZ8yzyIlAPZ9oi/QShtmtrQVh8KaYnDMXJBF
y07h1J2YPWPASxq1XEuHfJbNKoL5/TjQLZxn5tpPuMNM8F2nbSSAbxXnPui4JiMH
wDo/DnSMUTWuOxlKkT1COl+GpiZCI5PUW7jEwB9WR6fXnmB6351ueMP5vYxD/ts1
msb8BxrNZ+rKJv2ZzX3ucFaO/uSMM5m7WV5HNzOdaUyDtNq0IIzTjnqfWI/pdvju
pvXoJ1vqnX9LrYzVQDPHgcsLcOhqoROBYfCxtjRBQm/7OCw8wZtaYo99aFd/inWj
381SH4WQqYJbIYEIgB6XrBbPftFjr7+qrzHxkexpcNFXchRMVGmAg6kr6bIY8789
LEsDpizsy8LwA1BTCKU4wq6xhsNRRM5lJlbbCm+hoAY2Xs/E/XLzlQhbbMUq2AWe
6zQKh6ylfhycJ7J2FXs7d439WAoXud0DT+igX29yIRd53qn1+OblcXFTv2qAkPFC
tZSeVe0pCu8dq6opzYY9hhV/dCmRyHGjbAP8a6RK4x5zjv4jtFfi9EOVzpC3sJKo
k7s203PCepC7LK71MLR1aTUAp1h7vEn/be9rumtFnvWp75F0YNd+1Kay0mNFIV68
9I+xigQ9OsFfs0d91+gFhDSYximgJSEOz7ZkgcEPSNWMgjThKWaBEUHMAtrHeBUq
xpWu7okqHpxWE48A8nsYIhqIpT5wUACyjh3joW9SU6BT8a0PFH4H5JbUPn5F5BUf
qdV1BHVfQVHBmghkgna6CJWV5LU/K3Dvx7+bD5u1hYLTWY16zXSgWCuxtW0fKU4z
TNlBB22m5O31eRr1MYfetUSfT/Bo0oirHAR9Vn0ES+jGGPxRsx2F6d2NAVDyIo+e
HxdeX6+7nCaxo7TwT8MciLuU/BMlTkBtxUcYCC9aJmPTXbZWf34tJ23JpFg/zb+g
6pwPJBvE+svM80grdJiVxjQCpxE2h3TBOu6s6IFcn65x2MJLiZNS9Cptr404iYhD
LeM7yHjqETW4cszysVArPsQu8IYcDDpZeVWXF+AJ75VZKe71yoIPQkK6EUeXf2oK
UcbyB1egLRwV0Ig6xVRUXNcMeK6D02hcTdiqQLhXq8SkWm42M6NVGdyyQn8cyQ88
z07GzgPS3EnWRuJa6ykzkgnSJTFh4iZ0gbh4619AGpOFIzP/Cg8iBpnHewN5p9NM
ILKst5Uf6GxxGkO6T51YaXb/oEXYxgV5k61RHRLv+m1bhJolfC4Mt1goDJsHk51L
5h4k0SV6TjpJC1C4c8pzr3SmXo+gc2VwK0tcjKkXUME2OlloXZMzXsjx2Ad/Sex3
iX7TBELi0oOhmx2utsYqgNZ0sluUhOJYbmsObKqO69aniyCSrQLcMAcDnU8PynFq
vrzNHjyXjFXFW0clZaTEnm7leb6vTfHea5ZLy/7isu3BZF2TX6cLSZNFU+EQcwpA
yLOQjFjbxMjxeyWjJM5ZbsscQEUTgfFEg0ALjr1noknPpPDUqVz0cGrboPkY0Vme
nDOjqzcqeqeINzPhvskjrJdp3NwlqUTIm3Bun8nPZMx+UHGshSkQT8SbLZ8v0MoG
0w9Oht5Jpgk/zxL/kwCLIUlVHLnNoAX6/Np9fm4tCYqB41tCaPVo/vzwnmrvgNer
VNMWFBBFerOU+ofYzDmZWrZBKEiPSA/2hbsvR3bIuQeEFTENrJOP/k5+smq8MCkf
CIH/ifSzJcoN2QDTkFXajNFZT5avTA3ug00PWMXLKfrKuQr/OxZPZL94xhBd8ZaU
NR6KmcqbkFI4s58Sz86RqALcw1PoiAkDSyhubd1ylI8rsvnxUynz2Nl/Uy1H8gv+
dYmsn4vxaWaONR7Ap6SqB1NoBU2y9E8lsuvEEfSHeSF2DXTvEaQoXQEeyqEnum66
fmX+4BXD3/DrCLmJynVQ2sFU2CS2qj2cZS3CTDBK82zB5k747I4pAHwidNXD/B/Z
pQ7uDtGgvwZifaV6/08AiHnwtm1L+VYtl28MoD/FKt1j1vVK5NTJEMPlRtV/Mbm/
4hI7uQYI0yCZ82DAp0+E1FwxgKZpOiyLGKK4Qxa5Q+nNrY63M11JiK4jdWiiMvJz
4YXWJC87kpRIrO/vjwdcVAkUklz7EhbzwJCnJpzwHSdjzUi62YhDFOMLZpl0Hhtr
6sI6yWFCerV3p7ryV/CpWHzI/mOu70JOZq3NoRXLcqawnjM1S6Mhl9xXLFec6g7S
4UWeeBFYt2HCQDHMOG8ETO46XPStttGVa3ICjSEJ2BLCFy2dnRDvL/EaCXy0diQi
j5yqtdmP+EuwBCK9UMqO/eonF1i/MsQElEoKrRXlJoX5rXMMyEZzDdwISvafasHZ
URjYng1fLJKtkayrTgJ4RHHJzxlb8gI32nYbJRVST743A7wQQoggSC3C5LPl3xzo
Fyq9NX/CH7VGbMTGb0oEitxaYabqnIwLEaPK07QDmtRK5l80tH7hxuTrCcMnQzO4
oORVyzu+CvXhbVdAb00GkZFTuw2vrSSD2wVhhTuHF1wLkEHVkE6RngRw1P1GZrZy
fSKH/UzqZIdQNIwHw+e8g6mA90lG0qGBS4qDCmUWVd6GCALeRrwCwe1BEuwcgnrl
OJDCAuhtQVDUVioj4mA/UWUEkQxQ1Pv3cIZR9O7P1F33UspkcImwUTW2p84vmPka
itwcGlPzwH/oz2wvMrLSURfI1fgQjQK8IjbvPORd+2LVZe/U91jHgmtpb5nZ48DI
DnJ/b0VbmTfYwZeifOpOC5D2KHRA0VJ2G8LPONFZVugqtabJQjkDRlOZmyG8ZP1R
SG/ZVt3sZpyTOAm3slsOwxJAf4flYM6q3SirBHRSpZQiJZShG30lfHF6Me/B61iW
0s/I/U+1G4isv6TJ8NLzlG3eYOTPkEO5sHLyG0O+FiRnOnRrcRUZzT6xD0ZN1LKG
4Kbe2sGa55V+riDOLk1Vsh9A3H0CTJ0/CxrCZPIzbAZNgd6aUQO9adl4VA03tL+u
kay562L8x7J5Mfbt2qyi+U4/5bchqxluzR0+9h6Vxmc1CYbbXBdWzunZgF1dZI/y
U8h5zDyWzQCEcwvcCr9/wOhglMcQXdjIu+bwo5tm/U/hWK+mxxfMz335oB6wuSqv
aYUDlgrvQ8elw0FnWHR6bXnBH1CfCYPxYAISsQhcss648vVXy3xqjZrYrJGpn5dG
rVbyFHbTWlKFCbzP/J7xyXmbgI3ccOP4dS/c5X/pHYZ0+QXjllumi3JocFU6/G2E
OaneDjedEcd/JDIgCpB8kCggNLACqiQt3F82Z0eiHexz/eMIy9AFB2UgA5Zz3SHI
ZlfCPAu4bdzXYu0SIJqwfnZutY68k8EOi4Rw/DBnmc8SPrR3uPfB38esviwI9WsE
0x9588RuZWcbNX0iRFcHO6zD1xnehO+VkyEGTrbZtaw24NVouT4/tUXQrWOmLTyF
snCyZtq+KefJCSm7phrzSXedD9Bg5yEW5XdzSJqc1xD1hOX6XVh5nhEnd+lziYB0
xIPgS9GeGlY0gsRt6iDP9DwFyUgfVPIyzVJ2BYsX2PO7vqU8tsdgsvc97WOccx/C
ldJ8I94C0SbH7rWh2RH51PLKckgXYvvsFVscX0mWTzmdhCPcZ2lhbscwR/Oqk7IO
86KL3zvTfQm0WmnUvAJ0JplJVovMrGgemlXvdQkyAD+boxlvBj8krbz9cRH1W66c
rArgjlG1/3SWzS0clr26p8075/CjBspAzEzgKts/p7auhnlvJ/k86SPnNMELr/FR
n9zF1VmqeMas8cW5Ws52GkLprg4Gf7gMS2mOWn7ieqRUwLHQD/scR1EBzfGe9rJY
VR0baZ6DCQVLlUo8U0JWzLkNcA0if0dO459DReW/FGw=
`protect end_protected