`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 3584 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/9huKRhRMtvnNqb3Z+UU7TahEoHV+T8U3P3ufru7l1O
3DlgtZzb9QxCbOjthp9+wDkjygH0eUfDrEl1ovhZG63IRSP5AivbgSMLGmKo+m3U
mtYphghWBA+FOMsoWrFm/slhAlOLOGyFTWPnuaWjFcqM3tZBUmrcR8bSPjf/0RBl
k1K+Y5TauDD9Z3aHYlbRqaMXBiHnkxuk0NFY6onOHs7IecbHBn7BDnffoMOfYZWF
un41xM+CKR0oJ6mqkY60MX6JfVr67TF85Ri1I7DHEVj/vK9/yuCIhZCGOxUbMs7N
q+cGcAgZNpbKU1mqZ8OEZ2LlKeJ/dvgWqqFTQfhJtVx7cJvlaR12xnfFkW5lfsDW
VH25P4d2Zlq9omur+3U2PvGLHq35Mbd5QvAUWo++3PmPa1t4/AnYBkEzSdQInitZ
iSJwswbgGuI3VxuwaJc2Jj1hfe00Q9VI7zKRfA6KQ5hHH7/IzLUXBCmXZ02KthW6
ITQBc5D1Mb+8PxlJYPGvyPhalS9IcV4W1L4xKhbB7tQL4crOqbolv6RcFxELdh2Z
DCmT1dp0jCCQ85qKGfr1luSmwFcWcC7252r/Rn7HJh3LO2ZwGeZT540ipo/F92jO
zjk9+Td6Kv9UNWhVcgq7VXQDzj8jZEnPMfstlmMdNSXzOOEPVee42Xv7TdrQg6Gt
jM/de0PvSbkGGX144b+1OjMpzolQdI/djET8oCj7fFaAK6+Aa+8nI8bmDNLsbDyY
zWxNfvnVDD/hNyEm9b7dHe70agLUrFaS411oKrdL6PdQ8ZBW4saGq+sziRZOVRdP
gw6PYcxCHvIrguu9oX42HHAkaZldonyyVlqvB+UkBWRpHeGrj5Q1WtZanso2Z+uf
2vBgIFQGL5Obj0KT1/vRNjNVsd1/tMgdyWWvtTSAm/lL6w7ZS+7BlmZY3i5LmwE0
rXE6GOPUVQKfR2WEy1PuOiEsO4IlKUyghrUVCEZuDlJ7HwiA8u7Y3Fapt1iWRrHR
HmrPIsiTKfGuSEx6a64gD+tmPiUOHlep6YKjyyGEzNOa31BuioAaZNfwRbijtzgq
N9xCynlV5AJV6UIlt3s0lZFZW3Lb6fqivauubckegq4/93qTUYUvwJuGd9kd1EWr
5E6H/u2fDK5p4at9mUounURrT3CVnRW2geDRnVanuOhCmfZ1fjHXpICs3/nR5EoJ
VMcNB0WjbGleia1+rpA2tjqa2Nij+52Md8r3mlzAjMHmECpLyI8IDAyijxhL2SW6
UOaPXM5K1AU9ScGiZokArPGCoHt5YG4HUeddNpvS707VxsnVzdR38atXsWYBL/b+
EsQGnYgVe93VbrzDdv+CKzy7D/gCien+Ct8FFC7hhAsP6D4SDgX2uYboTqY8Fkv+
bMm44b3NgetuDI2xuhMhec1qceiAjuWSLX0HxLo+hjz3tb+W/ssMkg3GcdNs+ULq
cppO/WaGQGKYUKUyMdFTeWSnytj0mXb9eIAnLl8iLJtoJ0PkjgZreQI5Z9NHj0id
m4fCyh1hfaSkKw/ymyWgP9ADLwELLlxRAss8WrJ0Q9jML9LEppJPSKkt/tZYulEu
zO4FOm6vprInWc9jrtFqSW97tdxVZosxmcIIfulNmbz2GBzfZqxBp7vWBpy6d6Rj
NydeXYeWcT9n3CO5Hp6RRgHRDwxPHFQ9490HhEIgRNAOf8HUqPRZrwbUZm7dz7q4
JeWeP3WoTbQzPNLGOzXguv+qsDoewCOpF4iVO+FbArezlagcKCo6wSjLyRpkIrOX
5CjJMs2wtxbCwms98sC29m0KcbWGzQtn8D6XCFMo8FZ1wsR7vLKw5liSmwtQK+Ab
Z5S2BPP/iI8jFTaRIhSeq3FtnR/Or38cj5prhdjrJ1i/UY/ztUbn3OuN5kXb+zVu
gJ63nOhHfpR8NmzWfYcpEt1orye4lfrMGBpgg2Y0mB5/uWNQfj0tkieEvF1CxsG0
QmNKfN6osARLtSGnuadaPZ4sqzkds9Pj/P4tN1ztKFl+wHWSHnDUfSEDBsT7rcxR
6GkYnGXnSRpSRNOa2E9ZwIH7Ik9kEBGu5eL8gGKliVrYS9bf+yKBl2A6Q+ZCJ+B9
W+pNsv4eA/s/ASO+ayTShbAOB1w1ENia6aHI1F34mvusK0ErpcJ4rymhbPaLHvhy
bxwGggtVOQeoJTgPHo2uNBDtz6OTPeJ/1VrInMQuoBYPfSVG0Rg5rQmUr1RyPPRR
5BCIxD38Hdbxe9P2iku5a7JWhwS8fFRWFJgWxLTISSxU1yhUOPCDaSPeHdY4PPzN
LsQ+jGqmlB73csAXdTYaNoQM4Aj5jsMO2+PIaenNPSA4EG2s5gX0IFs0WkuJhCbz
gBHtk1Dzw1kSHaSyxTtmjFn9PBwpS6TnwWtb2zp60YM1Wst+KH4sNPOBxKKmb8n4
pBwU6Cxk8S8RZfsy4MqgCsG0NoJBtdTQW/VPdIidQ9kNIyWP4pSc1pb2Q0Kz4ilN
083ViFICfSx3B+8UD2V8f3f5PeaOvE109uAiONNR/eWGkA4IcT2+PxWNpEbfrxDb
g/ZQqMRH0O3wVgr9ah41w8nt5m3lvGIrYGMKSwQDbzvoFzhZ9UFS8Q/bfdhFHIGV
rIHDd8I08Oac9NDKLP3NnfSMQmLQGWfDrj5dWNWVGp+9if3AfCBWSrJIDb6lkvrY
0yOTx5FJ7hRWGZ5vdUqqY37EKQzzHMPOqhiQVQAM9dfkFBqG/dPCQfBA8NOpKQ/3
yzGx/ikGe0GTArrmWwcOVbrUyMZanu0niHFVTpcz8JhLtlRsKAa/rjsfBLznDEDy
zBR0OjyvWycyPWnlAfZVX+qorotB15WOOSVs9c7zPaljH9i0Q40tmY0wtMxMsMho
9CWMbIpf49Aq4giUQFdGRiqZi2Q+d3hDC27G8O3S17GeMJrq6tK6ZUZIaHK+VhVS
+o3W78/o345VS0MTkaabUugR/Zem/tBJ+wcb1uDgm/92m+r9iN8nr1Acola0SjLl
YQjLEu+hus3sJwdTSk7DlXV8Tm6zrA7jah/O7DhhtNYMAQuaBQnEpGB531n/fAfZ
QonqTEt6gmwTXxDgKNlNYwuCsSNzLxHyqeIo5DgWZfmbZHhsJvwT7NtG8/Cm/y6e
JhspUIy/5lj69XQwmRLZs8et3Gye2Yf2IZI5NC0EXrGI1lwkmcA2PUMICcTHJCW+
VudAdOCqmN4kInlBYIED59mgTMsXyJRFx472trlg3LTpphYCey7qQl0uMevTFmEx
hNS7F9vKRSWH99YmGsgbCqAwwhQWtye3zu9Ne9yzhwlKWcFz892wTCECVTz5OuJh
dEcGxN5ktED092B9gJQ9vT8qGXJRLDUaJ3so0JceXbl/Zt2uHEgG+tndPNz84PLW
vvZpkuFV/F5TYcVD/JuqL3V8H7m7O+TAnb+aboB7/yXUBk2EXSuoQN92z2lk0xId
oXStbRNvpnTwY5b54H3v3Uvww1tyu5sGMJ++rU5ohDOhu9Aq/RuQsyNn3dqDxTNT
VeaXNyccE3ZRequnWtCibswly9X6BDkB5a/q+sRskK/FYFfxaVLMM7FzmadHM2ik
eH4mKhXO9xSt7dTstbO59SN2wV7WeHKdkz32JgGCBbxUUFavE1KDCURriXxHrZXF
QY17+V4wvirI1IwHChrrH7d9mBOY/ppKBW9ex9lKje8CjCVEbfBEA6pyhBaJ4VPG
qF2Tf3hts8RMk3Sl3w4yPsFr8cG7TwIrM9gW//NvUY5o/uj5lgQCFPaSTAvZVksY
bGef2EZI1porqxsMJtOk9fR3FTT74ThDFGYx7y2hTpRHdJagLAFoWnBfZFvrYlUz
UOCg3RfRwGGqsZfTp+ews6ggOeXgqWWSuSZ5BmejR206wNwxzxi6k0TB6evSL5TN
DsQKMuq75av5dbhAMjfnWp/dcMHOOPsmnkAJZhR56ImdTUW5NTnxyKT1x49VEoWh
9RfgXorizFWzpRxwRDplWr2+z8qAzwHzT4nQNJD+qsitGRfWbMW9XXGsXNK+dg3J
aFoMittOhMYuXXgOiQUH7p98/t1+tX/5r2pEukZAePksDuY3czU0uHzprvdy3mq1
ypyLyhXeAqnpQCQhlRvJtEsZltxGYjW18Jj+KWT8B64SMranwBM5YJ1jWYJPErN1
RpnORBU1FnYvO6Uy/7jZzMjq70wEoHWGbsACn+1XEjjRTlDil+Ln6Q0XnDks0nGp
5+CQAL/C8H4z3BXX2TTtNe8MLXm2M4UnTXCRSBDmPsTm+7Zg4S2MumifWFIyd59k
kcWNyLcbEDeW0xtep0ZoPkZGNojp7Z1KcR/WwcCs+ksvH9yn+yyuvrMzkm8X2iXj
fwCCIsWqSkkTa6nJjeQEP+qmcDLnY0+k0ZEfJhJnWtMkkMkfY+yaO+hrTwa08BjS
JZAAOnevXNFv+FDyONbhSbkfsPPfVuWsRW4fNB3gFF17KpTqEowGrLZv+MKfAtsS
XUZSNrgVLiwXXKy/w3eSKp2sN9gZW8gp05RloNW1s+/FrVC7amLOzd+lslQ1e4m7
zOf1KdSzyIjMkzlKzPR/ir4Lm17hLo9MlfVGJL95YgSbP0uj5xau5lKnlZ73JdRn
nDgZqTyipnPGaR2rFHaJqxvNYza+PB+EAblHXjy4wzU2OEqi3WkMMVuFSxs/lgMp
AHBTJ1uJ5Z1IeVIN5kMHWuF982p3mI/NSAXg0TrStYTimST4/FTJF6G0Rk7J9A5n
hgJybRDeoojg6VxPC8bnad6fO5obOND5QeVpMBU90Yo=
`protect end_protected