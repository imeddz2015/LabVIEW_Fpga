`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 1888 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/9huKRhRMtvnNqb3Z+UU7TahEoHV+T8U3P3ufru7l1O
3DlgtZzb9QxCbOjthp9+wDkjygH0eUfDrEl1ovhZG63grgAd/N1nvegdohFYVoZv
KE4b2+TdTuSnLSOMGd/fRfIPjJlqNhcp8J0YJj/uwHEXHglInM4VlAiNb0oRRPLd
ijMOIaRKZFU/mOqMhBaSk2vPs9CcWtJV/jb26hMkCCc5jDeUjoxDd9enWMjiJ3Ty
0TWvIiEqKhP2geBCyO8rFia3M9wQ517tSHpE4auEFLufzitTrNFnbZazmkXnGjcy
ADJcY2ur673I342Me9llNfEhEUEyCLztQQhDH/LCbCkWsIUXDpEf2/gq4OybLwgA
3tH1WS7ZCJqmIdrUd9GcunUHeVmp8dnQ8ylC/lZQPCZSMS3ULkb8Lrem93x6v5oO
WnYJXbvQy8i3VEH/zny8TwTKGGWYA503cIPlOiOJS+HqY0Ga4AvL23Z2udTWMLT2
lz1FUnmSjfJNvqlv5Afahggp4QbJpz7K/xomepei551ERHqSFULE50dZojsp+ip+
KNyJEANgyKSX2nE/WCf1GhBhNE0/8IZR3bzQkarUhVdogmXZ/9RjiPjpkWttflhj
FQ5l6sf1zRR0hWDj1mHD8gO5dFAbTBMRBq+mwLNIBTDyrP0GxEw3gxrCcuHTySuq
gxBd2WB2JPefccGd1PJaPyBefUi+eL/A/yf+WAiqZq8de5MmMC2b4S2IxF+qX7+B
xdCWSXi4zqTNRaTvQzlwo0ne7gCRTraYrlYJWD2c6J5jcoM7+er58E714SvVbUAy
PBcrgiMebRIHij9MDxzuWDQInYxlxgxPrTzkFeDouQCsb+Ht83eLP9THFI0vmgFi
P4ah0CGlNGalAzZ/UBRelo9q8x26sLLzqnqpKb9/3PmicSkdIEIZ3HSeZlqFnOil
vlv529CSw40fyFyAyRQNellVQdKQrz0+Cq1NBtwJ2XL/0qA322LYpZFByBGaywRG
rTY5juMlahymu86W/NbjiELVueN/chk5mmDEinEQlMKsbn0lmFuyfAuK/efvImBn
el8y8Zhy0nSUrXM82XfxIBKPycm+9ZKEbEl6gTQEKI2h/ZY/LuYl7wSO+x3boyc1
Z8a063a7ZaniK9Jr+x0+RMP+DksQ3wP6lIOPmugoxLmGoisNgHqCdScAg4EYaWsN
FzE1CdmuVaSHLZw4KKNxHbMrVL5nbIMxBO+dnxBmiMF7GcN2UR+47Nx3b9ik7QmY
zOXxa5ecR1+O58DHIGI8vKejezqogTo1hT4zVfgdrQGH6LOKgP7mtvtv6W/mtKKs
UJeLeJAPou7Stqgd9orIhAfbdS769N9/YoZsiKziRd1VB20quCx5zblEU9dYqldT
+0eMxzZmy+EdOWx0NsmWUwNdgUegypIXyscXKncrC3Umv9AoMhbEbQ9ATsMK8res
jmQ9a9FcSm6idl1TlaLETs2ClxwxG7iKwRapurdFp9FszAaW2FhEXd9ZJANtpNBZ
6SI2RIM9bT6TktGolecImdqNHPdV+FyEwwWwbfvsYelyMkPKM9P2+nJqJAxZtaMN
aVpj+zEN3YRYsJMY70sw0j9kgpK55sWcFPwctHxqL0b6B2PpOU486NsN/akSJ2DR
zjXjW2ToP4wBP9xiL3sGl5h4lkMNJ1GRcpnrLjVq1JMy6QpwXbhy2tihPUva5JKi
92bdJLb9mkXdWq4uY4aoVOkrL+AIlIjxXJ3KeXed6gc2x2spBv5lmYDckTQGEoH8
E0I5P5CFLXwIXxw/aM9fyxzMKQQLreBfBLFeO6RBdoSNmlZl92LouC2Lo8C3Fz8e
8Cs+XaCPRE0c5I6715v1v6MmqkaqCXJ8Agky33afhnJeHBMmhmFgF9112iMhsnXr
Pt4/H7G/a2Ct1iQlhz8G96jDk1N9CSKoyYIGXgBWe5naChhBG+SwTXJONY4AAb1Q
VqPXhfx4uw1J8gn/zHjy+YOGiysn9HSTNEnO8/1m7QJSYuezgxLPHkikdwwfVtCX
6DmwWVUz+eVtDW56ARvkol4Mstskw5OEnKrmztNRZ+R5x40vTUveohwNL1zwzlW1
HRBIbz0nXkPRS1r2dEyKAkEeR0b8y6Wkb2do3ARfMXsoDXXCMuFJR36I3P5j+Qxg
k653QREsSKd40gFJpUgROrZDNOP6QaCc5r6RtSI8am5uIl0kNVdt9MXCwebOxn9m
bEL29/axTaWSmsMkJWCRwnV2lCs/9S82HFGMKM0QnLThiUfqnxjWxSdniaP/mIwy
LI/g4Ho8C8pXeNk///LFsdkDp2Mz9dVc9EF1va6SrgdjhLpXT5eN6uhIfOg1H2/W
xq66psq9bWVJpjc9cc9EgZM7XWjo9heTxQe0GwCKX3kVjx0BBFXL7al7QxQJdivg
UoZQy9KxGN2ODW8MDzDXq6iFYpS2cFATztH7rHB7USWB/gFrR//XeVIau67BBr3t
jIcilX99Aar79Y4a5Ziw0A==
`protect end_protected