`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 19456 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/9huKRhRMtvnNqb3Z+UU7TahEoHV+T8U3P3ufru7l1O
3DlgtZzb9QxCbOjthp9+wDkjygH0eUfDrEl1ovhZG60ixD9IMnqfMsh2gQTQ4BxX
QpR6osdETy3uneml6t3LFW4QQHsaJbYlVWazL5sKyWXxGX6bCwZ4tJiruHvjnUu6
qvVUery9ASPWM1O2W/OtHIqub6MTc/9LEhawWdsh+ZXvL/0Dj3wA3Qg05ZNwneHE
PQ9ZVpXEzFZJ7NnDtJAaEkS2YlkBPAq9kPUdUBcLP16X7Bp2o22sSlu73xC2J4OC
iDcFzyDGBnoHBSsjqzFdccgH5LNEkF7Wwvplsu/jH3lgvKWhPYhWiMRuEXrxRFQX
9WAjZ5bPs/qR9cvoMEJMFe9JXMp+7gJCHBHPh1GYHIv9D21JnrlAjYfvL1IJ4+ff
ev0DTCa3auo6LZcMU9YJ1AxgZlNTaeGQ4Z21yl6Yx5j8LxVAtUBd+ba49GDn57WL
hzQCEnfjTq8SfgrdS+qShB+Gw3m/O5arZcKXbZUkUMjaYlbx0+2DK/9rPSFbQl1z
xTzL8EX3Ps4XlPJ8rPUSB+OkdTMK28lm+IQTVVxJ0VUCcDcbqeMd4sXR0eQSZra1
2/n4YCzLI5l70CqYOJOUJ6V76EEZX77RyzAv6ck2u4hIzavtEv4tsOVFWakR8gph
HzpXU2uQD7lbjtNzXjwCkml3pM+OsxWvbzR3VfwSfuMD7pelrbfjJpmJADsFiebi
Rizl1uBUHkOx9WLZ9wQTe6sxyVRuK6Omp0qD4dW1butliwOAhFMTeKs0B/NPyqXV
Fl4oE8FwNZYGqok1YW99IMqLfFjpQeuVKjt+flAma21iJnhBNMzFYOsK71bvVj0m
SM5t/bxj9IxC9Ef15TVFAWPHfLfJB3C9wi6mf4Hes0Wxsnz55X7SbMEFji9Ds7LX
KNa2vogOfCB8poEjfoZwF0njLgTqMBwSxeKvkdai3SpzK1MVEisbDzOlj3o9p+13
OCVeLs/NG7nAuImqHsIimmj7t1RmjImMlFbaiGNkOP8UHLUdoTcReLf0/KyEL6oZ
jcSVQMjvNmGNl4Lg+APLZak+fCpVgpVDpA8WsBft9yHMhS/JH1XFEciKgNfcuI6K
oDJS0SdMdiGJgnsPCjwKuGq88XwRu2P8txnBIGy4uXq59Cwy5Ts31Gitt7VcNnna
3KsRqlBaPpGwQJrv+3bYpwrY2fHBBmwWnbtFQfsesgB4nDeUpEMSuvPYR2nlhwEL
fmBFFNz+jxaMj0+4v6/H0b1rufeuUWy6QKpHMnG4G842JP6nTBbmHrEwmnoYv+Jt
E9uPW4c1LR2UsDhl5vLI99/Qwupq4qSstNJI61/dUX3TRGfq7ZgeFtr7yOZX7BzH
7ihezRs4uSDOp0YFxlPKdXtZwzxg3J/uYa6K1tSWvEHHMAwCPwlmvu3RB56BU9rZ
YCPtAl/x7ucvLhb7W6Z6q4ACPtqjociGecaHtfjeJm0I1SHQWL36r5+ctPED4LI/
8rqyGGZ6eYgHwTeTxnAkluxl9ClB48UDprGzLPk8CbxMrUfsPmnKkb1P/MZwCs1n
kXXCgQdrt5lsOuN99O9JuMhbXxMPqNbPX8luWeg6Pj3VV61D830+72nb8yFOZ9CZ
lRoZkVcc0Ui0EVpYQBhSmOppHVazCGYZfpPxFLfUdEmUSln0eyluKjA9PRm/vdgi
3IQkqFFoiMlSYXvRUyhGpSRC8YJ53LFAEGN1PlFlSDrkj+aHa9f8Z1n1E6d3KYPi
34GJuhBfbeWnkpPlTNaOXmJG2C8tPlu4DWscO5fpHdKxxZu1yrKMd266vYy9elVP
r2MFbfteqQeOMSxXjpbmPt6NEUHN8dQUBTBLLyd4olfnj6A1hCgPxm/SRLOOAUmA
CkTkFWlQgaNhrqP0KwKgDeKDfPDJTlZsakPZrKmqcRyIxgLQcj4+bIUfyowxyify
3TH9Tob9WYnxLZiiDbeRPxl4DjNIvuF9zct40bhlTb1Hu4GHhkkxBzrOBVUOFQuA
vFI+FuQBT2QsUrOVW5H7EHXXffG3YuhAsnidqzNUdMX1B5uy9wn7Yu2zw9Lmkb/Y
aPHswFQgy4Whm+LSKDJJWP+tNOq//zmLeReyQJsUR86FrmCYuu2ZGNTKD+f/tuxo
YfAAv4CasPJujyE6to3wMorNqJ5Vcyi8/B1YmJuO0f0b7t3Jk6yW8pBuyyckr+5v
2oa1P2JTiGTfsNongSKz9mBWUXe4w7gVpnuP1SzqscDYpMtAhkYzKbbFayqUPINd
vuddXfyfyFCfx327ggrolhOCIJeEdq6/WOD2WdK53fHFDB6fSouhK6nUCLOpgivs
gJUxKRhDcjcyZkWjJI48UGv6VGb1bNbk2bqJDQmzP4wBoZRvGzgRdHcpL3lxFUiN
sxVhlZ/J4i2weMmt+I6QE5gniwqtEPEpwAQANc5bCvHURHUZ23ryFD4GZm5BBCp/
RS5w3e67F/ZcjRJTUKqt2Qnr50OaWaS6/a5uv2J87xAEfkJKksgQgO4Uc0ht0p80
1qa1BevRb9mgsd+yB7arfR8Uf/sojHluVXLHhWoLiqj80MTV9s4UKBmuL5YVhMrM
bhQRXN7OwHIoQqfJNiVG4FaZrXfFdcbHZUAAgSuEPc67FllfuXy/elzOGGznYLZE
G5JVpA2OapZbV/Nmmt04BJ1MrqQvpXreyYYBmKhi383JGy1FC0W5uNYCy5qvy1I1
DCh0B8xIS+f5Rf0D0xiYrLOg+vE6vv1FfdaeUE7DdZE4eJAN5Rie4c5yWvDHhq6v
SgOetQSBKVvRWganOQnCDaxWiRZUoM27wkfGvmu4JE2pwUBHbhybBGT9LjLIZh3j
8sQ1JtL8yffvtCMBDsnRwND7z31gLPDCNf0SHbUH0BiX6bJseKpgDgk0ttnwFguz
9Z5fxXkaL8T60l4utJ+AKxN7EStjhi+w6JGkZ6HGQiCyLSKyiZbqU4S3U6GdVvSo
zoKDsohcToa2HJ+7+8bKFQikkdR171gLNlGFdNxWPrX1M6eQpjc+3A3tqTcEI3mR
zUI0LQhaHN/TyTvk660+Aw4GjZcuVRBtdYCeL57ZDBzkSc7hoYTnmwzp1fakT9Ci
jeCFrrCFHsmpGO+nWcE2YnjJasjMvC47SbB7tTdQSXsKw7jjrq0C94kKzcdcKpUB
22u3OFBcXZbSHOKon+thRhaQgBRDnIY/eUvF9Zud91QStAXpCXZieVly75eQUn0+
MBGnSQvj8MQXKCtpobfARFoJKToTA1Aq2GwMwZlj2fBDBjVuaSmFzqfXSEzFYwX2
mXIaf1ifrIXCySkRi+icYopy0wiOqR0JaFF6GOIsI9u1SsXQVsMgtAnGf0BCr/lD
GEyR8Bl2L1faiKA5a5SqSRlbvx2SLKXLk7P/i0S7yepIOajguhoN9aOgPoWpht1X
reV+HiPr1VyRMctMIhC+l6n9GqMgS/4k3GuB/MYZnTFm+tT8vVH8vGhzdBuu9vuW
mISQ7A5/ZBlUQTM6VdmEW1NuSLkaws5OoH4DDBadS6hGA1tGp3liGgGn85tM0Esq
yftBEB1IWedZHrp4Uja2zHP7eYh6XDkvJ0PsOXCQSuh67Sn7Xf3pH9lz6LSY0cDu
gWo08gRF0nvmfIm2EHrppbNcJe8mIJGNrB7CjHrAv/Cd1fXY26LLfQi44sdSZYlH
wQB6npZ8ELIFNMrdrj6qfnCelEC67ANSbGLigtk9gBUmHJux0XbqWuK165WFCMtv
jXxC6hOtpy6wu8X1yg1bEdipByZ1/2xXmf9cpioHMzVoZdEDCH2zkDm3CSA5xCRh
cnybenZOnBL59+0864A0/8BKyGYAgiZTdJYHk4h0MF0msBqaebhhXMKvNctj0qHQ
pUo622aBxPVOj78RF7E8CbIjHS2k6/SbPXmIwoEyNrFAZcSjY7H8AsMLYeXnpFS6
5eclTFANAdHm40reugdU5iHI6UXHdVMMmALw4sekXQw306u8IKc1lf8FX29CBNcw
oslGGlsYapVf9iTmschcoGVZJEyjdo1sqeo/Kti1NUWWzgU7SoKnzCojX0Somlf+
pSLLsVwQLFs1kQYZvkCq0la1wYT+bWmPpIdOax2qVlRU5sbbiNl3BvyeR51TNxYI
v20j2HfXyifmJ7fy3uTOCAGlrjKSePvHNMEIx0j9ugRN1gDmmmQLhTn/TGyUS8L2
D9qLAxMvIX2Ksf2i1aValtWal9l4whsUmXUbGjEFqoMV8NnZfxA283tey1nm1o4U
t50rZHb4oTjDV/zpDyIXEhU182ckwbXG+KBGS0IWSeJD9h+OckH8sfnm55nkxxTN
PKoZO4e8IoMd9snHZz69VBpXG/g3zk5TB8d3APeQyrvZPSvx/v3L3jksZix+RqXj
eW+JDiSm4rM62f+m4vCupeuhdbJ8yQAO61ziM2T5VFtm++XtNfTzBA29WvUR9++Q
kCq9jkEmSaVP2ASx85vZSHYD4PMnvaMjTEXtNaprhXlNcU4AUS/V3AW/AwV9IBYk
FqGGzqkFAkN0cle4Gjep/ZstbqZbCpXHBWK6xojq/Jix6DKJh89NJeytfQzyIfB/
KkRhHrJeUWkTSFewA5F+55wU2QuaS7Kh8GwaI0jnCdoO3C6I2IUm5s+c4sMC43XX
yx3AG6duvjaaAMQVDtJRZ/gAu1p533Dv9gsEX35ndlGmvbonZFTHzhTLEeS3QSfE
zH9uk4F0ibxXcKXRFdKVe5xbWxecSKhKkJ7Kg3nMuyXNT7oVoddMsh2MtYMQgGvi
Htur9wvjz6yaiPLHVonKK7iwRY6d+6K9pDJeXgvK5xzGICAwelhUKKAJuRxEawk6
9Y2LeM0UqLBrW5CsA+t7klxRbtQvegxPruE7XTjngCK5/tSKQMhmoAlFtf/Izn26
77Ecn2oemBrN825wyFVcMFojEtaq3s5gnPC+PdzIUc6sd0depu5J1RxCqRaCmQ3s
1lBpgClr0yF7TP9y0UN/JA86A+xvSLLyx6uztyrIwYF7NiEEaMRePeZWAePKzt4u
1pej38VkFVu92qDkJW3BjBKkDD3EE6UkmLfGb71nV6sarJIMm29d31gYoR/GGlqQ
xnZs5vtLxyV/nW9WjNhTV+YRg77btS61vkij/Ra2a5OgQ8flXKWHRFgdMH6O52fu
EdYN+WJfaallD4aOPZvm4d9co1NYnEeuCC6T9eCHAMhdO6SbSscS8vbUwmGckZRO
lbcSzK/79ZjshqgADulZEbizSQ7A3h4J2UtRR7+rsjeIr0g1zQaiX2k6nwGOuIes
PwjQlDwsy5uyhpP8hNvlmDSpsQEPAih82U+eNT7n0Q08MvzKeKbctoWQeX9FAvlU
46ZpO9WR2w5ose7HzuSVXW1etEaKvVvmC/Yi0LTgn9fdE2N/W0h0kl+xihUmCuTL
OEjz4YOcW5SudxDjk9KQATPg7U2A/SINoUEOwCP9Q+mZchG0BHBJbMc69dwY05Hj
ZLLgsERDY2nHF1GKkOAI5kwbSt/P3Ct8PAcIMo7Ys9PUFn/k4YQKKmVzXVaJDymA
0ADtq0afj+giNb3tIUDXhzBPa2fRmyXyf9SWRKk9fdLqYn8O/TxgfT2PcX6VvTKJ
I+wJCyO6dBaQtNwcLdUmNSLPcfAty2EIsjGCyLMoa6THkuIhshb1iEtGBigAtSJ8
3geXibwBfYutycxVrnARkJTgN0VKyINhiibyQ0pfAZ/q5sljOC9i8npsS/FNVmh1
9QCfEWnkDCTNlFR0xMSUcwKVH2Sgf6iseFTSjLV4kfDpOMFnm7EVZG3RtEFxaNlc
qr6Xk9uYYAGAcLCmwQOORSPirR5eS7ZhEuLh2vEBeu0v9RbXruPHKHjdpOzJXFhq
EE/ynDPoGk6ETjrNyR/07sSZbVEDEXqsbaZaKqMpp4vT/rtdrGQtUaIH1obeA0z5
7vtwdOBIyyy6jcjkCpSlkU6AgnVvKz+jjAu/ox8O/VdCpDmUu2B3DJknGmgP2+5P
eW7qHvtCAAfBb9LWNUqY/gaUcvr0yTg128KmUcRbG1yzmGzquwpM/QHBCtZIeDyM
N97PoIo35RnPahBX6NuNBKnTXgaaXhhlpU4iCxcbUoF4MlIlIbxCwIokmgQCj+Li
mFKxJZxJ/WNwIqjYq6cd5mYlYpIWS+QcgOMK1NGgTULrorFN+HoelgR/6OMbEt/9
pJho6WGrp7pGJTORH501xt/dmhCL/45iH5RQqLUtnZ/0gcHFJUGORRgJr8BQvHXU
TtYp9mQ+gqFL/xgAn81I5Tu1Djs92cMfEuizY+KfMzgXdufe49Qye/DxOOMus1TM
pnKTyunAsMjK3GfKp8EIkAk+dsGzFeV69r4jECA3Y0JssmSvfxWKVTEy50+cZbZq
+DySAh1xKt5rrxizQoKgGU5s0x7eR+zT6VA3gaIoE1odAOAkoRDgznsgvcrtxv1p
YgAXeCFKaRLpkYZHh2gwbVpZWVTBRvawJn8cFPZDL5YeI6/BVFfEZYg755A5dVnQ
Jf4/AZGV70BpD9+c8l8sjM5CgZ+KjFB4h7dPvuOBthwpLm3vOxLZoHAJbInpu6UM
xfiycY47yUTMgAOy8w995wxHZ97Ix0dtvLKtpXVa70O6MBB91zk0wQz3wAY6ECLG
k3j/VRqqJKAkLzH2OIX3seh12szhQtk7FlmYErutOXJ9a79WxyPMAB1J1TvmsLkm
9LysUP4G5sCC8pj+fkdn/QYra/ds85fqBJ0GpBU8cSvrDBoEvy1buDpOdgCfGi58
3kcf9btWSroGrFA4tGMtRhbrnQTNF7/xpLFCaKdv3kJHtxSvTxDmjuezeKr4DgT/
OiyAbZsMvTIbzVLvmjvFchW/lFdqbLO1y8BG8nNGt6f+Myxfo2h/+bgIaGaTZFJv
fXx6Got8KZkbJWaa0VCm4r2C1WDGk4xXBmWGffu33o8qX+LxLuk+X/yjYmGmQLpL
4GzrQa4Ws3yWu1bBTiaiK7+dsNdIBKxMbxnGj+7F+ScRjQvLw1weVb/YtAN4C2O1
er/Ha1RN5FsPw1fmXUih8FUfofd1T/v5VCI65UatEW8HsR5z0zq89Gh26G0NN8qB
EJsasH2qz5Jl5olqvdBOKcohhY4T/djl86RzPpm24SvOQJKOcigIK5CJaH2pB+PL
GriCyqMKOr9fc+MYlfBpWOv2vK4T/aeTgtI7UeMcEx55XD+c86atAdZBnRx62SRO
/9YhfuDShx7/IAelHD5xTaWhtjnZykDDydG1MxPYbLnBnKhyCch9RjVuvNzJGwee
N57WRfnzP25AcyGJnCjBksu7VF0Bqw6jS+VDVCXtrQVdoHfTmn5XVn85I/6avMpm
ZN8yXMXsJcOLqlES+tX0rbTxNS6Rj8PESy7P3Uq/zgEarZ+KpG+nBoWMeOJ3DEqr
ZslPrnm7brgsNZHwFFDEF618BfVLEYS/iqVcp4feRc/tOu97IQmBN/Pn4MM335Vq
KJox5X7WQo6792I0Canhm6IpQxeOOFIPSc+QCBMJ9dKmpW1cVgW4b+1HOJ4D2a6L
mWuir86koqgH0g0WW9Dvw6wzl4Y1c7iMaVW7VnL8pmpXCKNfReBDR+L4Dc6UnFNO
5EhGsEs0Xys38g3obV/YYiQlLsmiUVdgxLHtC+9vL/v6XV7BBWOFgLRSCFsnooAY
ryyQxr4ElW8k7IioRJhSafJlvv55cYEPPVTeubtH8JMMdarQarKo34RnYvmxuFWg
kwfPoTBczOGyAMZEm3b0WS3Sf82S1hgS8vJlhE0xwIAq0cbLBWDYo9WpRaz6dNEH
M7sq4r5FqwbqVubn20JreLbutC0aqcemKPt32+nPvNrWz9BLVc9MJ5KSMGLz2SvR
f2KYibUemIQxfN7oj15YwVfmNFG46ety/7o+PXVepSusVwMlgm62Ygfw0g6Jg9As
oRzN9OaWS9gOOAayl7fQYuvHbGnwsZurlwh+NEXDCb0vRSDNERg40+eng67+VaTs
X9PQdZUspiIfhxSCxAnlxKRW69w6lGM4OOpXQ1//2JUCouK8bITExSioCIUKo70L
gERzl7GrRZdmG0F5TOnelQbe03XC4lsZ2+pEEtGiuZlPvARuXFP0qePem0ikYx7L
gcdmPUyvuH9obMKC4VgLNKLsOUUrq/pDvSh/UY8kKyj8YIJ7TyIkwVlXba60nm7x
iabJ3iqhkGKp6jkoq7XYCBLpu6e0hy4VuEm3m7fYJ7JXTZp+pSF0h9fGtwYioLJt
6sbp8FCJkDNf9emouTPDT4tYAPIE+0HLtjFyAyDAP3eF5Pzq65rBx+9xe9AvB8xn
HG3D9moLgy5SDlhND3qqHZT/02mN8cRhxTdRt0oSS4OOvwmhO9RGDVVzW7KSMHv5
X1b2t24JW0PAFWtiKUfwoX9YdzeVJw9FIQK/x096+6b+bIHLb1lZ2c28n6szBlXw
ZGKrLJc6Ny92MD3jHuVrkF8B8WuNXiTsj9Kw9c9yZpfoPuiblYm90GYEcQHkkARR
JsEwraKdk7qWjwiMVFC4te2v0GSfga4N0Q6nhxreBrN/tXhB3DHD2x5x1+RBcVrg
O5B/7OPcZJyAoIa8aU7HdT8mkfaCQd5cXS3ydMTqsgBiDnCTxg8dtoubE/n8sYuG
unxD12iU6q0Ls+xF3XHK6Yd7VbHALPl+RW/lRJDH+AbGwntmRIkljwjY2klsPo0M
vfefXCcs8PyGIoQRd6wAMz2EMgUIJa8JIIwH0CeWva/IsupKhDOiWzuP8mFvLAoa
0LTer4UhO5JB5N8ESgjf7pcyGA227irMDTsDmH4Q4AE+Wg9u3n1O6kenk3Naf2W0
SoUHkezPeJYt8u/hT496AhYQ1h+mR+LwJ7paJsh9zzXgKokLFjVMH2SEHSDJOEif
lJNo2lS1ecKQ3BMkzyhG8JMspG/M1f0dcQRBvgFU6DonOQFF+JBNlGpZrKl/9lfo
SiVnCuCSWTs2caiBCWNDpu9DlQssSph3J0eKTWYVcY/0BaD6JpO02E/aFWa8JvZm
1qjHbRFMeKsogsb9w6DjwtiXLwqOBaaeHP6X8Y5T6eztVMX2jdsxlaO/pc1mc4QJ
SGPQghjPqT/3lcNBH03rR5knmTIYbEOnNN/lYz1q0ZH+kF2X1DOcxIO4lptFgseY
Mrnr/l1iJEydE0aaT1g8dbfG1cKQXfEKLXnEV15BhqG60+LxcjvXUijkTLNFSNlv
fCx/24ngmLbTWRl4ak9S4Uyh/uTdcCpPatfj80c9c+TqAWTlX+Ua54afUkRtj7d8
mFvQTF/Wvwu3BDZkW+MqUXFHGPxWYhFKN0ZxZ+xPlrKOkcmOAfltlvL/nFGXCx3K
On2C/Deif3H2AY9X6cO+f6cn5F319L75yJt6cydHfHaWgZ9lXm1NMZ/MSv+GXqPc
UlE33fP6hjsUSfogTdYpJC8fycyayenoOcT9rKQNjypltg1p4H1yDdPfqVV5Mjzw
eaCs9FcYgFkpxLxAma3ZOC2GNYMk+hSmqaC1nI5jkDqKEmBpbNKb7L/VZ+PigX2o
olk9TxNczAJmi3461QLZVQvZqn3HYvFwkXiKgMZUQ0kBFqtj/a2ZawvfAhw8laAw
O+CKp8e01yU9eddUx6e9E8OrXr0JuV3hH1SurM+Hg3s41RFRGH0B8x8ViVNzvMe4
gkqu3HfzbKikESXtllXOskbGrKFmk7xX20gJOMo5Ff0AgL79RI3eGO0rQ9abHHYf
UhUF6u1exYyYAvPMlDbRP8HePWQ1sobrPTejqKVrgkdQSewM41hAQd5fZfFa0qwv
JXHMPw9XdMFJMNLGuTvqA+Tsa73acikxFtLU+QFoEGUOQes4cNL99wCIk81JcAQ/
LbqXvctPrD5MaSeafZQZTwftwP5ND5VLPnJ5EOI2DSZQpLcrw4+TAoPlBYNcJePE
pdo1yyxylbTfdsZvl5sRvMlu2VKre1Po3JebPCMSMJWy4odaSusY2uoP+VOrtA3P
H8Qh9mrj9GK8i/H+iBkbl6k2W9aYhU03yrlnzQe8ZYs/Mo1LTvIEOypB0CA8wt/v
C7fz/hD44lcZYUGPkICNQ65gGe6AlS9dTC1S0KxGE6mg/Bm0rI0kIswIVn6hX9AA
dgdW8bn+4dblEbKudpspTGUUx+tMS7dh3wY/lWuyWB5mVhQPO/fO2GqRiJ1s+ZGr
w/LLB+3do51Fa7hK1jDH7AG1bF6cmYCY+lommAGabLqslqkpMdi44/DwQhEsvEel
Tjc/e53ZYLb4a7XRr11+91FZtX1c6KzhGNnuCnMvQZMmbODYdwtVHX7IUK6Hxl2U
zLFv6mMakWSu+lWddWNAD+uaVYo2cBpq4hcxaONxVPzJoCwHRKPnRmuN8DTDODeA
gRNUaqYN7mMNseS19NxwOFWAmUVCfUnzD/8IYH/F4iY23oh/20TFJKTQ0HoWdWdR
YZt9oXI4wQMb09IoyXRu8mI0E9RTRnAbDoVaTgkiSFDW3e/kIqJuWDQbDjN2ZWAS
81Qn1iUzXL7QR/wsiO5RnS2+aziCljZhDEW52KJGc84qypnsbB3sqfkX59BiBvoZ
ZNyY4d+TPk5iaAFNYWKMgdogeG5MEHOBYhLlnee17dnk2XlL5aJKw/wVJ1YmhStD
Wp8oOnFqoFAtc5sbpPB4VMEeBYsgplkRFkHS5C6evPz+Xd0ZpLFybMX2SrIK3B+m
oPt/w5YAQj9kwnrcIiqEIMgCYdzpQ+VaRwBpdmGnC3iKs/lWD9n0bI8B/+e7/oiH
n39w3IEk4VdCBKb4qIjO/xWIv5gOe6/j9WiSwao+Q7opL+1k+3PWPJt7nk5Z4W5U
B2Z523AXWlt/L4zLmpFIiKEHmTLTGNCU2fTjfe/fNhEwUGBUwRrNhy/LOd7z78i5
6c1kQDjs3C0J0cxGJhnFIEYTJSLSDJSro/dtgorifW3JjpV0/3hk8MJfo5DIyOaK
lLt3ZGEmFqV3X5EExTTePltC8plTpB479UenYKNboyRyNs5gcA+VWOYAJYqJ7IUi
U47cBHvxXgv/v5ji+b0dK6g7R3d3SJBHp1XS93ktEiErJWA7s/mmjmyPBrlv3jrb
aXmaJKL1NhSZWkZ3Ok8FY6ClOVNWp0eEY711XRufnLgJ+j5MskRZqbHEP6xqVE8J
Lr8WxUp4Lm49aygjSlxqF/9EaSe70hW6Cp0UElVtyahcIugeyiOa8bYiladsQT/k
37kykH5uvRrGWZGrgxoY9emzXw+HeOmwZZxUOoqq8HxGr6Tb8kYTrlK31vNefRyS
ERMzRWI4lbp7PFj+iPInGSL6syMMqklrz3L0uHaNv53y6BfVB7MbjxpUtBQ/mciB
alGEOGOLtLYxAVXYSQQtRnWSg3E/awy803FDyco8ssa3oG3diSEu2vWBPnp1YYt5
45zucPWPyupiewoyoYMmhfen9WjJgeO7gH8r2rODe4kuHSYxE7yA9lrdCGE7fQmX
k2VOQEEAo5IeIBkEERrhece59htAJh0P7jcgpgvM2rMwjcm6wK3T5l959kiUyKxB
BMn+/+WlBlRO9W2VN9ounVlajZcbGZ9LWydlSpVdnr1M0sTsYhgQyE8Rn1nhZjbm
pK9qLJlYz2lObwGEmdaI2kyM/iyvIpLWXvUg/RSxQG/cu95QTtBTRFPDObAUmS3H
n1+XWS5dX3i7lnMggQBpbQrhPPOq376sHOw8PloDu7i2qeWst/7z+kdjrBw7BnX7
1fexPjFPK585ZX6W9ayPjZ2a2HIy7WuKhnZd1V0zMyyavOPq0VZzfnM88u5A42SB
ps6tER1fPJCQT1NKHoE5eY8W/y2snK9t97Xdstk7BNWbZvSZvkl4grlxH6WmW4ZI
o8lODYJ03lw/xa9tov7k3MEgpy2sjeMmgA/kC8YVb0M5OGH/wZKPaYOW4ITkUQqf
JqwX/oPCnL3RptrMMEXoWD5RkOr40h3akt+CIE3w8magnh5s9PL11P+K+DSWI6ru
VOS5YKPumKrsr14HfO3oVR5XUhxmZIEPkdoH8zgAUDouZVr2fslQ8try4XezKqI1
xtf9y0qO6mKbKoywxNYwDh7Ncu2kyaVZbApcj4qPLrKexsFlhIzY6g+WGa30kcQz
Oi8nhTie9wX1mfsExbwUcqsnW1B74+hKOujjpIjKr6KfsMepzePaTEq3jd9zPPgm
CojfOphPVmb84Kj6DQJvY396yt0Qxaft3EZcNXkmpA1GGCtfPW39sfqav+HfHz8n
0XRZy3050eOEipP950btsJ5ys81lEQOVR65hlNTxA4CcanCS40a5fOBY1RR97pPM
qG4TcxaTVP6fs/Uvcx/giAcZSJFphxuUgFrVl1iX9Hv6VVaBaVaewiWp7O2VkIc8
JM94IMTZb+J2CSYXpEdkd6cCHAo/UhRdTC/F5xDgL1BkfM0gzeJ/CdcpSLV4aRNn
LeVyOtNja84h9csPwMq9feXrhpaULTi+0ZayuqSKhyBeS0HgUp1ZBhMVS8dmLLOQ
EzZd4Dk6rF1iTEIkohweClYolh5tgy9cLPi00ZBmEH9jTkco0IRMKWZ3LP8Uq8F4
XhDEE6Gzf2nxZgGwepPzLWmGigDwZ59mMT36NVJKbQLTtUbqaRszEos1uWJT1uFi
04OTnYJ4FJX3RzFuxi6obtsatylXLxS9HmPBKmBRB0pwuH3RMH6JyIFy1ek7QUSr
p2PxzPCZGowQ75K3WGAcG2tHP6/D1aROtncDkBUnw8HaV9lEIvsblrMqsm/XYdsP
rLj7k/ukmitH9OeE7u3YYD8f07zHQ6cEH9gtakij9xZzwti+peWOB00dbPw26X4+
+f2EvA/JYDoIFGMVJxPns+lJasG7RL4HEfPHGVLIdCuG6EGFYjbEng/nb09sxwtg
+24k1L1h73uUIh+9zCr+ZdHMmjdB5VREYoAoG8lgkA4OmVWroGjhDqYkMukDL2jo
BoN7panCC7CPC6Gcl6M1KY7quOJDkZ6uTJTsZ15VbRlVzttQBKJHs7+zcaV/dJAE
oSwf6Ogv0nWPUS2EfgZv6QJQAB4voofcC2i0sJyHDxC83LfKa5Lv2Mo1LG5+hv6S
sGJDGBsWnAADJtI8KMn5IN5WvGDD+5PLQu/o4ptzVKNXoacsjEX6VjTFKDxj4xmB
Cce2FOTBWxyj69XSgrK+t6V5sAITAByuZmjRac68YfMnEVk9VxL+F7qDz5WZr6sd
nMuokEQUee5HxSlqgS1saQlyUNxxBr/DFfx7M9N8w1Yr5Q4gVWu2fOhe8FFFjkXm
s1Q1l3TKr8gbKL8BEO7AwEEoNer7W8tOdoSJqI8MQd0ZB/z/GOd2QzIqGK0ml1/u
g18tmkC4TDPYhSPZ4QIhQyAutdQlOGv+DHLJcZhOkOrkK4WL1y1+W8li2O4v0PgP
x4ehUuhlLcQ2vRlaReahUIf7BI98mfeBCzDNj3J/7lNklPzYJlJs52GAvvmzPJOp
MBefACW6PfY3WjR/EzprdSWo4UjhsL2MmXkYkJODHhAcLHBdNjgk/b2kVdm2/yvX
hkjMhV4w8hRr/bPSzNEQ/M2Q/d18dJL15C2mmAxAl7mBqlIxr/ANC+4KchSf9jU5
jd1EpDYJW98okZgQAcQaUcpcE/smiVJHmdy+MMsxNFCm3OCR3/chvjBDsWsafbEE
cxlAgj0Yw49pZaVMDo2Abw9zE1MJNO+FsV+tZQoYOKqB0EFqK2z6zMulN6Pbtc0V
MuLEZjBWIu6jSNx1UZd/zfR2PjVct+J3VmWlV6v+wAaSyGVJBsp2rAbrOpixsy7L
Jh9wsX0A2KWBGwQAjJrrH9ORtoeQCSs0FsvrUvr9NviKIihb3FG0cth23dwxlL6i
PxQIi/djYxboAFXIfJ3EFaNETYMOQRBHiLAaB4bbpEgLD+1rtesNrQNCZO4R78vq
omne0/K/dsu+qs6smPJ/K+wY88SKAZVb1pnRBoIe5Xt/WO5QajTyEcHdXC2eldsr
QjKV9QM4kp3QskKN10LE5JPRjHhNySJMtyGuY18r6TpnV12vsTN+7GfR5M0415rS
7D3pAK/TAZDswELZFEHc8ncEnEkiul8jOKnkOGX4OtdJpCbBKAdABKbOBaez1o3N
gszdrO2GqM5AjnRxfCZU6U9QVABgARCY5yvfMBqtABfIX0SySc3FWpG+FZP+TLmB
M0QR7SqpvdGHMopa/zVJ0Vji1BbPqUhfUCkrBL6O9aX2AOHJEMei232GuGxTrAVU
Xuk35fDxNti1XWVOpL770dGBR2QJaWiU6BvQxXgBc+xgAertvzhHH1ZAn4GV2eXl
mXRUKWQeWxzs0Q3J2qd7xZuaqORIAo/f/M99NZvK4JYsJhfmIhXO+VbLGdjEKkpV
fGxWhVe6gdqyMLHRem5FCGmRbEFag2rs0DfMPEmxR/BoKuVGKL4txcaONHpMPR00
W8DFUn7ZNDHs2zayf1xP+JSeePItbRBrlywMfNgveJ9ADxMjWQlfr9aGiIpgySbe
wKtWHHeJwFhkj5NuihNJfA53VjRz6wB39EqHbjbBTTWPVV45Xgpxkvg5FmbcQ76z
jmBsw+PqQ0fzKiSZ5/Vj2O7/NwHEDDhjhUXmdtwyUVrHfm0LMySwNhjg3LvclhrE
r5a3i3T2a3jC5wkAEkFPRJDW1/OuZPbvb1Cget5PZWy2z3AI3OjejAbO2ijXotju
mGVYD9CtHS1QG8Hd6UHBAef/N3DusSzqT+Rsc2HG3pg+SDyGVj5DY/ohKjbFVPbm
G3iYlpYZi2kKQjSXacwT7nmdkT//EkhNDSITvky3OYHO9VfQTD4lGkoi2Ropzdsv
z/hq/dB5jqjl+TBLm+/jflPxRsud2nNm33XMB4pQsNW1b8FmmOij3sWElMGXpVC1
c2/DIi43ECSXUtxyCjr1exTwBWNs5ZIbS7J2pQZ/VS8hmB23CpBU3KSeDoNLWyn/
EX8P6TsYXkiQj2T5qXDrIS3CbVzDC9iJ2mNFriWocRfgaBFv5kYcYqres1KoveUc
8RcXt/hha79CxxaOWjs4hf/Akr9Falqw7MG6+exuiRaqyubMFdaBbsYYQQv6vhBX
IIldpgdk1WutOTLeCEuaXpwD/11aEfV2fmjy8c0POtYg6UFx9ny7dDeTaroYYxz8
v0T3WHqCml+T7gnHq0qDJVc8575N8PwmI+yr8E007VqnRQW2oeJESX9oqoOG9p5c
J2PqecBxGcgqjmgqABskYgZ7OSCCsT0A0FWQstX7Z3NWoW5MRzIz5ruc0NDkYEbf
qEmqULGMdjLhPq9+sNCfrbM1ekmwk9PVXwFOSElRJ8nGP0k+KVtxu2S3sgpoHBAP
giWaIKdGkSuqtc6t9kXBO+aASGDLKWJX0kmxAy7ANVYwgXgWD4aOca0DLs6CIbKI
Pg4kxSRoyRO/EYHMpKEpXdVeXAIGSUOH02zKUEt72Zo3eYTOgG2zTUjOs3uVitiD
IYVXavvK7QNm4EklG1WWZ9OJl3rkQf0679WvpsyonF4MYpxzlYADvFpPklg6uhZJ
yIL7ruI7cx0o+u3JnhvjVJKCgQmH1tWd8lipD/y9RuQ/4JUgVTeLEF3jtWREq50e
qZsBL4mNkbgiXnTjEtsQwlkITW+e1Slk2tzHwe/xPMIXdHwHGYrfOYEpNkSwlaqW
F8XaVxdnM0u+5Oebpqn+0KowfyKfaOT5E4wCsgHrSOOsS7RO/4rGbWQ2Zku4j2NG
2dgzoO+a1utyMIJZRn74Pogsv06tVwC7bj4EXUEllTAM8GA1ovdSO0G5l9RXfmis
X8LaJ0lifgYjPLgtH94xUAiRK4/xScCXe9iaxqGxNKKIqOemB4ZoRODd9Hu6+fD3
qf/WbrUpbdiErnrGqsy41gCdxv3xjwAe5NmVPQdSSHxRjt04SGtaGy4Yl6pIFbG9
7810MN/KpYuuijp/e/SX1gjVQMCCmTVN268qm8KNyGZk3OAZ2AmgyoYQwJTUoiyH
w8ELOKphkBcwNcvm5//P98adHx+3RYIR7MPFn++sSG4u9SEs54pSKNqmjPH02W+b
MysXnym6kKszgyN5Ygn/DmCr4m2oC4Fh7LY/WhFQ8jKvj7HQqdt/0Uxl4qJEMnO+
PkY4yD6OX9zX6f1j4mqD5SRAHLGYtKu80KpiwHrzjS+144FBBPafiTPr14evYSbe
G7kPWqeN92USYXYxX0Oy/LwftuXYEQ0n7coA8OPC2OOqwtICyxd7EXsL15cKa5/V
INHB5C1X/6k2sLD1FSqh/7gpA0p5WJVit81gCF9Wl2B0cphIPUSdberzRYY8OMMY
R12OxdZtDpl/X3lG867Bu2zxaR0wQFF2IdSI/NFXznw4+X2WKfkx48CkTI5t6itD
YCsdplCI2AGY7TcaEwUucIcUY+ytwAmg43uBxxsXS+Gr0nZxuwIT3T43uGHxO4tc
Sexj5clt28ycRX7saVP4+z/H7GOFHI276rFso1PS2wwkTgP5A4lfIhS007lm050Y
94ZbQnEjnCO0zaGbN3HbRZZuwlrNOXWldU8APp9vxWn9q3prQOSPfQsQJUWeJZSl
JMgE6ritsaw0xLblQ6vDQNldmR96ueLtTOVC+mibRfnZN/6Wv79nG5/cr5R0f63c
XdxnMpibISwhQkK+EifwO7PtHUtghm1tWNqoWoQKUMoFo4pG0zsBc7qhsBkgsqn+
PWfMJbztwGMR/voDtRrQtIe8BTl9oP9uwe986tAh1Fm6Qeot+rX+FZMYxwhD0wuI
uB5V6R58FeS6ZL2iDqbWrdDmO/9V0Mu6o8b1rAvpr7at44Xd6a9ZrovX+JZIyaFL
VJKAK8Xf1WFZnJCQAhyFJXPeoafYPAcYHuGTRtOkyyjLHau53mRLgMiJlPmXDfH3
76dgkfsN4xCWc59n9n1W4WB/QAyrxKOim7UegtnWE9nrzr7VkfhHLYxZ6bjXFF9Y
iGw705FRbusvVj/mWT/Az4FR0YFPLCXraHB0arOybCpO2KC2kD8w5dB69tkjIoxd
5GGLvlTn/fqLy9nSOHtd8k2ibnnLwYdKVw59KizXFykB5zdYagMdRcAbV+/HThsc
raNkqlYfGvpvIt5+HFqn5wDXtXzrzgtdwRxdyc/8BIjo4+N6hZI2u552OeAkv/WR
A8Scg1gHggBNCPDJ7IPj3fvQjbunp43nhCvaI1JxVf4ASNDUo+TbYmtHB7h+HRTk
3Tgo3uwpfZ7HJlod2PfskzmR8Xibs9GfYhJ2eizavQ0rYIh2/ipoItXkDaRp6jMp
eMr2ziqR1FNObte7q2Qh+Sne/gZZ4tQv9IQob4LbQcAgReUzpTVVX7qE8eVroaNu
jACNuVILh7+euulxZyqNOAeRvllN6ENMf/rJsJsLXkPoWu4k7+aLY0/ItDfGs8pk
OanTWr0B0l9VcG3EUhGbBhYJnLBZuxmosxyunbN5slW0fEUoBlyxoswMCyTKMlcF
DjUN6YRiBkGTY2Fl5In4PMxRFRGIuBGvEHOG1TnEEH5fGiS+WvGLLYBNmKyvyXaa
mIuVn2SLDd1mptcl3D53iTaJ+lgDX02aeNhseBeRI/9oE6xWIFsuzKQJLM/zo/0q
znzBrBATuq9Jt8WNqsBrGNUMk7OxIc6AWttUeb0Khg8D4aUCcY3yFXH2UIZIrf+v
m8XB2BPMtGY3gQfjQsPH8xGqWL+KvLS3WDDFthehPZYkIk1UKGW61EoeR6tvkWbU
GYQLVB5iOTQvzH2s4FTk6quSO7IYVuVhd2Os+VvP9XU0RtW3XD7sTp5cSS769+Z1
ryFdIhhzle4bg/kb9UGJniAo5Nnfb+xl5uZ84p0A13d5rtuMYF47e5AMZQR165Eu
Sr5LD0gRjpbX2vsmP3eHPIOLZxWCaatPCZtetgfZmaLoL40LtcQd/ifFBLAgSbXH
z1JJVx9CZVyD4sAPmZtrxnz6MgIU9VvivO1dOBchnLkb5fq5w/AYQc5kontcy4Dm
JAyvAWBLtSat8u0C/THRHGbDPfz8I6wFsjoagSFbigqs+lK20qvEAkSp82ycJ9VU
EQeKHhDV8fF4wFXCtO7KREVgdiYbClFhMrzBZzpt6qMA8AJVRTcUiKYeHUhxanEY
Ms8CTn2ccuRWl0cCm9BtmyfvF/D3CJlfjxLWNi1LYooQqs/FU00kiazaS5oC1PXu
a84fMwMcK3bwS9KW9AK2Key2prjOfm25dNry1CHM4t0KMTXHCZqcDVSQZd/yMuvZ
quzTQ3YkY/md4pKue8iP27xr6vljwJgD0onSTZTuT+JWfDK938rJjF/yGg474q38
34ezBmmZIeWhEmbHcsfONieNZWj2zK3/Dg/uwq4MNB+BZNjeTI6tUtCqxEmR+Aph
mB3Fomo/0hw1M57iN20HxCjmvrd2tEGHhAJ7imHd1nInOXT1lw8fIsKiCYwPhZc+
F6hI14w0B3iE4EmefFvTM9KWgyqPQYXsGp5wuSlh8KsSVw96pbmhHYYXvwJFYwR2
1fIS6dbE9EybRB2w8LlxJFs58GGD1A1ieWmrGx8UqvkdlSj2CtnTYoA5/6SLuTr2
xQpfp8j4AZ/8QdANKrzmOHebu2Gmtq03fQrZIcYK8LN2rigmEDX5V+9RctqUpNb1
oNwoqmjwdaix1rXlfHsnwtgiPaYeCS+d/vZBNeUdsnI1QjtEoSC7jT2PHm1Tab/T
ep0UEipni+hnX0wOEgIzHAo81fmxiUdc2gdlNhHnGXh1ABzenqbU4kYqq19bsybo
3LyH13tHxYhJEVaCDWp/V627xr3WIDKWx+MHH+6Q+ylu1zVECtASwahaVaS4EHxY
xiEJuoKZgtLdt/Kp2dqJ6gkfoE4JJB2ygghrI6c/63+rShydwxsyP4BPVnZmnSPa
VZAnVWxHG4vrewri4BjtdskunYbWCl778tZmrp0YJNgHWjfPMy1PQbrcN5BAwT2s
7tfb22x8TyWxMih40hLvT6y5BZuFmZuekXEfVAUuCNo/RHg8t2lqb+XmZiIx1H5+
VsbOQcyJSDge8zdsgDYr4Q3z9/J0uihsHHX6p5Rhnp6S3hA4uluuiM5cTiuPraLy
0wYCAQuJzx7dq4wDECf9NLlMgSLUTtETVbUrxA6w+d5OgliyPiIxuuvcM+qtVwEo
bJlfDKgl4QcghjbuK1AUv9OlSU8R+aLc0ptVe/QP4r9K765HSPYpUedM+EPt+Paf
aTgz1ulSOP1p4g8NyY0AYQ8BAqzfzQyh8S+IJGxJSEFTVoKqzE6prCs71dO6m2nF
5q9OcxeSmoF/xPPLVuDHw0fawUnYJPWiR1Vn+V1wjdmGma0T7BoxpIJlyCUHfN8A
Bet9ut6TnD2fjb/d3SuQVawO567eseaUxd1lM8iDnmXZ3PK54sP8JiW+stRnkaT+
oqgsK1cEPfkP2w7f45ewL7T3TboH3IlAG8+oDChC/4Umnj916u+Ew0iE9HvPoxt3
JyT3ULhq9lSLJbZIKRr5PKja1d6gNl/n+0E6ZZ+/pimxCbclCRKO4iJYV/gYQxuW
UofZxtzJbsZIfAcrd18I3DHkJmuJ3SZrMKHzwqlO1C6X48DdlVwvxNh7PJt6yDhI
O7K+qfK2RB9cZfN/x8DfmoEtl0jSKWPVR7AFLoapEFgCodpxih0kzN48/wav5VjA
We8XCkmuggJxv351IscRAvP9FFTdLaAI6+6iS5altAlYQ98JVazABjZHBHA8YDfB
tGs8d6ql2J+mx1qSdqmWqze4B1tBylskLd5eC0Tu/8AggOsR8nr1JazUbuhd2TDn
z5S2mvUeFcagyjdbceVS48gGsl9wpaXoBaiGFH9jSAeNi7S2+SIBj+5AuE70QYW1
l1aegAankOi7zlz3a8gj+PrWqJxv3Xpw7V0zMdZ79IbnPSTiudMw4N6fpCm+VSm9
8f3UI1KSULkcxa0DkVltWbrVPo0wvxBJNHh4vwVCBoYrnrRBON28xEVzxjYGN9+9
wahtOw8xKAvSAlWSeN6K9NhE4YBQh5Xjy8DY8BamOhP/2bUi2GycLQLFmIHTnhUU
shnbXB5DXWnCzk5o+XkwilsObXWr32PdM3BIYoM2qQX81gUU1TGDgTQAsLgxm53r
xX74xwZQ/ZM1iCHRtqt/BypHG+zVVBcc5p4GNbhn4teDH/chjURq+CfdIl5BfedC
ohgDMTYW4G2iw2U1S+QpPm7QrXU38rTQy8XNz2JfLvx7etfBeTtXSBHH26srI7rP
8wdn2V7esTGSajm13OEk0ZCySkTjWfeDA+hFWIOJPMGPltZuGgaSOM6NKYVZWq1x
5iO99Td3AZtWawVmipuvbmOnhB1ZMBNtZzGIShXNFVXmEeIF/m/W2FzOnv7DPokQ
o15PBlN1bLx9/DLk2yeu9UNpHEQon/yhS+BsTaqpxJC5NYq+vh8TP/UcyD5O3qKz
cc+LEFIgaH/C1uBWgeJWt7vUNpLURAqeOEAPvKDBxKvIPusF96JH07xJQg07zKWX
FsxK/lf92syyYb+O0hDGfXOlmJP89ifM62nzK6jGNdHrur3HEuRHb7qDVRtCeoPg
pkhTKyBAoxgK3UqcxbbCvMu1loOe0sGaqIxLZiztL6GM+nIyMsaUAP6jo8l7cQqO
pRI3nNgRhN4F22eTgFe6p13/+P/C2g0nKM0i3KCoYUJX9Kunsd1Dg/NxcWvwiZ7j
WE2IITxv732YUVaTiDmFRWrHlaUaemEs1+WWL3DU4P990rUXuWRwrpcQcBs917yS
GIe4pR3tXnWxR5Rl6qgsSc8S29S+8YbyoK3Q5Mvbr/wLq1OrUB5IQJdLdTKtKM6F
rJRfagzr2biD6Y/Q6ySQMK7dw2DjssrVlN4RPMvT4AvSzdhKL24Iij2cxVpjLHAo
gxgfmKyIIQqK6VFWWE607UEyhjLYzQb3QtyyyygwYjrX1R9yYsfP1lORLUXei2OC
KXlSqyai3CFoaw0I6aNoBAOKzmlXOwyFDCbki8wT+24DZBjb0AeWihmN67n5hHsw
wRFPIJWDNlgUazqPLCLtMic0cJKNBtD3+T74XO5KpbYOPPnNMQMmnCQqCgn77H8L
ZCZ2PHTO6ty8s4d7pZcogYDSad9KGs5i9vOm+wAqS5aO2Pqf4zinxca8UoUaeInt
GwcE9HXKjtvFz0Ks0XuanH8J9KSARN8V4SOMXw1FMpPbha7mgWtWDAT8j0yR8QkI
J6xCXYGNuB8nyW8QqaFEqc9abxe8uBF4Cs/rgo7RoxBKjvsI06EETC7iwJeNvEF7
98wgoDXVlIjeTH70cKo6JPc0QkVCKNoI4jfo1QJuOrd8q/mUcbm6fnsMSs678M1Q
w6W0rgOQPQLkxoxQ3vph8+6MeHJTuQFk6NG3+AmdwHCpsegjd2fJs7QEXTwEA4d5
ML5wK0bH6zVhsXmA64F69GAd0BlAn1ZWPaI2wVFYaXWTcKqYJvZCJ0XSSZYRvcar
eJWuVfd6YpIonWIas3dq1wuwTOzZOXZZDBAmGyHQlh6RMfw+BkJcnNE5mQooi+/v
YftMauOowOa1GYBjUde6SJGjcuFPx0FZCDEPuy3Ms8riRonph9xmhZfQSQuxH6nf
Y81Lur/vJJ7b2EY8iozNCHJFTgdh7vv4woWe2eywzgHEAG0Kz9atlh5Yk48ZC1Il
l30evXJWpBCbzOBHXvr5hrXeH5VoDWmzpXFyZ5wlIqfo+ru73za+QhjUCz0hDeOP
anLkjOiu1GfW+Are8uhepD7894BToiJRWltcSzciOx3Wc0Y01CfqPg7oi8bvdgPz
3UFmOXa4vM350jOCTXDDQ11tEgLyg2PPB6LGSD6kXf0Ddz/WkXHu9hKqRm7m6tvU
vHEItqrwTBAz+H215hq3aa+WZY2yu5I1UT0DbpONpxwmWBVST3Mfhl1Gmag6exuP
b9xYyrFjjQ+zyDsZmhuHontab2SSbASvh0vhnivRxsjitGoMbNLKrB+O/PTYidpx
3AyxOf0F+swOedX+wk9IeqUA8G8/U1uTJCB9XRtFn6i9T+I27Co06rjn1rrPzTJl
lufHiGIXWdt4I8awWZVw5JeP4USWsa0iRtUvBntePFoyv3x0Tc8nTeBlp2eciVcW
pLBSjBE4QW2/bs75IbjneU0psYw90P8YJWPr7tU8gIcRSq6CoS1cCcdG+8P69iYD
tXy18kkbS7UoDX7Ncu9/hNp67DAR/DhntbNpCUPvu1gsneivAj3WmE+ueIfBBmQH
M3Q9AyOANS7yfrHZs8bDrGPdopgkn2t2rUKU79g8DwPw6HT3eUJWduxyi48tdtoZ
beroEmkIIj0dnf8YKHcd9i4g6sgVPUKAx0ICaTXtUBG3swAhaG1x69OGczBmbuXS
IvKpP5bgmeaoHxAnTW+DvBnW3wvAdLlR3ovGrP3rUn0yeLyM11fwOgFVRBOTTOJx
zU9eDxVY+5H7hpBDy2z9aLmdEUlFoai+xv36ndwr2FA+i7iFRYV4HhmYjoWGUGaJ
zL30n8oessCDJaX3R/JPIgaTFlZ49HdXt7CjPXlQkQppT83arMGe29ILeREhtM62
FK/D8ZeHZPE/qCBRFxHcJO0D6/D+2H4glpFv7OyKF/AoG7BFwsVqI1/loBUS9j9H
T1Nktgp09o1YWXf7ZXab5Z11KzD8c/nd4EnGT3aOf7jsgftoc+aK5UPZQ+pBH9KV
02WDQG/aGZ5U1upkzd2YCwPaYLHzpdUizZw4r+HT1uXt7eKI7MMoABGZTzndoxvB
/vCbaBSuMwNG+cWEwC9pFUU4i3HcVQfjBvA+OYIXAYcn4dB7yO51xRaelaJMWoOy
fRB/jd+KIacBQsXdBJW0Q+gTwol9tJHJ8BcQefQZ/xwm+pdi1O8AHezT/C53oMpE
k+kOdIMf+vuoJCufSc5R6gwL6H/x7li4Z1nLXUYp3pBwEMmeHbgJVRHH8OQq2TvN
fUXOB8D5ZOYEnnktrdCMpaL/BHBA4MOvGQ1ZeMFV3RLr0RuB7PQEhCArDclYJTgm
nKU3GgU7Ymyno9cKaEf+AIl59Md+7jlZkGD9HvDMoDRO2bHhGsZJxB/VPl28gz06
uULCntwJvMl0HxjJ+rpDQrmXr/yLf4ueonTbfI1sEyH/r+rYDAoMIlOw7MEyJfKw
nV403vHSxwxGsjMcVsoYTWaW5NM6Ay/2Viq1jC4oMHO+O0QwHp00wlyUTbVX7vfz
3r/sN5qFEN+gQ9O2rZ1r0ChSFNG/iZQTfbYM4URomZ7797ivG/kO2uYMb0dGwUmt
TeTYMHWp26uMHLGjHWT9by7/Kj9pFilhOtTjuZBq5UalLMP9xg13Z/arkEmLqjy4
uZfeNFkBeRWiDwmBHbx5463ISn++GZwMmDSVeGonTzviU77BWVUxuN8J/VGcEG2l
st1Za3FZ9v5BRdYZp9KZktkoB9rss0JpMJy7CU4vG5v8nBc4PLB47hzRjgwpyymK
Atl0saD32AVjFIMgD6FRguLzda1WEq/hUGpQz7afZWHzp7Alc9d4IGI+s1HryLjH
uxV5yt9tIp6WOZkBeWlnG/xG8nZX+ThK+h8r0X5JcNnw8lNHUQGOv/zGGI3+XHx3
mQk+rTjuOGPpsMfCXLz+B+MG7mgwIOzZIJqpjjWvxNS+O7RnKhxixwIF4ptLNCIw
lMIqmVubDR67mIQ2k+lTPEnZ6vGJ7rlUa2bkjQ54N+OH6ajqLGo6PnqzVbUGYM7w
DXiC2wWIRSTJXCkPLCgB5wMSM6mn67MxYxSySkya2BpuXE80gA/t64zYqHIGji5E
p8Zmxl/3ULHwOQyA4YSn989gH6q5uljHgD6EpJA/Li9nOuDL1Z4oUNZV+glrTHDp
E7SRmgIoXMTc2Ra7zjoTk0bALd4CgdZQGg2OmnmBt5CeKMpAF48+vTLDCuUHnGm3
HnhsUCnDLzVzAhgnxkzISqDR1BJlKNT4Cjctv6hkUPNwNdvZvx3cf1COoIYue0f7
YAVbmqZpXHc9ZQ+Xw/FIdRTkkZ0SnbaMVXTVrG9S9vA79nInYti35bLGsAiuckpa
JyYoQ68fVCRcbWrK07j84wMcGPOzPx6+/pXSSdTnXnsC0ch78FvBYcTnd5o8m88v
uKMn3ldHVvbexgjLMNZ4MaMYOIgXYG+PPkV4qSEX2s2nfOn3eF9Vu76u/ruDKpyC
3bxLdP+7INepKOqEzYovY/1UD08ZDuMP3Vc9+ZZP9kfb9wkgpXedOhzmOUfCMA2h
V0MC1ibCvJeb1BWnhvLyeMU8cmBp1qaz69CHux9XNSMttrZ64YeHq/M4FgDWNgZF
AlU/RzT/5sMRiQ8zwJRRXTC8RioNsPhnq5LJVCmFIkyJFUqJ2AvArs8CbUp/Pfqq
2ajzSTYupf8aFy9ots69TH7LPzueWUrma7aHzkqwStXM6pdqnacpgWMwPYmsoeUl
/A+KxE77bSD2aLAvJZ/xym00/Kg3lyI8cdjN7LC+s5mr112eNyKQJFyzR7cBwe0i
iX1yC6UuqQ7xI2vYFHBrb1pMYGF+WCOcchTA/Ep5ixCIDYk+8YdGwjRfnXjO3X2I
9DfaBfg82Ebh5cE0Ljx6+tQsepunJzJ1M0Lty0iJNhQe++omMjwxSZp+8jxiOmmm
lG80F2p9H+xYka6Sm+l0mcRSPC2CFXzFsyOPnyqbvuyf9vTW/sWpCY9sjv2N++QI
ncatXioH1n7mh6TeFu4/EgApPzgU7lekSAIMPd+7x/59ZZ65zpNzN8j7TbAiCGnV
eduUcQaWG8XCh6jqeOcQo1hUIiph4i247rOUvO6W/PC7gaZcBIgGCuhOUTj/PaX2
tiMG5XKxNF8Z0sG38WlcQIu00eqT3aG1NKCeVLQMvnbuUDQLmQUJFfVsCa66L/bT
BKlB3ycQqfVWu/flc/4F+8zHm0+JazHwv/aGo8jNe461FI71e3TCn3evk4r5rBvu
2HPmFTPagS9o0Gv3GaQASvGEtikmkv2Vk/jlz0+o5lE84clX7ieslZjsVTKV6VT7
zagfD7bsh1PK4E7W2slR5UET7Eenc2kEHFzNiKK+JOYDVGr25KPmxSAq6qNVocZR
9eyMFVMUdpuPvFGpjcAePC0498PPrro3HZ8wF8+nTaxqBQXFaMd9QHflncm00l0g
4ipU1YH4KMFmIPIO177avffFlQkJYljMQ/WsZcJI0q3pzY0bA8SRHujRtv9cteDl
+dQjbY+66nXAFAuOq6ogf32MvgQiv6TLgeRtde5gjfXrMe2JQDvs8EHb4KtoSmEz
v8ToSbtuqsil63e6nFKEbD40PWr199/08V4r/6pY9Y8tDUfxKVK9UmFYhF+jFk73
CqRMCeNkD+A9FdG8+pdjZT0nCmxYJv2i+twyF2zYvf4WWpGVufxbBEWmII6wmyPD
dShgcn4fM3tbdVvJHTznqMXGqGHUv/U6vvCn2zDj1VMBvovuszgI6lh3K1lh1UqF
SSEdft0Ey0PUpW5t9PptGkbrGY9dYocvZ0+2eAXuBYitwk8bkTXbWLeX3mOWBLTO
xDTT7maGu/NDiLb8oSzrwHulqZrYriRXK8qjxWJ5x2qp9DlMAF4fBd4j7MPhyW1O
tKYF7/5pTckoKgA4+dZdYCntIR2jexXGPZGeOnVH3q6XF4DlviUON13aAdkloPnj
ir5bvEvvBONAwJr+Dqv785mT3GEpKdfaQUKprxU8jJ9VdqjsKt3S6tvHoFnSvNL3
WeWpKuNRVlBGd8JhaInXOOPlV/YVsorrmiX+6Da7jRiHG7T4dBkzLtjIGdbVOokw
HO9CpWPaq42QA8/Qsmhk4IJiqHlrWqGaWjDtq1yhDMBMLY20Wn3mPDBgCRkQeDEW
7br8D3lFumvz25+VHypraQ2dZsSW2qAVlPf9EKxX/c56kYBQHrieJn8mUV7epfOi
wd5tcbC64beFQxxPcTG9tHt9Ra+TE8yRbNB/tOSJJ5wkkoPzU+IdhFKGVU1NuUUS
YkyVpTtf55xMcW+jIo7i03K05z4+IcajbPAAhjCYxnkh7qEw3YojvmHOJbPfMnph
Re1vr7eHRZ9fcJi0bsmLwg==
`protect end_protected