`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 17696 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/9huKRhRMtvnNqb3Z+UU7TahEoHV+T8U3P3ufru7l1O
3DlgtZzb9QxCbOjthp9+wDkjygH0eUfDrEl1ovhZG61DbJ3DCQMvvM4ie4vgV5Hn
5rMWe15uAcAh6Pqh++3vLFQEnj8BNM6nd9fDuSD+Qz9ncFeR7rB5wiPmtPwZVG2y
SjSeB2LtiB54saPuUiCn95emvyhOtCenO1I6dJdY//gdach0qMaHZwpcMPA2aYIM
sfKfAmR3lMM1kLfBesnzo27YLRBcvSYOjdA8th5VKkQmYcAWt8XXGiKI4T1pMsnH
xTFHgSzHGQ3/ZpeF587hssGPZY6UIoTbWXf5HrnJ6tmPFfivjwQWwSWel98XJ2ga
5ACVhNmAikQF35HliGwa0QsfFHJf++ZwIpHQPqX1FoIX7GA1H68D6Hsc2GjlhXPe
xyrouoysEeULSUJ6j2kWpOmPS1kG7260nOxxLQwZ7TUzoVtzl9JID2MSjy/1Ues+
NBX87rQKAy08kj9oelCqFbB6NJW1RC3FiqtsXiV1v46W28SScHqm3kNwyRFomWaG
K5LilbLP7lEv6cIFFMIuR9JhQlHPS0I3/ym3IPO/7vLoWbXS7Fe9NHYzPXYAmB2I
P19z6diTdIcAHCg01zTsxZrwGnbuLhF6bcYu3V3qt12E2+z7QF//vyAgh9L1ntyR
cRhOBXnImDBjTait8guhwAgiwUPbbKEj8YnGSwmeesLLE8TwQu0x8aEybP4WC1Fi
hwOSS5t2o4+BlcRjKoou14/lGUNCmOkrX7mHQVv3XsuPcFsVWmNgm2TAWSAhbqbm
LKhUu3G9fABlqQBka6spMM30ImFdsMe28JBskU0hYbwaTplOtebtYOW1XLN0p27u
lr3MSY5y6j70P0W7BTFh+734EatZnB9w0U2ZYTKltYo3adY3Lmrxi48zNsmb+n0e
K+BGsWbNgi4f6cgTTKuRXVeC59Em8DcHYQmj6VCWzrnphlsNCgrwBEgH28JXk3A0
mETuq4alEl5aOu5/PJPqfRx3EEfqA+RR1v+q4t5p0xpqo5Wi4Ag6r71f0sz0J6jm
kMPbm+09YP5iXeUDsrc5vJCAzuIr6FyKFwgLmpZwFO/Zo3y8k/F19wmiW2j6xMR/
EMRg11o/0a6ZPX78wiLfUbncK+PMcXZoCPiOnT20KU3Z14ljb2XwynLw9uq/VR/0
z6rpBX9HocwauEckzQ5GNYBCF5BNjrUhkXHQpauGh6DdCVOLXypo9SSsQHrjWeD6
wMkZuBcMDOZD9JLCd44s8/pxFDF/u+70cdKhB0FXNf6qRBYbLYP+rF6ju4fTf3um
/lGj4vO70MqWz2u036Wn2tw0tCWNwwGMqmcmCGlHsMXXabOoCfueIifnYxeFrXV+
d8BQlHdl6VxJ/uPTQQEKeTqmwJ8GaW7xzkS3MJe47CoRkXFgM2b4OGGl+wSgxoet
seIXHE+73gYg2dM/XO5+/uzG1VdX5F3AwKbXl4UiXDLKG9CEROfqOrE6piFCV6/P
wCvC6OdnvVHg8tvKERSG6NXRtl8OT/1LvfJXGTwrKS+Gn45m7NWzzCNAB/otKZ4+
kbLz3UdINfJ6mSQX89gZuEGCHdjorJEHTzSBQW0ZGlXamBoskm5uL+GG9QAcP2PV
PeEo7r/WShl+EocODeRPZrd12kqfWM24YRPMTJN0f6rryONNDU4zXAmLNFpJ0QAo
4IlQIf7n4EfRie5nYlVkAxXh9bXtPiFWZbdui3WdoBswC0OVGsNNBbowa72vg3Xn
anPRQcnwZ6aITj6ugR0hgzpuieJyxqDD0zOd3mZYgYKA2Kwtb/+PrcT9Oqug8v2G
ZMJekhxLVSeoenEJCtFlPH95ATtr3DdIsxlx76wy/FOeyA6cmfbFl1GYMzw7ETLI
0YsGx5TYMm6ddzX2LS1DChZPuJoR+J00tBU4qvhK0IayreuiHQFQqwlbSLV2R4YW
4PYtGg6l73zqvUgw/l5ii6GXrFK4tLSzKRHb8+jq2dVTCGArrzXC0GZ0PCNZVtxU
xhhoYG18/4rdSZGRBrb0Ibb8E73Vzsm1fH/p0g2CELrDGdNmtx/WDOp/JQuDRebC
ZAOExvn2A02Wxru+OwxejhVLpnvKKw0g1IRE7yUjFWVvy3b/aYw+YvtZtsqzhnWW
l2mejsIoaDMFk+Vu3CUDOIBdhoUeIVtLzvnrmlhAeOJ285TT/IOqcWj6igfohoJR
eIPhEvFww4gV/MS899qmjCMjOMywlpHP/lr9+a5vlxqa+1qSyVLqLjs3C5E3FKJt
fqqJdsyCKMMODSaQHop9/cAhAMljeC0nuOVzD+kJK7fT15NVI0PCquy+nQ/PuUP6
BkRlkhSE0V8rljeGclB1lwiF3aAJ5qn2/2zXw+7x7wtuJJdo6EEvCJwzThCZ+mKC
tN6UAS6DRatarhxw4mYxz7amykTAsX5Y3+Gi0kgu1fvF+Vgack5NsYFqSsBg2pGm
TogksgCZ4abAi1O01YQ+8oIxujy5b8aJ6OinCSTM/Xq1AoKfJxiDPfdq2FTiPLK6
ZQrf+Chj89dfbjP1QaY74SG/v/mMCYpcI9ucspX6lLlaNL21Uca425m6Z4m/+ZEM
HFLFO8XHs2V8gY54iv3dnRG08dxR/fmKruuSHAw5X70Ti6jT9olFYMfrvLw3vIg5
DwSWOAcu+9KPuURIaO42jnN4iPJ0e5/Tv8TJFPxogzKjbgE3ax5cm3KMEgn9iQNN
dLbJA0XYlI6LYCjvz+Ku/mGgPGYNyEs6ZraZCnzh2/zz90GSOVbDppt/N3OCPJ84
aL9nuvIlKXH2dU3Md8yb1hmJNkFRDfs9jcN2cw7OC+36MZ4zC/pzH9qYnEwJJovW
KTdBRnayEvb57Q+D2k51bhxrgrw1/Vh9Y8oeQTXM2WtV8/jYu+p+VcmAsBgnr1h3
W52HDmty5bQmpjCIgsr+dt4rooIOvdQVKYm5M/dSMEkOkKrbYbXQjXCOZ67mfIca
oioD8JEthygsFJohYg+hniSnGpY+irj4pgYohyOxxEo9oqLNqNVRyDQ8VD7B+OD1
pHjGTCL9YMFG09jQ83Snt5wAaXLIwCQnLpoCbfNTYeHcXN/mFWiF/L48Qx4VQ7qb
faKtyLKdMVswxiK1FgHTH6v4e/2YbZMK7bHfQ6+wFMuSjnsnbsGHBSo2wH59jTSy
Cm++bZhyo+A7Ub/1q1cBsUrZ3b3bVi0bexgSHarrg8+ZWxa4anxOjAhMTBTEIncJ
kY/tX6zqAejco8LltAzqZUOUdsDhb9gSofid3lEBjwOssRaj10NDPsV/TSvlXtfK
8/94EctF2d3mAXnmhVPcp+zOrijFmxu3VluseDZSaizmwvs3xd8TJPEGHZjNIbxP
xnu2H81H1fEuefTG9OwTVpczhYwnRBUexqqPlCYx3W1/NU5TQEKMFqynACJYfblV
SMGmOP8shPQ35eARL6kh83OVjYjRhcGw3bKUSmMkHYwI/Z2Zb/Xy8dJDJXKZaa7D
20j/l3X3QBc1ZRCZN9rFAGN5fQg8erUXrbKpBJ5dOxw13s4hpPTyktIexjNkLgzC
0i8nWsG0RFyjjsusu+7SJZH7Xpe0+XOO+1N+JvxiD1fiy145VQHrD6O4K/ysNiBl
tNN3H7EIhX5Nz0SxjWuMPkY4IDpKeav7I8RlOqMfRh8glWQRS9sOO1dFJsc+dERp
j0IVdomjh3WpR4GerYZiA3dSfcXZmNGeSafGngfGsha6i4DRXV/ZRGYbrljle/2/
gPd1zcyhfxtsxiuSug6Pkm1wCDv1A5IRjRaR42/FSbBNSgVc6JgLPdw/EE91uzeG
SNKL4hN66HzDC22NKDljyzrv2g0hzQTrbNMLShg/iAJJJKoU0kIaceUqzEdxJtuV
egOSDm/L+OWOJpwioCr3jEQT0HVjcRRkyFM5pAuv672O/VxM7vdx34WYugqHDOFp
N3SzUaaLz9vcvt/ylRMyG/8ei+T7kf5MJ0W8AR9DO1ETDSwERr63DLC2V3Mh1CvU
YgAPAaRbFv0asIS8QfWLSgESudUsNdPvp6ipGdktUyO1Xk6vM0VXwFvUqnq5RSa+
xMZlJkb+lagx2T0aTJYJD1JwEiC4oLPtyIK9ikbN/sQDYrXC0gtlrDhyzmH6kkmX
EoyDHMJcKSQD9cEyPpHEe7aa35eu1o8IPANgzMTMd2vX6uHaekMK14jchJPy+cc5
YdR+NpI2/sUgGSdPTcoOlBsRwWrkBK/0qtRtgsIXMtoAOvTavo30Jk4CX9Cy8whR
ZoMJ7B035FtHl6Cb6V6t4xAtRGgTKRI4f62Jtu2sN/K8f9X7vcL0CFEfnj7jzuTb
k+JZMNRbqd/4q1f5BfMVNQqo3CaIVfzj81cIh1gXV9xXJ2vgjFMgZukyJgdVdykz
z9O8X5eDt8I154wkuCQPEnV6Cn9/ASR8RcZv+MvfRVwTtKBOpHHmNRSo8y8LxZqv
KrMr4rcfQExx7k827M4RimxGeTNBGn5GMgLhRRbJqYCpx7KpTYe1cUdMzbkbM+tq
xFBTPpSVD8HRn+6b/z2SXlXUrOgZ5V/x2X84womIpoBOM8MOG8VQoI11zueNVvxp
IHV2lfnYwmQxvpJiakzfNtjzIUm9BMGauPhTK/dQYfu0oL/KeCT8mAiKzsZ8wzq8
6I/5gfbslO4yyXkrI2f82iijiAdhz6TF5oq6CD1FkBO8mlHFCRI9lJwB9IokAYPS
XMW3/UXpoz1Bm1jl6jsX7Wws2XRRubf/YWHk3kEuT17o2fLu8UQ56jIL8k3eWOtG
se/qQrOY9jAnbIzbOZ6oVzkd7ZfhgWqPBam+QHSpXjaAEDBKY25+s58Qg7oas3ND
anrlU+9NWKsG9ztm/+s7mNbfG4bw9j9Ywf2LjNE72PkUKHn6dqeC/kUSalbOlGhz
xk5olnmEq9H+ZXCTWRmy1go0zw1MzI0rMH5WzKGFTm5K73J6WgbGAzEt2eSEb7RO
yFlXWH68WzKpY56v1D9lR87pYKByA+iwbcDTOU+nHF+qazKXSylunN/umQGVJjFV
MQVsv61TxjQBLtvf+Qsf/KUkxm7zNH9XEaklUTqXMFBX1zzStQS6yw+TFrU4XSAe
rxs42WJzWHALAa21PxeIjr/ICijSLUuMQ3nSvnibSZFK1uN1KQ1ViT3jXsAiHmtP
DiUgEip58msshSlXt94NX3lLS61HES+vgMv3tvgRbUxbQe7d45pk+Tqg1c97iM3/
09PTg9FbVxMrU4g6ExdR0RNytcwszQd/qV0tuaZtHqRMTQGwtc4d/wRL4SN/6OfE
k9JZspAhiFQbfsahOHieCrcvT0T4zWG6Og9pvibs+23ydKpj7sm5w2VKq7zWzC3M
KP939oIFcnKQMmS/9E3xx84sczCWKfjqoBvQMLRXy9f5ZfQfyg0FGwUHd/IB0eZN
HFDMDce7Ki/d8sK/R3MRNYdbGF73WrN3OVAy1zV/8YKBNoLtFydNZB2fKyT29ifU
Ht5I+RJd3Brx/eYbR4OprbpOsPLhXq6FCmPD1R+8tqKIDD+F7IxTBTG5G1V2oXLm
8v+uQo4EPutQ9rUBU4yrS2tid/Eve/90MUnkyJXn6C3HYEflFb/+xFlBQ7s1Yyfm
hsbLH5WJdrKu3GfKY04wM7HNtUfhgFX98GVxzedRLRn882jjU3FlGIxYo3CFjCNl
RuKDpc3ffYdbHGsg5pL2JyuLFKIWZKDR5/M4b3dxpotC7AmYcnGic1EG56hMxDUP
EB34NFVwqooPrL1lzSjNJpZmr5rNK+1Fac2btKCAvaQ+zAmYMIzkb/lAuOl8QIh3
Qx2FcWYlvLHjbpVldn7ol3Xskc+8hN+WBeCJKWF3A+HWXZfh5AedZGfwEj0IRvG1
DSkKM0tBl7txNBWdzNZp/RC4ysPYRzbWZFF5VUm1vSLP2kmHI8nfw2QfMQmf3bKh
DoPJ45tbijLPXX7dET5myeCfBe8XAHaB5S+AwhV8GsnFQLLcIZZTUuZ5y/MH3wHk
mf/cmbaxs7xT+8DcXiR00I3BTmCuNGRVVHi3mPUJgCkX2vuwoGPa0Duvyg+Ng+Wp
GltEm5yb9ilCI/6vhC6MGkhes7c3A9dO4zpmzFR3Fv7yF9jHZLm9Mml4GmQZ1DXr
sneIQO6KPzmA+SdC1Sct2EO6AMW82ZhmoL6TRogZPHFLq2vZGz13NJ7iCJ2uHe5n
QwRHZ2Z4XUyzmyCdCeFpBSH0RLeN0fo6pqIadeDQkxsirvtYVnztjwE8qtcszTJI
0h8fnZ6GitoOK/eDkZURHd8IBMYehqMlXPnNy7Fhfnokl02dzYNpyVIUrsPBJ/1h
NJjByl7JRqOY99VhnllUeeesxug5Y4LaK5WEGnnp3bTv7dsLZOyDpjEdsDDQGPpp
ex1DYry9WyBOEkuaqkAuWh/ohSnDY8rHVO1o34IOOE4bd4SFqFnmrNZYBmfmoobf
dw/BuZ+tTOC6JTqyELGurdiOehlJ4Xl8L+zmG6SaU+haMn+1nldGxL9J26e4a+qG
d+3fusSirYCcOxHvPo3J+wjMge851SCYr/Fx2xZFMlavSMpoE1s53NssaysG7RAz
4uEiwNv03GRtw/91phEXm4v772EFtnfn0w8xEOoZyOfF24y3FER7hwARIGvQIBeC
yBtR6V2YWHGgOQVxnvBRHg04IlYDO53tDW+6WCDNt14jeduAM8/gQlDkprFcU/xF
XKDgJh6SEXoHgW/yw3mI149giIDgnZG5YMvfIXN0r0RT4azGP44zM5jymY8YV05H
Cy3fGqgygwpWYP93uYgM8DOdUMPrJRnJj6gfpb3rZRHBvsr29FgRwRz81Xigb/bq
8fhVG3dR+l2R0419cilLGuhVXW8oGkrFNvVW0LR6KY/qJqbqIMH/Vn/9T2jP7I0B
RzR1x+PIAcGQPl7FhKtXG4hSPwXs9qnUlGQK5a9iEI2P2Z7xZuZohZLhm8DZ1YF5
dZCebJxyW8e/gqpIzZtKThIKqCuW+PNJIHR/svHPMuRCJYeJghpnoVNBLIpje0p3
kEDgBBUY1C2YC1UHI9C+pLuNPwCU+Ekz5yWxjXLqe5gmcyvuuIA5csFIh7jDydm2
BQMtqXLe4tRQeaab0G7SX+J2kg28oJ0y19IedFKaA9CFTwB/5xxPyTFzrZyIFUQP
/9jBo/8pxGhypYKJgDSbWJnDqEh/NpZK7bK1Wf0THojy/WLUlSL/A+q9H8q50Gbe
/oFjk6nbBzs3ayLuWX2jPTtvCjPJnw+1DwXJJ0gIcvwh52R3Kzi9lY+6AtQH65+X
WqkLCMfe+am0mqvyGMPp+5ZHS4fCni1ZVGGXPCfpO90Anh9v5LnRThE07uAwdNYL
bYNOC5jL9rqN3TupeGrZP1fjxQmEdo8q1MYPxb1wktSY9uFz+7/232D81rNaC157
avsy5+fujkxr5rSa0ZP/Nl80MtpbBezDrshaf6sXY5DqkbHG7E5qq9ZBIwrz2mqQ
KN15RbXB0JBD9HwSGt2STP/ry/RCl02mfesikOEBeKeBAkzhJbRXBx1T579WKJFQ
iiUvqypMp5KLC8zNw/HYNt9HZJVutFL3Fh2iffW8N5Tv7wekxpV4J4IzYIyNNj1G
T4jhzczTyVgZhh5R2PLDVg+9sri2JM4PyHtOLVt9s5lej0KHaUAW2KrwsQJwaeUk
sDLKjO4f0JiXjnRd0l4VyumFbbTTafycgsoEkcn2XyXn9ne8sJvj60b0zLm78KQy
EGuX0WggAXxQ49fRGW3sLEnrrRRrSidUL1AwOfY5Sxearoefl+/6MWL5OJqTqcCT
bcj7uBDwjv+snlfYXOmKsdHJddkW8SZZVf5dgKUG8cqNHWu+sQj472sS8p/9yLhL
cfLhHwEWgReURDvVkc+8g9nnkr6yJO5NNouot6pmihxhl/BmC2DBeWO1d/SKfuCk
TtpKSmBAyx7KP2QjpuVsyB0BvTP74FCVx5f3EPROlHhNbqpGhBNlTmYiWgVahabE
JnhXmQQ2qYXrODk+MtHgMwwC0Vq4YgXS9haOLWNtCT8gyWDXXjMFhpUavli7j/dY
uVsgpQ99FOy89Debli4DMlyG3pOjF1Doqha98ndomTt38ZIBVvEwS9pA8ghw4lML
EHDmRw7ebcmQZTTeZV8Um6a3pyQ/ZpylxJ6MqgSC1tN/fzmS6QriGXJ/fsf/vqBT
iZsF8M2mIVHhFL+Ewb+hh8BDrSUM/pnYu5ezYeGYaw8FG7oifxIijfKRQtK+w/mf
8lqSAAdPZB2OA9h7XTID4WfnP/2lJLAK9zl+QVbfXaKY/HBt9GQe4jJ1T2V6CoCW
sYTss4SaFiMGDaIciFNnCLGBzqy9utfDdyUELqjSjhfX1mza1GUBxscRLNd6Xwu0
zJYAv76t4Fc6QD2G2wAPTk4Cef8KGTg/RKIyP2AYMXJMsntqZFJ9K8apNSDi3KVL
5nGsDRqnltVZ3jAgtWV2mbFPmC63p08Uq8zRbhUT17qSHMIbGR8g9fpQPv9ZjVPg
HLDk68Erdou50zvpgMDa/YQWLVTKTzvbQ/L0RR5TowCb7hWLu8nVJe+SVmzXWQqa
45qh3CYncw5bltgeFVZEyK954k/OY3U7u18YyTQlOAZPBtVTor0/zqeScmXna8vP
n4do2ucNrnpWDACgKoRpdwdrB/A9/mGDwj9rLrBrr6NdFkP7z2osd2YZ2viXXH9E
SzJDFbP5/K2XYvUEkGEOi9kzv5BY1oUOFH33q7tdcdJdr5kSxxAQLvLry/0oBcGN
+aK+PU7hi/AKK5Pm+ME8VVGz27EE0AmAYrFShflgsYimd/mSCi06IsAMD3va0KqG
6g5IVhrJRjWvFBDQy+25Wx6Qfh+PFxucbN3KolG3SK73W74CwdOc2ALv7RSCTfvk
W54iQX70zt81Qykmcnz0Wt13DzEsmNlT878YMsaVuH9fTwi8fvo7ifMsAYX8voBQ
1rTdTGjwhRpGOowz4bXTWNsxbXgSLUn6pRz4VK2r33bQEOwj++FHOvd8/ygT3/l0
G/6QUJtjHL7W4jj6Y5n80Bph2MB5mC5TvLs0wwUm1M30Cg9zislKh7eVDDgH1DvK
ebQ/EeNPHkR4CcJ5H3paA/Tqt1JleW+5Ex6oL6+huk2VSi3JytMKhOfInl36d2zG
wUfSfBAO74gjac39Tj1P77x42PT/h58vfTA3R071QUP4BJYzKvO2rHzHTLjwWCk7
yQ08OFpdpp/QJY3gZfAKiriIWPDqnE/K0qRSqVS3JQxmEX29Ou99bmvhEofhm2ba
kVh51FD/bD/yNeMxFw3Zlkgy2k+IizMWx1bRzvvdI6Lql/wWmxUToGihR8ro6+SD
rbdzM2NJAztQZ0u/HoTFgwpp0vAwIHzDwR9ey6rd66I0mO0BqEaS5XOfGjN0SDU/
2MlwUsHo7Ib/LMR078skB3yuIbPhjE8tpFw6ceN+SUIYy9lbgxFah/F9pB2OsinR
IDboRpoSSPoKGub5APJnrozP1tCjXwRX967pWlbwHoA6/gnDZ0Qxp0dkzqPeVVlg
hIu1fFR4inMth9AqxPQIvkiARmKL/OUTz5B3HwA7jrKgkEfR8rRUwWSN+0ZQ4Vmw
R85IU9aStOsM9nozwM0TwZ/+D3I47bCFUI68Hu1p8vKTH8A/gtFnBjzuZhEMS8HT
LEuC36vroId8hEFrj35Uc67Y0DoZNXl8hiHulWcLZD0UImZ1K5MIZrF8GWAWgr/u
DEvKE5AXzNnUFXhEXnvOecFMxYBclFk59QcPFJfTbXFlmetJYe8n9UUJ11EN9yBC
cDE3EXTateg6Z1nv8U/cMdRko8uA7CjOfqhUu2S6ZhTzrZFT2ge84nwNvBBqp//L
Edc9GYKdLtquMvfDlFHOfBuhCb2h+0QxcHzoOVw1BROnmE7Oxye8+R+eJCpjeHo1
qAdDjwLH3r1Et2I9umqTw6eE367ofv+mIwAjb384OXj0sfbFmRO5mkgM+NSkuTRn
dyXUrkbHOmJZ6y/tGJqKgo/wNePZQWumUebfoqJ4sk62/xg5Dzf31y56pwDPI1Dj
+zPOOP6DTx5yX9wc/cBUXXhA/pPNGSrU3HVgduGO3Ur6B8cTFwYPM4AzjOMOxYB2
sAmiwhMORQGIqODMkpCMJUft0ES+IDuAXAOY8o7p66sYpUk38nWPxE290vrWt3mv
QbgkpgYY9IAk5CQX08hIxi6u1NN5qe4AEOjAVdwjDCc2wmFNxTAlamLW/9W1S/YH
tgXk7BMzXl4hLeHmyUylvnV+PSzzxMeF6u08wE7opSRoyx4Ni6uf2s/EHFM5cQR4
lZmra1sCF8N92+sKZRPxE+tPvhyJ29ELiFTupQVIcs3NV9JJTvan8LZuEkDPLN8B
7T2FXoJgHF7guaLoUUWFLWERfpgqGr3X8UROSw5EU1NP8JOWVCWk75vljmgaMSd2
mr4e5FFcbnRA6Ozp/zyYxy0HC/UyA8svNdA0Xw1yy4J2Yy3ja8dPos//sdSCrZ8e
O6f/yHEo4ro1uxyjg6UM8jIJGLdA9pT0n88qb+0TW+Bo+0cdJisAVwBLYosxxVvm
k3lbjGTuPYtTPKhDW0qXJRENAj+Q16eCUHGZu1XTmd1ZRYnvSLG1PSfEpMRuTrom
8SiO3yUb54E595VwzKrNGDMfB8Hh2ptEzt4gfWSqS4+dkFqOPS3FQY2NlGjgBFh3
+nzmCyu4sC6N/93pzU8tZsldDoSlAgR1G9R2eUIP32iQ472paPq5fOQxyvsewkQ5
rhdV4uTAwhtSjDqDaGzCXyjbGtRsRWjdxKF1ZpR+zCbLubS0gXJCskbIkW0klIif
dSEBjHJ6GkwayYJx9O0yTojCUrsTSpl3+cEcEuGX0jHjYNOxxDDhsx+u5noKEQ+E
t7dJeOE4JWgs5GSS5bNmo0jNcH1Z6Mkq2kDkeRddwT2F8CqE78WIsU1wXXyzXE5o
wHvMBrciNvsBX2fWemeb9c3r5opHaGSKt9n1mhmIU3ccDCKYZO68h7xCpVDfVEfh
Kgy3AEf0PML6AJ7OIhWq6pPmzA5d32OAq7+8lclH/B8ilFCl2UWRwZ8tUy/QNpEa
0mDqAC7PzUHkW2xEesKX2IxN17lECjUC4FyE+KHFKByiKikJ0IusQDvuH/ZkKxj/
vO9b+h23tUxTUIzwc6+zMMQj68bmDkJ9DBtpjyqR0HigFQhmRIOCmo+9u+uOzNQw
Tuj9pZ1JLIqEsMtWnZwGqCyuT6CqtT7hyYIgtQSdR+2OWQqKFMiHj15rs7Te3hjn
SkRfa43m2OcKTA6dNM2Yr6clSllwcb/TuXATSpJzQK6cJ26bpCTvPu3QRHbo+93U
p6rUCBWqpZ7/ON6EN0jofFOplkOYzFF/Rlz45SNY/WJD3sGeCGK/4JALXwo7qRdc
qI9bpFGOsv81U+Ae8KM8bP/8LzaHa8vXfjy9ROV3JV7DUBXpKIsGH0aDvHgKCAlC
Akq431tewPprxOtP5UZgtEa9vHrYCiqsJNVzeODgpJzh9WTPxBdIbrdfaGTtnLfK
bicnPW3mjq6BmR6JuImqELX7nVCytgtIytpF4ImguVYPeNlJzBpOBdcGnRxyghKf
o9TsgrBWKIr/4PMuGBImcc2NESiQDNzYI2zB9QyqAAeLDrrbEUpVlKWeu+EU3Vqy
MAsxcFfkQbdBBTfAmkjGUSbXi4aQYJf2K5JxhjqrQ9GRUqKRiGiDdbMIEgptVLWs
dJsJ1vU2uEP26qHFM/DEIii3ip0xudTutGXZ31mPrDAf3b1pk9krym6DBWgFjSxP
1SU8IIQvpOslH5+vf3mbcJalkYVhP5GA3fdM+kliQjlL4qaXhUMELq7G1E+Xhfwr
RH802IDipjH0Z6qH0xdrYITWpDuWmtKCTWJtjDrnyubuNFjQI06DeRN5LS+Ace5E
NxxfUTi9W/c327xRbL0kgVIvvu+nE2HmNe7/uJ0Co+AxXAuZOlZ4UYSSZHyvF/M5
ph/ERIp4Glbayai/GSK9W8ZgqLjiWHYRT1RafhHrpnJouMAtdyQrn/TPlJr90Z0/
65HV7gAVngJtP1VO6axbXSTQhyJOBAG/EPYeKtVi453CX/CAvhzYW+Uuym0aiPQK
AGeKDDWJpZ3JyaSZapp9P0MP84L2RIqCJkzfxF3sS3kPi+yiJTjo9h62EH51rLNP
RzmVix91haiIe42GQlnyX79CtM+1O3UE26Uxf+Kaw7Een1ovJUkS+NzWFC2PL8iG
7mBFHdwNLG359gQnMGksmfwiwttSIMTVpDmlPd9s2YzccFZuP1Eg4U1DAztF0eni
AeyIJEvLSfG2AImEIlcWevWr204Gnurvso97n8G/7pu0sXQpXS2yYEpyExzaN+rH
4ARJvdYaGcJno7JD0jBmE2glPbn4TjMQhoUxJz4hS39R4UpjzNQyfPIXRnO8zQSL
uRPIiokgao2G1FTXNYVc4D6SKAEBTA4l01lD7JzkixuTtfm1nWqyiwV2L8jgYIdJ
a5XjR5NYAU1rHecfroPmzhvbYrfW4axJWo4LLDnrIteXH8kVc9Of8r4VJVZLicaj
bwDrScadG0H6ALfLZSJH8MHZtwImXgJkzMa2ZTV+ayDWSPnzzuQjXXiXMtXj7RxJ
IjgK2kZaKg/rR7HXTa//uHFyIR145C6q7CZjUi+yNrGoU/7ouppR0F9OoY9Z9B41
JCw6Lc7XuHvIa7UjdZN6m1ryTgrav5TN3QwLSxN6AHxX4EnEIkzMhfaLcNrF47et
VChF5tyxu4J95qlgDH+PO3MJP1/N6uaZYfpjxgxe81EsFwGJMNwZoslswnAQFt0j
WgJzzgUdjoB9FyUIgcZtoNysCO2mZWgONywUpJizdsSZhYDWybutiG76KgnlAHae
Wc+z3r8GDBli12jHHGt98BlidmrxT4k+XOSNrdJaAU7KGSHfE731xquXAXD9HIbB
P7VfeEP3l06OjpW/tcgu/oTqnEEi+9uf3CyyF2niWSXyWhHa2vRN58k6F0SP9bzF
I1KcXfGLuUxVwBxeMvgEODS+BSMVhiN04QCn9QQkRcqOgEy3gJZSw9LoxobhHTua
MdX8CqMrJQHbg27I1QfPBlonmyHW6F6Yb4ONsNlA5O3VSiQtM5agZUR87MrLSN69
FSKDqmQmAwzqWPpova/LUv88YhhoUUiceucSy/PqF/Oj3JDOKSgi9HN39UuMt4Zb
Si8Hs25WuDVl9mnBYjQV1HObbRbJFVXBWvx3py8FNi4LuhFvLFwn93fAQJP6RBWt
RBNV8wYjtxsdyj5NKKp6GXq1l0Ig1PMHc1i1zihgBHTU7COSJN8Bxgn9FeJ3s3cY
B8iiOYVjM1KB3dC75jrFVoABAb9yQx8YYw8ruEQAMLWe9f7Wxknzm1uTkMMK5Am8
0dOz/UaIykdht7gEhZhtfcIusceHihrvUO80qznO1qeDeN/4Z8o3NNJBMGAT02zI
9h+dEhdnaFoNsuSgY973rzX47oPwq1MAxKHmTSG3JKxaVBAZFedQsXtxNnEcxm9I
JdROmcFM1VjxHt7R0CMkBugU2uaWWIxiQjERnGAckDvlwoliaPTqiXz6RQxDWS+v
fW5cg55iRlXvNollYZCZIBh06B5IlcvVIk+uaDV2bcz+/tcq3LERPVns9Lk/gjih
ziXDvKsgi8u7WEoyzAavhwX6SFmWM+njF/dFul4eaq6BQjqBDLlRj9Jju5KC2U+r
KOQqXfGzm5OFVFL/wXFWfyXZOKOf5JLhTvySC40NU0K70RU++jOLtMpoEU8AvFjx
SdM6yP4y3u192G1uxqLasK+FqVysy8/8ic3cv3qbhoOPGnJpIJz0zDW3NrSkJ12+
B4ypCH8GQNpaLyzo1T5j7AJfTa5ldWUAFmMwVMl0h/FnnscE2sP6xF1EdGeXMTS8
30pX9UrJU5tnCB9bHPQVoccf+HiiCvKCsCZe13oBxCV7roTB3vvchBZdqkJA8sEM
sFjutq33hTxtr92Yw5G8VLNZV0itPv3gUAZor9T+hT60OWTISiF8IrxsE0RTssxj
59Sv1pPMpaCrM5uG8GhpvyJ3Vvgyb3u3kbKVIkJy0dndJkwlts7v+Hkmo3XKuKPE
YCGbOxqw3LESZq9BzrYiXyQQOTb+H8wws5Oj+UmIB4kl9F/FS0K11Abn8hKnGT7t
hE8GLX9wj6GjR7b/Sbl6DPaRSSVnJqYPhxPMXN+hPM3OxvFLdcPS4IWPhQEp7MYk
GhOUUCqaJciOO0WXxdCDjxR2UGgiUaRpkKUZuQDoNSXd5y405RdIkiPss1oFQUXM
C13uT9RSxIeav36/yKEk+eiSGATDReiE0Dz884d3k3eQy7sGo9qbStamX2gXhLKk
DB5F+2LZaytTBskkMm1EZ9w7E7VQWgto7WixfeQGDkq4mIBXBJe1+dSrdYA63FQX
fs/2X4w9krQJw8N6JXqX+DfyIiBiSp2oYoITLTPU/y+eLzvU/C+2SV6iNJNLrQ/7
SI610w+SBJ5Bax4lR6aojwC66taa9BMqDvq/AbUGoNZu9khrRT9sIVPZ0oG/LsoK
GPrrTYKnrGJeoulVMbo12lxFfPxOYwUlXGSsqTstxp2SvNxQQvQBjUl+ZrbcLuUR
tSS65q2Ajw7kPEVdcxADYR4J3ssSGQd2zW00yvkLd50BY8vDI0TuRgouF5t5tyDW
bTCY3dCKyFWIPLG+B+ZmIulY/orRsMBX69FFWXx0mFwb17Mb5gc7sq71o8Fxxxoa
AQ2eADY+dGBww8stq9zAH7l8xQYW5lCBFwk5yPxLn8IvYBnm079FXzK+tzLLQYh9
egwfcasJ+tXMcsNV29KD716kiuQvYYiTSWkTDectsKJDBYS8YwUYU38UBklZElRb
kdnomTvInu6Sp+qiIV5pffMdoMCvtgbDMOKxnMKvxDtYV1Zsx9JQtvlCTnJzGrIQ
7XBo2zNyrqa5B0tcJorlb+iWTpSau7dtN+cb8JFdFirqJ26K+r3JwkDk0M+Ot0uJ
Ii0Lvty+UMPVEUtZIhuIp1OeDJzePK0CgqXNkSTSFc+rYMxuSDm/zYevIjyO2pfP
KD4gsz2quOh8wt0TBiWHu8M4vt/Tehg7f4kJIBUEQvv2/qnkTH3bX9flLUOc/Cjb
XBBVyczMB4CgFhKJAhn4/AI3UaHcyryXuLfgw7dwvtOpPrEJrBdpN+FLYZoy4hhX
N9cvlwXKTY6Hxix+Wp7lOi1GaRi4Gg5OOTICUiF6mGIQNzMywYwayOlVinRiA3R/
hnhD07bi32QZwFkCWGK/Au0wCNgoNZTX1TwaOrOX8heNhcNuYy7cMF4EdBoDp+Fy
rNozV+jHyDWUVMGU87jGoN70zhyIaVgij3nicZqz8y60aswUM3aM5srfGfrs8j97
9pqRSrZXBCMTXRlBHsTXq6GgFdjXjCitci15C75d6arKAub1jO/4jKb2oqn1XW7S
hqMfWGBWfARRh/Cf0MT7JPs/0Dd8prB8AYBoY+UbutiNwM3fev888IasYth74ouX
UEkiA4DFWajj6NnVsHjGk2qHjlY8DnJxR4spboImwejavI9jIHQyEMlP6d7DuzrP
KkjHT/g+IZccW4NyZBjQVgzzTyOfkEN788zYktINWysEF0ToMlBU+8XREGJlB2e5
OcVDXq0QS2Va2JmI5rz5ZzmJ+cha8Dg6QwMVD0M+p1+tyaoGohHye9WrA6jQJRNX
dkxHLjx3ayF5yUhc6zN0z4+rkEmdsU76Z1A2vVKzHTzbMiFDptv1+eWroT463rta
JtPtFNpuekUoG8EBJTQ1pliLwC5F/6VYoTNHu1xWtbfjT09NhZVPPpMzYjOWu+dt
zPO4Pe+p9NFR84oRDcL5bFx6Pna6pMNqLchh9skq8lDzHln+jwDn0EKHqmBaN35y
7soeo5jORDEeCudmQiO3gj3iac/lQBI9yHGaBscLR2U1Y0vmeV2Z0FppxJZB/tmt
6i1uLgLKRcSACQh418FgqlyyQSRm4+f+5uacvMcyqkHBwUl8yualkj3K1cHsXfva
ZVcpSWm1mx/hpS2O+RitX7G30ZJwpLlCKnlpzchO/bH6MK378VGSaaiuvB003Dck
nnTuDidMUwqB8keR8awug2GQ374W1lcm1Z9dftw31ufd1GyTXMJ0ExY3Ttps0nRk
LQSt+vSmNxX6oNsVFN3+W1eKC7bPKPm2VMdM3lzy9s9TWI7zVOnODKYwLw+fnLZM
TXF146l2QewvMoMPhiLxIZc0pELNdp/DrI5wew52HJO4y99at9h5o17sYveDShuR
OJa+rhGaQr5609WDxudX3nouoCtaFQ3WfbDORaPrawr5+VnMPqlgHVUfnb+EQRHb
tWIHkswGuCZVb04BQQoIlefv+x6OgwKBMHIj7yMDZryAf5pGN62OsmQ5Z0M9QNW9
rvgQzvh17WZBq6gSUlBSa6FmbcH0KYvMHGPuWZjY8+b1pswVAi6/MqYyPzmkejZz
dBeSH5JNPnAUuPwAYYlNyRj/fbvW93jQnrcROUxY69n7REgAEI1ohyfeJ+Y3VrJz
XZtJGxCX25f0l051UN4wBBKU7Cgk4ny2VTBWdCcuOTcEb10EcDdmky+u06wxriLI
W/q79UHv8ORqJnGi/Ry/zxHj8DcmSUkV3VGja7RrV54JxqqMKJfuLDhZTHaep4PB
8I5r/E8YIbsyFM1UMK97heaoFLRla180q3Hrt4p0x0i0Uixk/cSzSyGvgsPSHk9s
GuBG08j0ew6dZBw18fGtIifO8TpN6iuPDz7tnMLRUUNzAeANpshLSLTFUWZ+Q6R9
YUvsd0fBmWwVxiT7dEuOa8Q9TGHqsn4k3FdhqLdOLHV23fVI817fZ6jFTUDtYWmA
qusONdGid97IOZLXHPTY7Z9gRPbmwCsu4j+xJ3Z4abcGeEKCsOObrL0dBbdK1nsh
O5pa4Z5eX6TCpCG/s29YqMoUZ2ZitwU0kEKr5HP+V7+3x+pOPnkgHXb1z8/XWLHm
YOXjThbgzUJTNwpW4UEBFJZq9bEkQVfH9SVuYuUMTj4tWgtQoH+rzjd2V865zMIp
Iq/Hul64usISx2+yhLjEtITr/BQfjN52c7SK8wdVNp4hpsDEFcm7lrBHViwqSO3b
4cxDUk9XfkKFQQwVKKk1qXW7ued4ntslFPOvuZMSdefoYUVum1lGM+o+YNx0F4jh
doC0aRi3EP+kEwYq2OfPUScpnUoSMGeUOxrGx4PFdEQJmeyC9vagp4LTwaEEnrBt
ofXq6d5XTOvgteA+pOmPJbjw3fwMtIwu9gUyQmztIu3l01OYVuNoSKq60LAjGuXS
Fbyos5FpNzfiUTdxsIPRFX7cbLQO0KTx8jFzGMHBGdUKQKP3AJoupXLM5/YroQhH
kdmsRXmXCQaDL9JdeA2v7I7WuWWfyjB5vneNQMjGeBJImDr9h/pObXi0jQSwmELi
fkBsrvCQFPJc56uWUOHNSL3A8cqXo7pyxn4uJUv/+3Bj2Bln9O9kKBOSakqTvNSt
OietXvZgnP19Mr5Fr1gDvNeiuVquce8+zeDRPT5l+hugkh0WcYhu/lZmRBydJCdq
srJUhK/dpTGREfyxmq4v8GjqTZSOi1TolSaPs/FkZdrTEyPRngaVx3UjleIR5wKw
rQ+gYVOR4R1RtSuBE7wU51CX74wSrx5H4cKf05w5FrUmyrlNbCjOvjuatr2hMJxM
sJKsaTVD7KzaiiqYKKCyNziiSbHzrdbIQG7RyNhsbkgg8GvnEXOPy44ub89tbxPI
ytII77iaBYc7VqT4KNdCsiPe/cU1DHGqNL38YWRBlTwGaENzr6GjR7UfEAwrBDbY
MC+DktR9c8toOW4FJc+BrPuIHbkv9UbEIeMO5Z8Du1KP0lGaTm2GcsqZD19cVJXw
EpGlg+1fKwxdjVPlihkGiJTFiBSy5TpqpiDYnY5l+A4vbdvtBDGbzHA4OiEeXHLK
JHh0cP6whh1kZMEmZqmWVz4wZb12qTg7qHoaitOzYc1Tv5YE/3SUPTj7q83JE1VZ
6fzOkE2OhyyVJXB09QeRU5dnn6zy8Qlj8AMtJjce+DR6zP1v/Sk1sr5JQ/H5pdXw
quqaYnMelWkdyDZfNGqQd295ufPJ1GAStuzS9JNlaUzRXxe6Mt+Zu5M2xuZM/ZJA
OZypgFZzRcm3ZPvXwewZtnVMtDOKdiV1O7oSyMxDski+7BHpudYaP1+HWwMf42PN
d6JErQlbsLF3rsyTCuGYPSZAz6bXVk04xFX29aoYGBW6mAJNcRp9f0ogozecbPWD
P4BnAVntwpleLvWaUcKRT2LRiQG+Proc1CXuaY1518gE/D+tIe31cErFgk9C/oG+
/kBbGD0Rnsyhgo2+krzCsLLt1lmTbj4GVNfKCP8ppFGNzRU5UWxsO3Ad++es5eXV
tSD+iDFqtpXj8JVBkcaC7mJlyoVMfSqzv9PxUIuMFh/b3zKZH2ogbVGcrJpl5g40
KTppO84kVKrLbcY6cISprds7je/aYm9xZ4q/zaMHvJkEL/r4hcBe25Bnh1OliniP
Oxg8COxMvKYJO5HMGHLKh1fi5kLiHCU/eHpL31IZQVqPjJjhWeB/xLwNwKj0rjLn
jhJ9YezBXqSk/EShhuTQ3MYLFWG5ULW14Krv/z/oYQ899bs8dYgGU4ofSCNpo6IJ
Xvj7w49DBYy3zBhq/+Kf7SkpE+fdcYp3vvrPh1n7wSO9DizL2AzIq7K+RewsVc/G
eveGoyj5SoPnPhtdlgx4wMpZrUEs8i1lMGHfBIZ3Rpmzlr1AX2/Pps/CbZSJ2ynC
4CzglmgEvKhYp5bwYtLnQCKtOZ5UDCmqja8TSKR9L1nywcxUog7p15nfsVJDIjrd
S8VqbuUi9ezIxJUWaGx0mOkozjQGql84WCnEyScHiBxjRC4vPeXxfogA7i9+xjqd
e2yLyv2EcXhKxBEr6DmpRAi6hHD7ckPxJLfxO/pLZXEuPLRPAv8QLXoiJ/wfU5b7
eDqmaeeP39er8xhzh4PSYVXoKrlVDGArfj7RLj0PvL2E7LBfZG855Ngj+2LuvSvT
hyWEXhJpq23K7fAK3tFWVO5eQ6foBiwUFYIzeXVipBh3iJPS3R94gCk63jANpi+P
VAcXm+DZYxXPEE9vfYiypaBHMhqa2mNhKACUuAvP/0x7kiBZbA66XKLSRGmf3oax
xA+oAN8rS0x259on3VBoD+nQjB44nkhwC3d2EHZ0QFtFIVhOS+PeRkXBPCYsJFB0
GxjCsO4TCIqplFqfhUCaXoKNf/LuYIxrSdNXyXRPucRA0I4jABTXUz+XeVvsbIje
8nMBozhEdWV1l+ninjldKbp9CCkVcMcbR7Gjvk4KPHpwMz1DZLTXIq+3Wpbe2QOK
M2ltcu/ZIWepY3XHvJBO7JstZy4il7YNu9lnjEcafQHfZweQiG0Go9zB9bIIAV0D
sfHrStROc9r91ZAH2PYqw89Rq+0yiwgR6P6qxMzWwm7KQsTI7iKc8FR72WzQUuHR
pTMP8CKgO6tPCmPdex5cczKs5kTuQO+W1QOhNEmRvye4bIL+6zBSlF+MGTcD1PKk
0XNIHM+NeDXoVXsiAJiQoBKiCIlMVNoNsWn8sIVUG4LXncQ8ZP96Hql496umoJxe
P3nwvh6CU04t5cFkASGCDuQ2y6J5jBeJR2THe6TUI0oTZtCrAHmEbhM7chyL65VD
C6O7biyBzj23WYZBvEnQlpsnHuYdzrQ6JoutoPChHKdv4dDR5kytlsu97OEBy1pm
3q3rauM6ShluLulMT6Z66ky/jnoa6UPOVKSBx8jZ/nHJ3uzNXeKX/blctOl5RNG5
np6WE1llOlddtvw2m2b7qg+Xbkflnn/DRJVMshOCtFcyPAUlkFO7ZfSJ8S36lge+
aS3cP6HsWL6TilK7q7zzFRaphRy/EEXxTsADpEO9juARlwua0YDLUbdVUrZ+XsnE
TV1co44xLHYnoJBS2vVX5LGJt38mT/N+E+mstP2zRGlS9+2k1isxyVG21sJqC42h
3z4Y4n0PQDOM1gqUAE0SPg/MqBapthJD/WbuOEjBVrdAMa/ZMlbwZ/d7+xXcOgyv
mP372nocm+ILsg6TZon+LXvK5BaFqehtWx3hck0Zq+HNRv/yuKxOZzd8BTpW+C9l
32G+JuMBN1m5oDkseDAltLPCnhL4izKsFXc9uSpqsYUHSn3HXI4905LxpxzKOPfX
HaqpgYrpYCj6U9J/sLqMASDzC1rjuUJIFVnKLQDUWKBqSCIjIm72PfzOOKWlSyZW
ZwQV1RCaQ/ZS5uwsY2G6seds8tBEtPD2GY7bVEgJcqNMHFoXVjxuQwZ3WPFTY9Fo
ONqhCBC19G3ZRINqb2s4DNxVPuEviknof6iEBx/9qqXjX0HdKWVZiAG6tVupMI0R
bHUp+mIW9l6WZFskSW1rYQquxgdha7wZBPRlbc943fUYt82gPJS/AcCMCxnBHfvX
mjO0VHdH0VWPAqov5JlY8+924Br8w6vPKIR8lEHSlu37bWt9JSE7AdzeIMi0J4rs
WL3tMtl8zS4cddpcZZen0VGFWR9GqCjEMlguZpknfwor/fsjRsfRsSOd5J8jThb+
rSupjMgmC7RLg3ez03pwJ6LaNik939fnVRyjy+HoQh7sOxZWXbqKqE6IUJI9hH3n
aa6mc9/Zq7COkb7nnOgkuppUbHN5BS5wLVbn/mr0cb9majk7o8r04VERDi+UjPI0
w558UBq3N1xie3RRhuOc1h9s9Cx3X5JgXzYpThjDidvrYgD91DO2ZYbUn8d5sqnj
v/n9ZxSRWVDk912pjIXpohkxcV0+waWoNkc2MdgaL2CfYri+tz145y15TrNEuFUE
/JeDHzhRZFAwk5YEeifD1sdZegtLbFb6vsgE7UsWTTcA1JRFI7bq75JNQ5uaxRsJ
qo/yQbQLayOaECBC6wgYMcvVQXjsN5dYoJFw+maYd4wvkJv10WlrXjX9H07Y015V
dx33IZJbNu6hqEcb/czzGqxNgn4jbI53cPg+L61IiB6/BNOHvdHmy9LwJz+3dL0G
TgxMHnXnVyRlIPqlIMzX5fukHQiOcFeiaRC/Xzk63CI2xzncPbIx0sGGWSrRvrNP
nKNLlAODHrmRmVSckD868zmnlbqPdV5q0uVbZwDNeVXOTetSkvQdNXiUwCwAjl3H
N9qv49zp4BXxz09iTHLEEbYfAL71vnD2gAOlxH2v4v/pJs0tMLOM1yV9kgFsjjpT
v7mt5mQzGeQIEffS0Crxbgh9Hh1uRIA4/9uAEbn32jy7arhlHppAZ15zewhCDu5g
EmJ75NupNtypRz2mA4U7K9HvtOP0TMYOiPAobwXBL3RAUpyaMOqjTuS5MZJHMWhN
f39ZqIJdD//zoxqSneoTMbbhiiHnPHCGI1xwbpRGTxX76m4GdVKHpeGSSUNHYk88
iaEHaD3zs83ayohgSBi8UHY9/jIYN8PiB6fuJtILhW2Cct3alQsy97b2xb50l1+3
aVZHedFOAcvZHwM8ne6Isv+QCTACY4xgkZ7mOkWgZnLofrOFK87i7hQfQ5naw4ZF
cB+iZi5sRs4JT8+PUUH8xLCU8TuIlINwvxrwEx27lNwEx21t+uiSaLF6+VbX8JRR
6xcnYd+8QP67Mykosa3OKLt7p7EYy+atsDWw+WvndZWbMypZdy85HM/uYhL8jNgj
UluG0st9uHkgUVGTk1StAPQp5djfcY7VvJqeHuA9pRMenGwWhxqh05SqIOUJWnld
pwTv9BeJ+iRRZWKs9326S1T0DZ2TRsOfc2o1906AKCNBIhncGtNCJNeiU+XKvwTM
/JaRGvdxwJSIshGrN8KB3inyHx/9udxVaox3rqpafJlkM7DKZnidFVd80K25r2fQ
sUbtuymb7ccCyy9ooMhiw7OVuTsxJEISqm5bNQqd1fczNVbMY0c84a+CQSkwm7od
kQZkuGRbv6lsj593B55OR/Gn8xQDYDnUT/WckvXjW4QgQF92+zqfCSqjwJlL8AiS
NkizRSHjYAGGrya2kxTFon9oXSrLOUtz0fcW0SQFDAfnU6315DrhCCcCNN9fI0gW
S864csGr9FUi5g2Mh4j0lRSIbVbcrIlOxECoHqfW5Vicj5iSOBuxWEfq4TvGWV5W
4jVS59Dvif5FjfA08qwjiFSSHHcSWLN7Yfc5bgXQagFuD1rwMtXBrRtY/Somh4rU
bBlnAB6ZGj/ikHKXZsu2PZSRSryjrLcLlnkQeCUcPeKIVuEpzmXn+b+pi0kdj5Xb
mM0xcNkPVBBTtE8WdQg4vOD0H4K9yIILe750ziAyEIbgEouMhoZZLJPPGPei5DQH
ixj7X1ix066dfP7eGolIsWdxpmRk2YfDVYCwu6K3bYYQKP9mFzaskKUn3ppOEc0F
r399XrfsGpd8Nds6DAbWKLHjgfl3/11OlDCTo9aDNTYrceexOxPQ76gVJ/TMlAS3
i7ogMKflS+ObTeGAnZb+MqQWtcejzNRKLjFk3NIOLsZfP6axgJesPSfI601hTfcd
/ZnhH0INbgkWT5atRXtv/uYaFbgQk60voH3osqshgptPwvPymwX0e5Y0TIUaV2mr
t+gB4RmQo4upjtvd6r2xJW9OIqTdb4vUFIYcKoLALGOokFfQOXSB0KUfuMqjGr6j
8arqZlqw+Lp4aIRmn4EQjFX/UWvElrgFWfHEmRgfjzslZPnm6zMTCXP3GGMfRgx6
Mwyf25KgmUTxJIUoV1Mnb36pv0TNz3uzAwTVmNz2YgU2djKWvRnEmT2hCKBjiCOX
2d6Ly56cH+uMJeJ+lp74l3wfAah04YcAAAppKjoqzarbAwDjnnOjqD4n0BY8cAYR
MTXguggbMo3sNCo6fHyhScN0vFsUNqNvT6Fs77Zi9CCTkMvqREKk9lRIPWWgzhAz
YNRyzzDShSwrf3FQ/5tFzUmPa6fRXwQPYneviBZ8anotdB5HqIcj2uA9qrUbkdAG
DfeF9T+btGiq3tbV+NCB/pM7Vd0Eyun6Ua2zrJ1JOS0jK43W+zF4lj0CSYeioKkS
7LSAwPv+1fVHT3KifzUPsegbO2UoMBqKpFFtSkR+4lk3QvmfU5txOl3dOVfFmG8/
aTDvDrgdVKmh6Axkz9SuyL0FWTvtT9CfWGTviU7i+8XSABjzxy6fuN6CcKSsE0p6
sr8kN5DLxKZwGjdBFW6Wc8rln2r8IA+ChgSYU7ta+WACg5q46k03xPFAgdO6ZrSS
5tfqlgFwxeY6Md0TABOR02ZtzhfWWfVKl02U/jD4KksmeZKfliq8Hn44Qf8iaI4V
yVNU6Z7ISSeXi0OXU4zqV2YeGs5LduzsfBAc3E1l1tXjQcDVnZrtNOuzTtoUXkri
8mBIcaXDD/BQDpm8HteCTPiknPAkegV/yBfiXt4tEJ66aoJDyoRn+zYZM+CKc6o/
VmpF62b/ul1BtpF6oZuGRXCc7z8JcuEP2fDLj+m8u9WwwqHD1rjyeQ4TJhCcNKnf
ZsPamhOGKyQw39Fg0cHlmrKWzbNO9VYgJeBzBimvZS+exF/8PsffYZ6gICATBG7/
7hW7Lw2MFLEC5Q5f1hOuxzFPfhMdQ8lQ3vh8575dS0mU+Xlq12NA9XDpjw1mTk1v
g6wq0iWemOSoM9czskYKJe7TVY0iaOut9hRF3luUQWg=
`protect end_protected