`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 9584 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/9huKRhRMtvnNqb3Z+UU7TahEoHV+T8U3P3ufru7l1O
3DlgtZzb9QxCbOjthp9+wDkjygH0eUfDrEl1ovhZG62fCGt+wVXB3C2rSVlS0/ih
0+t8njYVkoYZZBEzgq8iXtFDCk+RQFI0/U5TApCcO1BieBBrbtacNRxCAQYf904g
v1gv+tYK5az+mNMbTAuFHs526co+tkTuhPXORcavU5x/A0L6RfT8i74pT1TSXSEw
bPSXW03fqH7+JIC2YWT94beYvgzGB+XbZ2XSy12vCiBNDGZUUQMMe1n/mISTAoPs
sTcM8/nMPtgITAFCZ6X1J8N9GAvi3R9ZxEn1YJrdAXK1188iGQPMkwMS34VrXBud
5NYKuzXDIPwRk/L8HM2Z5amO3jbLx2FW7tcl+S8HTcXsW+6pEaDda+1tg1iS1uCm
JAyGp6RBg2mUOdgzdAqq6yf8gmted823rVg+VkCSuK9EfMAx0DDgTHFN+9r2sHn1
fVl795SgoagOQMfDhWHPFvCv1NfBA4X4yepDV9Fl6wLnvrBg7tYWosyl3OeNCZxZ
1FXEFNvfg2cfZotGRcsgFqg5PGrC4KKcaJW442RrFxWk/J82zlLz5fYZ73iVjoKg
OnfONkjjpdxfpw73z2bW68bYvbrpHFdZE61GV92VuGkBgjcNkPM+2M+THV+Uj9pO
dz9IQR9iIzJfhxdEx0Rp3s0ySw+D0JYxgEO3APhRQ8rKwXwsrPdeTtl2Pe+qRw60
9+1rlE70LdRn8eOX6kXyf068Ti7Kw3W3L5Z5IRUhXknpO30l1MUhQXnT2aiwEY8N
FuM7FGRQMpoetdi/aHg/iq9ZQhoA3bO76mc7lRIOhv1sVYATYENoJwLFYgir7Hws
C1tgUZ4Es2g1omanrtLJCR3mo2OuVVVg6NBF/8aX6UArh2mTn55NDLcAWzUMTrM4
lcTjcIXOUu10tT9E6aouaX61GE0mu9OqCJjustzBql/w5yUcH1arS3Vm4oxrgi6s
kfUMW9PAIhJJIM8iD6JxeiuwXMIcDJKlDTgWWA2h6LHfxgduDlEvCltD/zhz1A+r
AYnFD1+ijQ5+TnQjd3at0JcAseGICjWRNo/rFm9EJrHmUDLQWPu5q8T3P+uIQMlV
dIyPWYHTKurQ4RoVH/QCjiXuqwSCTIU1rONZbtGonYRftqms6LPEWqL/AstQrYWc
k3OXF3xi7AhU/rRu0ZhE6mXUGy/t1Q27mc+/wBbhy34OEOdPZyrwJAonvZIFNMsT
2P/+mRa2cAZxXlYsSEx7ELF7lrjt/Lo4mrAg2IPry1DtGD+2TudHQvC4ULYF1lmI
tqHONy01VxaVjghEQ97/HIJcRt2yizvAdHof5fIpe6qT3NOZIBif+JwvUtOxNXAf
lv0W9DPnf1o/2LzrOOoxlqzRODXBXgt8iJ+ZsHblGTgIKNAW4uOp/MAcZs1Cv4RO
CmZwj0IeoznqcOFYPXL6J2awncxup8a2ZnZhYOuACuX60RBZyIvFPwUWMCTn1SVW
Yc4t9sA5VAX2HE1WOi0OT1FXO2/0n3oomeP9JxmDMIKTyIdY/EBlW3mhNcAYXTLr
IpLTUdgAMgNJ9DkT2YcYApDuCsA9fXHuY2PmopW9NhWb8cLpmSn9VNlYwGYDXPsW
XOrVDsyrLiqK4Bj+1xaKm64ZJsW2Xm4D2F5DsYCASq1AwDYMqx+++5cBLpoMclH0
PygPAfxioe/Ty8pXSi/n0zJ/bFJ5aHsIOpw3Y+uAi3aqiMJ53W4HJs+ma6MVxk15
Yb0fRq3PD8twY66W8oGHhr/32Nu2YgzqRzlSN21job34xYGN7kSiDrXKW2JXnT3k
4ccoop5OKyEd7uoyvHZm077aPKFW+uBJVNCTMXc9U/epNut0ZH/TqHIvBqUq9FG3
jo0EVhqOXQZEbMiL2r6XDbVBPAwlybrYkZVlJVrHgtKLF7bPpKQWoV1un52+z0X/
WuDQVIhBO0gQxdnnfwFgzVX6LePTXODz41auv7vHbJGa6tc2EJ1KS5vj+aajAMRM
dPY13UliS6yztk7DE/iZIe/n81r/3DfkfgIDzyMsJV+edcTJmmLy4/injDpg76Ao
Uij97fNU+ebCwT5iWnDlHxOtuOhYDbt95PEpqBJCOxj758L4RAiHiWw8xCuJTZfJ
jiPmYGmyVJSgnwzfCN5SIXzd0nmEgNsnuI162IMh1gaN6TGABQlREJzur5OcUoSV
q7wI1Aj+jWJvaZ/gAKrbPWlRIn6FeUufa3dpkuTdUIoumYJ1U1+UeIkSK1E8JMGP
a5wgp/QEfGPAF/oMeVDcoXVvCSvoszdXL50ibA+lJnzUsBayibQYCnmHt7LPDw6p
I2c07zIS4vnBRkF68uAXPCanmNglPPqtjlw8YiiVbOfYtervcR2VMniZvEWEHJ2+
XA4vAIiYzYyrfQGlwvL4G0jpauuoZzW5QGHuYTZgeawtTEluyre6xPnGt4NqDHDj
q7n/tl+yllpCgW+/YToxkcgn7KBdwhwcVtMD1D5/f7sQrtb7ypFC2QdoEQFnGIvB
n8p4IbDJ7VouhLFE2NktRXyF6NDuq4KkYvBoCLH2GVduL99t/ZVWrRXf9tw10/am
yndMq2exw8Ep05ypO6xeJGfExVpee7uTjdwlbtnwK12EdpXFDFbTsjkWoM7DCG6l
V7D7CXt1/kQnZe5Pn0JZuJmKeNgN5OHbNWDcYvjBOOwcYhhoM/LSCeSt9Ny6ZCGh
i0JLFfaM0u+hJvwi1TaHW2/9rZd3xxtJZqtVSwZgXdDXXgIOd/1mMyUJdgWQqzIG
hSP3EuGMGJpKQJPHo/X2S4reoP8AZGpTuSnm/urfSorkJzm6ZLz0wIJLRLd3GR8Y
2qz1iKzBJtDLeDnLR1dqPThiqYBKuW5/WQIYybEjPgmjq/XQkvS+8rLsy5Agrb3a
kozrnLeRm+ITW5gJhU3SiZF8bC5hRgnndtyvD+3qVvC7qSOjTNc2gA4dEeRritPs
7V16Si5AZBRhZEBo7d56HZlJd31jbUUYCJfgSgZa6H9hklRU06SKjr9ovvcs2WsP
QvfzDZRKW+ML1OILtF+jOQ8kW6rGPxTi3nACt2RjDy3x5+MJUWAXtavxeujNgcgX
u+B2zSY5btL/f1jlUZr5pe6eRQG6FvnfqNlU0Wh0oAHvfaIZdIdNQQgkIX5g5jmR
Ue8e1aB7xQ90QWY+rYQSQF/Qy1ARjo8VJT0v5iacApi+YaKV7I9M8L296Goiqk5l
sPpUb46i96VIExhPIeSKSDdxpPR42pa+EqbJA7O0GUEpukOeYhMSif2MupEya5WM
GIj7G5VHtbLS9OGPTfK7tkYAIdXSaaUO3rHrrFVskSZKf8nfSDCrZAE80LRI4658
hOkW44Wkfdly6jihOKTCnXnmM8GNmVGcPZoP+VPtCiimLCZcT+dIDg8APZW0ULCM
z+zriNqmnbSAU0E/tRpm6dlZ6++shBF6YpWlk/xmv2zlmHax3U0JfN/77GSFdlXM
vgKGrpTO1RjmlT9laxtyXAYk6fbZZ2Lre5VK/zXudWAwiLvkQ0ld6udgioyZh2Mu
x/q02bImDpoXtp+yxodbTcFOCcfwi+I1K2N7aHW5NRGmhkwjWUF4QA55M/jxyeTo
1C8akq65d+o82ITE5li2s1X7KmFXCgJGesPtYlOhSMdscDoPfgTl9zwoO8AX00vD
TMI3NF2C+fushx0WxvCjXVscQKWntJb3qmqjrGhRYIqsxAViGWO+1UZkDZ3L1Boi
tyD2HVlWT6jjs+V3l/Xg8mvbUs9HiXmXxio+EGzG/vy3VvoPEkmQwXzhkwKNb9vJ
xO8g7QZDjxcfiosyHqMDrZNxN0Jcj31kue6lHRH+e4HdBMHQCK9lWU412CHlIfEv
IZkOwbEDRE5yRghXc4ubFPy16kJRHxIKM4ef7lYQ/mSuHxq9mc0PDlkWSGzlWVHT
Fyd7nbth75aym0tbJcIfXgtc2RogjDsPSEL4QTEQ9t+MCa/rXiCu17ReEBdB/KUu
6lptiiA7LFJeyqUSJ5d4CIaiGoKC76yWPV9WOYxS4NeuvduWiQ7pC8h4iu3UT/hx
xe69Wi8F30Lszre06i2i8xmFSEfE+9Ei2/IHOiMUD5OJOpwgSzKUZ3VwHYCEnv1l
0BKtXZyAaExbmlZPpA6XNsWHvp0XaViPi1720EYUzZRlyZlsF1uQih+cnEkenjti
Ip6jDObED7Ufdzr5OrdRr2GnrH6c4p/iK4OH+BglNQ9ap3lDrBI/f2YlP69kUkLj
r0jCvhRJq2cYQz+usV6CT3rFKsHp5ikmBxBkEsuw9zi31QgzbxdHJestvaPvLxg9
IRH+E5w6Ytjx87gpok90kUoqDMqlvjdFS2WGajvgrmrH4TR7lZ4gstadDiCMMKgx
ORuflJvQtc3rtI2Vgt+3a4IS6j7Xq7JoXhprAdDmWsPeYBOwGQ7e+DM4geru9044
ydw+WxRaGvriVeFrghR7CVNGIUkbDvCQS3lMZxfTKmCeX+wSs4sOdV3l6h2u3pWy
RV4w9W5a6+AvXDgqYDdFJd80eNzfWlH6Z13KpV2yQ7rHwQIM7rGkCcCWRAxDwMw5
IzObyKYObXTI7vhlvvMlazzrd/DkXfFLcy4TknglNO3rWuyhzpPWfIoHa4VC0Yya
2k15apWYxFbWhzQeUZ2nwTTkqQh4qaWsiJeAcfSw9qoNxvtNyJMJ8jLOmU3clGum
rAg4dDe+xYqRmBu16WT+lvQNBunRWCVgX44ec1OObxEu7ZVxfQY3Nprlj4IW2puf
Zod3GxwIXn7ueIflhACJq5xRgLmUhkXFRz3Oite91X3QGhHuViCfvZzHzbQDoVhc
PmH5u7/rKcCUcZXB3cTBfn9kRjEveN7xmO1BvqqIUzqwFDavrEhu8sxzFWxRr8Gz
rS3oT0qCtl7ly8+oENw4vjCekRYA6vySzvI/tCjipKMWJjs/t/73IowuNV32HbTL
eTlWtOWfqlk1I7M8WIwgYMp2MCEsGioath5KpJ9ZP32jZFNSkbj9d+cRBDi006IZ
HDryOdIN5YAZlAitddKxm/+4ctQf0pqy5CgcU8vmZfK7ao84TCewuR2w8y59Btqb
D3w5mZTLQNLkPA4L8VHWeG+s0XUiBfEuJQtOb1rgs+KZzemYiG29YIuWgucos1n6
qdgV8IduniBZSM1HidQl+Ea9JR0w6YGGy03a40XTq6UdF3Zc4GNxRn7QHj5ruo3s
/mCChgdX1zG8aUvDx/Hztyx2Jm3Y5tKnft3gzikEurSJ1y+vUEHaFT5UcwiZQ/W3
15vyo3pZthcE3zSdNE5tjJS9MQtt2n1LwcAjpqyjxeVGODJJZADyYOUN69Kc7R1a
3RTKFdvTDdadsZ8/oksi78xfLDsq71+HRla9X17dOfuqSqbhrru4Uc68NAkKhmUk
plvPXuR994ZzgoSc1fsYLU2AkSAD4jDsHlhmUC8gISj50uGzkwTb3uNb70y+rSKj
9hg8bcB8KWe9TwE0wrgGoiizHIm7ESVoiCSf7T+1LemMK8RL6mKumo98J3X79cSs
da1EF5KrtloCRYsGGt/krPCkwTolnVXxWCVZFgntgOYfIyDOrdsQUq9WG5SmMOfZ
6bKrRJ3X7idN7Zh5DOTq0fV9/HVc1p0AfhySFLO8YVP6uJQ7k/k8Pk9rnbh74kWA
L7TFXHONWWRuxxwZMBIPclUWBZJGr8wp/MJX1CPFNEWc3zYyiBSa/SVAe19HIRtT
WeIiNibe8fAyssMvirnbZnffdXSQ98/jJfTJcOmiwd3CDdrBuQEBNWuU4qh8q0WR
LcL+KOlOm9AcxprDHoMha48W8QkXLFlh405C6LnWmc+Cw8h1JKfQMMf8n3/0Es9K
kdX08gYZFYbfekw0QW316bqkYZGZTotcZ5NnSUPczBAAIXcvTbPwumeiBuHMiTGE
KSkKzQsGZQtLfKe5taihCElo4JpyidPda3pyZd+HMy6Bii85J8PJwa7V5drFjU1G
2SCkN1eOt83eYJpunK9m1lWbO7Qc11LWFQ2u/6GzYw5QMJiPxS1F7MpaPu2XpIk9
ds1cf6W/LUnkm94rsz/d5pE+NY1qGJFsxSMKWOPsd020igmu4buqhFZukGZ+CPBm
K02KSUCvK6qorFlG9wI+87t+3VIBL/hbPLojM9ftG4YMXNPNBT9fp8S5B4Q8eOQ6
xRenbh30flpusUQ+/VsSuPB8//RiT8RmFQcfS4ofDMixxT9gfWQSPXk2dhfh/IID
XBahBZAvvdA4SLzxWUmUoeJ4wEEb9et/OXCVxjqVpnUI2gmIScmXnCwVcoq4vlZV
9A1pywTruoHfNxKP9voloHMKYeETigYEQw9CogdJDjHNy6c/m6TyABwziKMFAjEP
sA3+SFEFFwx0HIIU3Zi+QPNbCpIAgxctvWhWeyELNj/BooFUE1N0SmR4YJNWg9fe
F3QWM8Wi/o98vICTBo9xGP+A5bo9jWWPANKVSHd69SICRggfR9mvdB0suSR1uCnL
Ch4/a9OiJ/WfHn+VnTyI3zPEfuC5TNGAF1CIUhZN+axxWBG6itSotKjZ/Mi5aQCM
3QKFe6xkvC2nl5fxfDQGBUl9EwoaUdrCieAcIXWmt0BQF3tAJ32hfKGsrZWfGg+4
ksYFeyoC74ycPLv78sd4uMLOsUSePBBPIfWv9df47cCQJDSdg7uYq9/SFuEhi/VR
BjUq6Bxby1ZvoH5gMTeA6+B7N2cnAkNdxdXuMbWS53toUbDreYrJ8hScOLy/xUGd
M5Y7kh1jkZrNs5MS+eoWTNxXXbK5A+4WYigfPaek18Qnp56+R6IkAKuiezmsqLWM
YhJVAS0nI4Q8upiguyV/cyhy+i8wd2ystrEhhVoEmsV+Wgn3+3QUNKTl0fVJMO+N
jpuD9Gbl2grNPv3l2xYCnHfrCWtWRIV4/0hMY0hPZHIcQZhWtNHmQ2qGgvHLku5b
dB0P12rAAHD+Tn4SsJ3Yd1UC2XjqnLZCxEUtIf2AKhl6rfLUSdeObQktA4rVIQMp
BSvsKA9eBzOX+jIV8JDEZdnqKrA+6OrGHjReB7LbfaSfh2HcQJV/P1KVKeYlUfW2
wkt5CJx9phLjDYSNhb3+F5q9bs7qzKcSFi3dkslxFtDW/0aArwz+3eoOAuBtXDWQ
B100JwsgkrpKfPHGX5f0zgp5RFvE9SO3ya6DhCYcoTw/UMhq1j88KXKDRwr4+0OJ
ylkOmegJw8GOPKCZMQqkBnm6I0FUyRyXVDmTTQVwitOrxLEhq+ztu2G91Ye3MJcj
MA9X6fFB9WJzvNENk6XKqsKXbncsQeUcvfONappnnmho2xsD+0ORWAWNpD43wJTL
5AkB+v9eX0udGoLSABIB114nnBeFmhg/kDILCiGtk8c985q6E3NaKazFoS5eW3fC
G1Y88wtywDtl642egyPXTdv+rjNGWq27TIayPThFBCjMjWYJpRbfwBtwuAY25y6B
oIQhaTn17GgqeCaTGvZP8sZrp6xpEBbCzzvJJIIzi5tkw9KHHJq73FgG76omnR5b
mbeNNjDXflqWIESxsE2R8XztHOjM2Z0t2JcZPYF7vbX4wpxtxT8Ee6AeJlnp3s6a
YBo41e1MgSbhM9bD7yepe1W87ftkCBu125Ue+fkI2LtD8xtivW8Vx0EJXDb/TD7r
fdVeIobolubhb9BdTPfOG8aBe+AYMdja4FdInmfXRNYTDjy6IyMM7XEeXlcfUabt
3WMoEY3SL6K6CtJiOGvEEva5XzSVzRdOl/y4N914hic/6cGOqcEz+MZH7QbSkb6i
tj7SGBXco5uhVKFZv5BcOe9izsVQr46qcsh9d7NYAveY71RWpV2B1bMZm9oSQjvQ
95k512X42Mg8/y8QlmwQuyga/Cy5dUGJjiHYoRPgb5rrjbpF8pCYKIiPYHW8+4FS
kWP3+E8SlXRPv3b3Jy976nkAkSPdKb2+Tj9vXGtT5vlse5YFIhEQ06E9SzJMemyU
i4olnztoC8FvQCaHIk3EqNQoHy82hQN6figXL3F5mfFjYI0Y+8HyQFhe6CbhbjOu
/P90wjNgA2+njoHLbGeAYorBzfCoKTjz31rojCmUYTGryAB2iey1ZrvdHtrCesqL
4mfXq0dUfWvQ/1wlPFQKUW3jAjbMivh9o1gPMObi3uwips4++N2RLaW3pB0Axxk6
7tFryB5qbdSzQo1dYUK6qZNv+/wT/lJ7eolrHPYlWKGBREzPuupJLnm8J4fA5fU2
h8O+x7wZ9hwizpTQ4E4UyrCcXXLLuvqk3AwCYIt4xaca/TIsv21CM5SQvk4soeT9
7NdNvoqSRpSHby1FGwrUh4sCBoCPfU9tEOcneHXPF9ln+Jg6NxB+WDO2yhSmd/KS
aiZTNsZcXBBHpcS5zmguyNJWnPfhS8H5BAO8CSL9fyiWm9HeCWqj90uObSCMkUHW
L5hOf/vDID+YptnrxJJrJZU25rEGMT7mDXpdzP8/OjVSH1XtMDl7iw/hUiqBhM+B
iWrjXt0Kpv7E/ulfoW2+rONTigvxPLZI7rPSIJBaCRagEIxe6+wxDbIHr3lZS0f+
RI5r4OPOUl7xzs7IXMiIfIQLd9Z78XM3ZPt+MYL0ayr7bKiKNPry1GIEa7p6b/GE
i+OQfPvNPUlUbbm48IhU+iYWacRwO8dlxOY/GeNAtWsZC4AKDRubR6ud5T48cw30
b5YVqelq/6aL2nj+HSVS/36Pd38JhubF3wuPyI6s9fBQZOEKavSathVy3bTLhTW2
gQmC45NVOri31RVrEMTO0aaSSkNxDDl7ps4wkctc8q2psrZ08XVE6E20sS6+r1wv
ow3vBUji85yk+doK/BcRYAp8Syx2tAT363+RZX+Fb255WxB2DZ5Xqgbo9GXdRzH0
rHrXqEU7zUGBLXupusctz66wV+sKLVP4p9SuBsbAxgElFryqSMBCzo3q3uccCD1n
s8xuWushbFXafiNGKIN0Oj1d3eg++mr/MSKrVgI8EZ+8Lqblf3sA2P+LgFBG01HR
3SCwXfD8eUEkF3JBzE7rwP86n4gDcyNfJkmy0OBYmfcE73CZGd30FzObSKJy4GXJ
NPkrKV++pypLrB5AD9O4JmyqhUhCBv6wQyhqAhWc+Y3OzComqzvhXNKqGZholjIT
hs4hWWMLBkzt7CEDarW5muFjppGX90+K7DlMzTtEVp0/dknRUb3OpHSLug7mf42L
Dq3RUBZWPngKby1AzO7Jc0izlIIdIwnU5N56oSd43tGQUy6UjFNoq1qOou5hHuQ8
Tvj20waLyBSGxpOkJBZXxqR0w0OWdykJJNusCtJyjDZ9A2qIe4UwKes+a2c659YR
1a+XSedOTfHsOl/IVM0dQ8BqvKDROv/Ylty9QEs9uxonhy1J1GOPU3lqApIHH1VF
G+WKa+s6poHN4ov0aVUrXFX7ak1AQ0YH5g6ISqfQX37nIO/XauRHiP9Q+2HV4OiR
khIsx6+NbHGavHVIBuiIuJLSAfRC+i3H3QsZA0y+uoLPc6G96ETajPOlxdWLbyGt
cN9MyXerhKXHNAfV2mJAKJbB+z01I3oNmHLTwt+R/Feh2+m7xOtjSKKjjPmXT4jS
O7XUqW24X5F5CXqttz5Q0bDaij6cF4pPxbEBH72LQCVgqLiHAIJf2QdJ5fJRb45C
YjU0UDlvJhC5eKsJQv1J1fEI68CM/spB7TFUcRO+QzMF6OfZt2CQZB7dkGnzEuwm
GME60BMj0UgyEIQUzwmWKyQJMvcsJZxPCd6DjY0gDkAqPCgxkr1bFnJTmekM4rte
rQLNn7KRAgBkmYVdtJxkyEBKL8siVke62+6AUfoVbDiGqc5jWfsWY+amuuPfKpcG
bLQ1hr4UuIgdXMs8+zlG170ILy5jhUMR/YtMlvjfE7226b54dxi27YuSSHzFpbj0
pndbTKSFnJ2VBr4B6BB6KQKndtbc/wwXu88HjY1vRBhiKfLcfyCVScfGPz39deYU
4luUJ61Z9M+GspAsR+TEgjd5/zWvqmQY0lK4/np5HR92J7fvvutNhzao0yha4t7r
CVBTn6AEpywjmOb4+/5ZEN8g2YQOotLboce1qbJHPL+qRD0hYaIH2TSkgto+ZcWU
jATqrbqgnl+PmLlMPsOzHMmxsggPTJ4RNxcO6f/tGmC30NL98BSNtzZqtAMTvXEa
orL8J2HYGdIg+OqNQy5wXdcRJBMeNNETX3WTEb7tFxrvt3KQQq7snKyZB8u08Xz2
aFneLNo76s+PyonuNRgVO7qv7AbO9ufdTb5JhvlEmBtmXSCtsnIVCPDyThSYU2/A
jzhJOf+APDsbNuUI6DfnRaUaQ13YLAxmFQ4CvnkhUZGRZESiNnczktxTW/blEy92
HkXDIkVkpcnqnpUKhCFATN5qyOIAI5dXKdTyTBXIyVvIRlLHsyuzCSm6LwjsCZsz
WqF4Zr4QF+Ht4eYvC9Xa17sqWk0CObZeMtk0QjwlJpe9WNrGEb4xotIrPRDYQ0t2
Lv2SsirUHD8H0RqLZUlxOetlJ8leFJNBuxiL+bmgFCyXJKY1RsP0J3FMG85m84ZB
5ZTSEEJVrs23j8pWesqftyqlmV2pSzieA7Lfw3RmYs20iNedJXs1sfHdTtvih2xt
U69/CeWSShoqAJ+Wzc9f7RTwoFEzUHtF8SEwQ0zz+dyHChOCQxGeG6361BYAofGg
CM9m1oCWFDB8M1/r89FxXmt10f2JvOJpYcWAHDc31R0SPXt2aNcVvnH6K6QSf3KA
+ZXkmp5Yxet0XQ5baTGFtFY4BXdCKO37mVHTyMDOOVinuOkXqCnuS6bGrITktNFX
fmnLZSmxceBsytJBID/BNOLcyxBzyWtLcsZWYhfF18nF+Bg9Fle1A4G+QhpXMEtO
FH4X2H1z+Kd48Hh/6fHdXupp/ikLNAK323fDdixcwe3hvxjHcWkXMEq5+wdvxhSl
6BMPfU5axN7/dK7HSYp8MTYitqQ0qXD6HPjeHFeEs0QTWs7RkMYsL1BbI9WgrCAn
MmYsGQjaBelHbzOSXr/YR8zL/zbmQqbBs2K6bDVGTeClUsgn4bXasa5rXbiuxLtL
ebH3Kmw8c60maiykx3fhhCtgjrwKjs2oTkc4D9FFHSwVwTKnkD98IgWVgjCl6ids
yarzQ1BVOjkB1m7rodt84RggWWqa1V+8ZDSjIEKp46lomRK5iNjy49eca7xhCV7D
N7Um0j3DjciaHGrELmbZ+B+PUATNpds6Yx2Bw4FKGMTpO5DE5hhu7fHwIb2tk1ds
u17GBkGxyHmaORHzuaajoBvgCaukXPWLy87AHqK1dX9gWNlgBpwBls50iuUP5tc0
Qn4T+1OZy6YpRHanqLaUnzSGPWO3Gd45AxTnJh9cLDTyBjjgmhFNhcoIbQO7yvPV
LeKfARX4N64hdd8WmZ1zWTmVcz4rQkTOI7j6CIy//iXLXkVA9A1Eq+U00RyjqVBt
F9tYc/3d88piNhbu8LcwLO27XC6k5nbdabX0Koypn6nuIIKGuHmiRlVB7g1NVnA1
YRakDltQ3rNt3uJIxTwxABCQWPHN+yK0MQDeAOeGz1m3VpOqtNx+clXKSkR2h9Ld
mULZDQRr0cS6LKcnS7tSjrmeGzOXETEoq0Izh6wet3l4UROkNWHJiBb21mw6jQ48
YYzsVwIK6i6wwG+hy7J+52jVHQvbpuBo5jP/osXOeYDY4wBjHeTGEgJKASFEJdlP
Be98CTpadCqcV3TiZdUIeTLRRIaD8MsqViZZklU214z2StUeEXARgVidqLmLfdJJ
vf0hTLEKf3ug8Cgn/Rs8ctGmYkKRAqCBBtqcyPOTPICVLvGmP6F6TmNAQB2ROKFM
IV9bJIOVKNHD+GXTR9NlYfC5SR0jTjEy8zlIYGxYNw8FETNKUVOnjKpCn2xUUuoz
uqXahPhnaHwRKs4KVZNsl+D4cEIG5ADvA9ajy8Wn6LFq30uI4IPiZ9x4HlYwKfKJ
p+kRzbrfkIhqgnILx7K64MSnU4qY9W/3PVQgtL51CCFaaGTCbSNFfvYlvuZ3cp3X
TcNaLwBACljL3QubZe22Fg9jXU0gE+pXPP7WgRLwRHjr4Oj/AUspd7eEI8py3lCo
K/ymh/fe7eaD3lH8RQlBIZ8BXTQFVIkg+WKT1YuethjngauNH3guBaaLnn0zqxdo
w4ie9oAMFp0pv//egcyyyf6LB1DdoWADDgcoHMk4xoVUfKIRYkYuTO3XpAyA3Wln
kGE3wNHlOid8r3cZ0xNHQT46NEnVVE0bDpGwLnnYwG/EEN/XAUPbAujxwSnEZvkC
MFUBXq0PfpBh/nIbdCWFCDjhUYAXFSuhDeGpHAT3STsMYabwIEEOwg3yAHOuOmB1
1uI+TVLcb3neeqqy/ZAmlVgeS4PII0ODjMHQzR78miKvpTRFmSbobBIWwCX2vjcy
FLLcizeoiWmnVMDFkyoYohkA11Hc4ef5YtifeUNNdT4PVHabN/vnarFii02JhK+X
INlUTd6kAwKkbOv1HGM5p+xhFDhKV6NdCAyaaZ6ADMoU9N7iHEt+uri7aObd97xg
JdCozD+jobHcLSuaiw6MfimrKOxjT52Y/Y3JY9Z9zskJ8cvFbii3cBqDXpCJmdrx
NRY/3vrcr7rdH2BSnitPBuHeXHN6nDzwnPhg4J2UNaukhptAfzoAdzzlBAsz85/R
cQI0Z8InDCLo1Jrf6NdFUHuPeauCYyuzeebur757HRrSU/HFjdOkUwycnyUkRk/X
Lhty7sHbkmmnCbtdSWh2kC4XD9LXZRuIobd4e6FtVSg=
`protect end_protected