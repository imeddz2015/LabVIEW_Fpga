`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 111152 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/9huKRhRMtvnNqb3Z+UU7TahEoHV+T8U3P3ufru7l1O
3DlgtZzb9QxCbOjthp9+wDkjygH0eUfDrEl1ovhZG62UfxSNOC/TPvAWh4pm5AyA
oZY45JQgYtONChd4CkB2g0zRokR4R+2OsDE4rBNTrTGWteTpnQUGHrAUSjog1Uat
ljrdSf5ei8Y2YmL5NNZlTrd8/7pMgrJWqtDmNgrisDLz4/1I8hWVlVOspA1shhDY
UhYfuNVSf8/8r8c/BQ7AzzWUDYJ4H8rzB+NMCQHlLA/DGYYb/fU8QPqM9RceR/t+
+2EXYApb9yA6dMcVR4AmOeBqXr+2fOqPnZU7ZKXXqsaf08yi6859/KLORGJNMLRv
sCI17/kTAkqu/Mq01bL+epv7COKBexye/lJiR6c43dktY/2c2lyYlP8CS99SpGWd
dDUeU9aLZE963As8EZ+w7mmoRBitP+2GIvWEiPxL9H7VCU1tr5uDnjR9TNAsXta8
eEtoe6jF/tsd75THpdZTU30wsiXnl1eaxR9+4XafNkS9nCvSsJOS2LMMqAqz/5Ar
eABMEYlxRJE41rq8x0H4DCGHgxE25hVrPO6/z1l2IcSBIv9CZh9zUVQ/JWcqWCES
375feNTqQRUUkp4WTjW+b2gCG1hdkRohg1aMOm/1daFuTiYT3CJdMjtakJ9LpTVm
QxdD9eVFgDJnH3Y1a7IPVQJoMU02DsLocdCvrkSOBcqrrpiTYcNJLKHNH/wU15Oz
cnKPiFEm5df7Fq8NrjCL4OT1qZZg+UtRd7mSFxVRxgvAjg+qQQgQKBpneyGXNhNC
Qb8Y86q97lwzinjvKayH2Asu4WII7Nby/Vn1/H4hHrYnFbt/cx9u/sivnqh4XUgi
47L0rV/AMC5j3WTZ6pVg2Nt8XSRGqa85iinayf1sLjSY2IINwO5fVQ25qmlz51VH
1u4bDcsL/clcS1Z+68nQq7JH/wUkrq3uaTMxOHhebzGWB2Zvjf8BNFxr3OOTPSeb
lyJWLTQjrFEyQBm7OYaKo3OfPDv0Sy671b7JS3zrhafguSEYeiG9byhB4GcFgkl7
Ka5U1iShNx9eRpRy8lOtr93ysgU0euwgyvmoD4ACsJzt0oO3O4E1Yq8AtrqbriQd
z9Vp2Lozas2M2THGq/+mG+shRUa5KN2ZvxLsYyLN0+OALiML5CsoH26/RdZSbttO
wMIrDMnB2FfDPffEWHJt9ONcaxyRTAm/Qj813s2M8FZwvnvF3O0i1oh481WNK/jn
1Gf5EfS3kSofyCWV3AbuI1Q1+MDr0mFcF/zoF3FdmGO71k/+oYLSVZIFxJDbUr6y
XBU/ihP1/4o9OEAhiEYAKGgoPy9JtLVjDzj4x1GJ3q7CmKKgmGniCJAspW1BY9/v
AXhK5UHUdZIFpzpH1CcpNFrDe5oT7leYn0htnokVHMRuKWs0gi4O62doXPPVGaFT
tm0hdWTGRRdJcuKJrsVVbBzluxZQ/vYRFQlNMaKQ0/uOstuFVeTkt8SZN2VciL1F
g/HeEfgRI+b2XxiM2KjajNjbphYfKNLOX3WZGR9JGoyQxGi9YcRHc6Ufy8Rj1+Ee
hkLQr00Y1Mawhi4W1+1umjZ7MY1rXWfAlE/Wb0Sii9NWMl6uKTuiozgMH9aTreC6
ZnOpxcY3kK6Di8W4LnOrPStWfGgASAUaV+0wl8MeKEWWH6919D8UeCmqYNOk4m9J
DFmyDWtaorN4pW7wTksebOeiG+xgelRpipsNErGg302jVmNB7MS/vNn+3jY268VL
a5dp/RjH1Y8P74RrdW6FVgXZfHKC23bglFT8noi/wJdIcxaqYN9mQNGfS0ufJugI
TB5FnKLVJZK+1viSRak8bF17Fj0H3FnofrLxXAvNGJTzTCoO40UvNxdaWBpACZMN
nqhVVu0hGVSyyieyQ474sPv0PWgkBkgg3SESveel46ddZe7vrFBouogb4ILFFKMp
t3rftsoKSdjk+BrWeV3NnbW4REX8uQ28oqxeM5WN9UiXp4mslGHfsRu/DuXe9rRo
GSUcSt1U+Wu54MHgewxaVksuVixN+MGgKo8G+R/1CA/ADsOQA7P4dFL7KQE5BfSx
NBUbyCgO1iBZtZgedagdWp/7ZH0yKGdHavja/oBMS9uv4X2uIIugHF+TojzAjIKC
eqHYnpiGiVcsCraSEDll5zkoT6zm/iOZWZDfqJqmkYiX8RjUfN+kh2nsgCKOk5Oh
2hMWhUD627yaj9bgMxyTQ8tOzkvATOQC9PNmHNcgoY9UsYkShy7VGHXMwH8adIyq
sCYG7cklo8pOagmEtVrNKXFL8J2cZ+rxOTlNQfhRH0OYuCGA2jW6lgBTr/1kJZwb
eHjChVz868HomNRI5AJ9za/zZki40kE2dqO/gnD3c3LtKHVSgC8nhCnhW7H+wITf
89q0p+8Pw7Q1vyY7+81allB5FD95km7I8ZjDXwip1vyoRIreZbPfT5EDbMGuFSsp
VkgdYVWDxci2t/yMTPSClH+kGb58w6f2oJ5H1/CrU3kl4Z4t4GbF7vxJByqvJk3x
Sl+Ul97Ii2QgSJy8SSs/bkRiPhcGazACBtOwF+KTls9kGPygXut9+HlNzTDcFFfQ
QRC523+jzrfx8s07dPfXK46CxbYXQHWL0szJEwJXt6o2DNxNXc0SMVdAJl21EXF8
5GQRXhZgpbJvj+0/iT69H6xjY48hOTESSmdXGo1xvq4qD5BkGxz5MZ/L1WtOYimj
2vhrHpwLxTBoZiQHa7oVAuiqVk7yb0FXOTGQk2b0bRbCJKDTR1N4FxNcC33gRBHX
caG/wa2cI/V/wKvaoP87BqiqLMdNsiNEMt2SYoJVSp24nMRvLVYwYF97ZDnlnkwd
LDAoWmKG6sNiHWx9lQOvIpYRJLy8DxbXzLUeG5tt1DENbbxnMmSuaIKZYzdPf8f3
mTvL8X9VeE6SINrEvltV3/Th1r3zoHP5jfYrMin3kvhS8Pf5F9XB9nUlsOJ4dgAY
LliswcEjxpsJendDG3phK4Hs31hylkfRO1go9FivCPSXmuJYtM0N2C1GiQ+72j5v
qm4fhh33Douom9EmddNaFS3bF3pxaK5cx8edZHvCFRLOHj8HNsSqrr2NsKKtpU0v
BUdge8EFVURUmUjGFTEVjM6zv00wtbsHpdIU3NZxFcQvK40s7LJAkYqs85cHl7V6
JMxL0zGEYrVmBFPcYFca3t7QR9W3Ppt7ft1A007FZ/dq3qrbCXrFI95+MBCYxOrt
LOD7Jt4NBKhr6l7XyCsaYLCZbmqOh+Q51XMzThhft169V3ZFE13u0WtLAMaOwzIl
dnIEpg5tajABZGqewkfqOFVncag1jH94Y9190P02IoWSMhpo61hWPtE2FOjoggNm
4wPKK/a/l7RAkuCQLlF9PimydqXyTM/PQjuGnJ2OHX0fJ+WadHw8HgiL5RVNPqIn
SAETqKYoWAG12b2nI+jgPNokT/h5F/f2V1NACrXjNPwzgRRdRjoYPJg9RNy6kMCR
Q9OFe96BAluO7CP2lj+RQp870OBRxTS9kTjrXqCZrfLBSNqEH9AAg/VvF8wxsiow
dXYpFSg1y4CiXhz0PIowoL5HekL2DAu2QLUJNrMdfUlE5mfBfg4oTLhYzHfxq84i
HGYBs83r/tg2aww6UQzpgwDDSPTMj+XrcTrHcm5wvxr15A9ACdXsUYx8TBie5vcW
u62IZ9tdo/iCo/UEUT66Wjzt5IzJV98EVcSo8xk3jPSS41997kYM18i28GDDDJ5P
dcXMKIhbM4KyFy+rOHFiR1tP6jX7oZ54iDYyYRBqlR1nefAWWGt6k4Uk15VLhl/X
VvxXzrG4LGp26dQNb4BD03Ejd7eSTYabSzOlFMl6ygIi8krpCnmoEqnAgmnYtVUJ
LbkWSGSno5SuJmCJUo141KI1XS3iTpXSbCJoodrXEYkAv7BQ6j8y4lAY2BasJ1qz
Jl9P8xlCIME1kqLDRhP+XTYrsIn//ZRnSbRhoqUUxgk7ySKEBPkqIRyISEMuBE7h
mduOCagbrezEP9RQBeB+ZQ2/q4FNExzpamF7YNOVpgCP58aajF3ojsXBCNI4JII7
xh2ga6TCcIzd2NL7ucIfazh/JV3+G3/IKYaqY5K8bZigLQYOAh2fliDrN3iojVqc
yUDDlgBfz8r//wp/BhaDrnGAfUCrICjenn7O7tPp5YlInhVHUM2vi5negX3gLKWZ
3L82j/mz8e7HgT1ijaHEy88hr3aastKEn1LsVav6buvbZemQoimCXIA05hPSdxi3
BZXZb2yMeLIgme7Jwfljv7POg0hFoyTkroRRJGJPsgG56bQPpnJnWjW0Sy4HYmXj
geG5Kt+tSRAPsis/cj1a/YZumwPxUhBnusvLcTASebFrVPuATn84GpfZllMUMYrM
kv+9UKNEjBTJFF20dtXi8SgORRzi/VyFQaGKCSp1TFkscNmrGNV2Y1hWyg2XZOch
5ph67DjU56SPNbXES3W5YZzWPh9W7FZwhulZVquWuwOnX0ptKn83TrTdf6xugoi8
V6rPJP/HRHNHHL5B5VLMsnlarfvQEJuje1J0pqQ9kY541W55UOWIyrdE5GjHA+UC
16u8R4b874jyN3+GX0LaByCB75RnZwn51FQQoiZK0DDQc5YLtSi1dZytvImy1wCo
rBCkrsTfYSPU+lG3mQqc9YCPpBh8EaNds1O9TYRNRcmBgTna5EP4IlDV3ibFiwMp
g+qmNxeeul9t/LW+FyRCyJrqyUk22JlrxNUKPjV4FcO4P+oExneeZp1bbFucL4UG
nt/Er1lh2Lm4eyNpcxsH0WOWo7VFNU27ZMan+uDWlmAuXgAqwGd0NN5Qv3iDlezA
l+iXB6cysd0Y3+TSVMiQL9cesmw3j4e/eK5BSfGySWRvWwA/yiJdRwmogKPPu8Cs
cmoOHiECaGZPytQEn8COLdKzcV6ZvZrPl5QjBG/g8rab45pRldYfPNaZBaErD2Uo
/5YGaRcKD16R8Jb/ui2FlXHG1vwTjuYJn3yGnHA2FbyZj6Dx1JyVN0svwUbGyZuH
+LPLkAW208hQsI0814kfr3gIKWRdhpk1gD1cM3BRO6k2oNngzz0h93hEcZnRdbiG
U5gLwWjxgkgQj5SVd5nl2Lkx/DvtputHnk3AN/l6ZIoQ4DdLy8Y7xf3sSpMgesFg
iai0Qr66wLjJ4ov3ua3/v1Y2wc77avN7KtSx980NxqendoS1tLWD3CNGlULsZFrg
mciWPIIb8gxI04cV+cH5zvGEuBmwTT5pKRZ+hcJ/GI/dllc4lb8Ws+5YfcbxMxyV
XTYhSUWlXa26LOKWBDYrBCQbgljycXhJAjCdjWe+WqM+Jeahv7qcqE6PybX+C9W5
rknzxNiXyKsrPM3zR2xbU/x7Z3Tb9vSs9virpZfKmq1kTiWvf3KVf+a9mYiHTaTn
jOHqtCO8D16afDBZDoH4i7dpTZ+rBh23bkg6ZrJc2ifXS9cWDD4NIkDYWZ1TE/hI
0Lh4Qk4+kzdtXzXAjSDNvqkTgoNzP1UHFquDgoT448MqOhFFZROZUumyL3xVbDKf
+KdDZSmGMbUjg6qE4ZSBuHgqHz5X0W04c+YlIns4Olc7vDuYzw18bJk0bUJcRKHE
Ocw+tbzy7MH0ruF8B0fMd89vu2PQSGBRHR7Grbks2ii2qegh2eSv+4dyglOE0VD/
fjsUpnkrFXnyHe2LfnUE0m2sVasYEfDR4XgZoEuKzepdMRMZU0BdGjN/wHoO0lxg
Yl8af8Smj3yVOl6WP0bylVwRGvYvaF8rISkxLDBq1VY5WyoDW3ux6uWgo9Exies9
y502iarrbjC4kUB84DVG7a+LzEr/CR/0T3Z5PY22sh5LYtqb20Xd5bjDqvz7XrZl
ncUtkTrb4Jvlsqgewp4oK4IWLK8eHN1Kq7ONMJz28iwK1qX8yKmIsRUGVGgXdmaw
gqip25V7JbpwdkjcjoSXsuoiYt1QajGMZyrC6FtG8whwaHE8WnfXo5MA2TYmIvw8
aW6iLR2YL02HlZjq6XFinliahkRw4BU0Y+xdiCvoO42VRWqzMOzIGMihZTCA1zVA
GxpUcUCl0sACJozk9oNyuhQyeiks4nXp/AoMnrb76mxIIu+VBQxlirx0ssBS77rJ
KiJpEiMbdW+WtsQQlMe1jI3HdokaUHAsEgcGmzs9BZYfhHmsEYJ8JLnkry8td8KQ
gaSHlYOBB8aPIbnaTXvhyBcap7mY8qNVY/xySVJyoU+uuZwjN3KRo2ra8bMjoPu3
/13S8ubac4O1X0tJGGhkNKOPNHB9UxBZFNDNyCyrM8Ra3C5sBdchNH21NX+PfSBv
FMDKwjxK80HQzZaF/cUmZOC6gFMOGRxZkh2zwIwi2Rl3UjgScbsJUN8/l27O+bLw
YWSTGClLh8J6Amq4Iux2vmSMClv+vn9qAeFMLCnAzy9XeJZr9JMwcFZLPSCUiyXQ
I2Ck3r49Kn7Nd3wTx13HAvjJPeq9enpCwmip774mvSjBpW2HGleg/LtPbZLc6l+J
Z7rgo3Ec3A++Y6zPntKVRUr+DNKNLERu4Tv4D82wu/i4ZNk+qvFkT6Uwgku98xfq
tCCvFTi+Y+YvFnvir4E5tz8eExXqh0mouIsGNF+et3Af9OWPGxJzLuIjyfiXsQDf
LmeKxdDd1O6o4IGnbMTLJP4L9Wmu87ElTgqr434l+iOj5DJwXi/4STjakhGlu5UJ
hAQyHPO0+U8v4cfo9k9KLH5jnjqiyX0Z4rZlUplw3sDgPlIulFmb9x16qutk1EQz
6AO6xdQVvf2wYfc9/3Uqvt+BsrhyPzxA83N/sJ65i9BO26iqMIk81PrsKtjwe1He
4yrf0xBuEb0FpVaS546SCrabBQzljWSYXmeGyvUFA4EK03C67NmISrxHEOMAHul2
/8JtU/Vngzm06ckEeJIIrvsSd0g8gENZtH1v8P82s0IVOSMwzQuLe0SfjvRRF3rW
j+CSbk/3/86jJFqWLPFnW/yAqMLlQLAa748Ep2BwkUJhW381JsiWqukVSEo80e4Y
jtmmxAU8sOm7A6gsM3i9r3uNCxGmygyT4EqOe968vpb4Y3k8/5MYg6RDcX1Qbzpg
xKp+HHjG8xH7KG/jIkU8t2W/2Qir2hVUecUOJWh31HHOalCsYfF0WHrByWkiBrRL
eCHy9KHGRPebDDrpHxWnQ8BGIb7cgHxAgrPRGS/CMggIPUhWJWfNcBQ9a1HLf5UC
dhDzAzBsEWUg2bNlqoCA8Neak6LHebzw5f0pDU+GT7s52qR+jeewd81YqUItp/yk
I37Er+VBRfQiVCaG0GYX/5lSWvXexb0dshaFD9iCxsdo6USQjjfIdJphkiT5BA0Q
PozmLP3rijPrqEoCeigc5SSkn/9MIY/TUc7KI7uVK3t5TnLMaueXr1Raf3VHMSTH
rYOYM73BFm9JeCUAlmzYhMbAUg8KvGg7HVOno8O5cjulGUO0n4B0J2ohTCvhS5SW
SlbQmwWqD01e2qsuxlrrwFFmLQCrMNB8WRSNWWtmqIAe4e1iF1pr73c9RdeZDXhb
zI4xEaw+HO0riue4gJFUWK6CpATn6U8mkXDZeC78BnUY8dyM96zcqnO6sSQgxbYc
uNvUID7ifnJv9cWyoAsBlk5a+THk6Pfse0HgwyxmLq5cXBca9/PMzW65cJTs+mcR
iUkagR3nkj8CiWqT9HCdZKHh3eAEBICDOxdD5FTnOBTGXkc5RojWBDXBAOCdveY4
GjfRdFUXH7Hy0aNnW8pepGROWSQT3ps0zK5iCX9TMUqcxYKO5TigPvDa6rVd72Xj
DWkYMxKWz5yZgl1QPxMIyqngTW+evUs7JvAI3xTV5jPxXORhGVbrGsyTkV6o25xv
qEKkVkZtrTA63pXR3LVJGnSM1/KKs0xPZky4Lu7SxjGmvk8ZjQDYDy0n8RaUBp2c
U5xW2DYns6QqWBdzOR2bP+OA40mibxsCvTbhtUQ5UEYlE1bIUVBAFvhyTDr6/iJI
fHe/08AADLbPKm2IWAP/jjTm05jMYnt1wMZ7gRgrM80El+YVkD0Lo5T02WOOzhC0
SfEhflx7np46jc1ifLVX6cR+zipxYNLqXkPRI8Vgl9WtFAwI8w82rQRw4u5UUHY9
4bfa4/lxD7I23LLBhQk1ibl++JxpZWOS6RXBcsNP7d5v/pTewwQXziK9AFa0o4Bs
qCiM5pohPhXOKfrfSzsqgcUqp8W0ZsTWWwSi/zSF5XiiZRsmNm5hdIzC2YiW2yg6
f4a6fwUfIDHJVD7M8M0AAsH3vGbctkE+rsFiZcf9+d1hU5iRR2vfj+Y/HcT3rd/e
vhKV+gAaQ+8O0qjY5i9DI6UOR5KLWgDLE1ZkbD7h7SkdCfpRSV4b1igdTxHCiiRL
qyRtNwEwyWX6BJodzgoGVHpBYVILiTcE3jTdZjNBZW4ZsKwS2bOGR/rtnqb0KNdU
TFTH/yB8bKv1oN06V2aDuYOr/KKgzQqVONqpsL89+PjFqPCqf39iNEfdJ0XM2B90
uGyqdMCJumfjjg46GrXAqUH/T2amoRd2UB8kbrMjZ6k72DSi4dWRWLBUSPH6xt2K
l6/7wZY9g0XzRvA2ggNHI7VnLil/umULo4Y3Wz3f0j6g5groeoSHdKTunR4xgHvA
LWdfDwkzoTcaBIwSQ8VJZAJ2y6kElC6Ih5XoW6wcXO04MQnljbATs1f6n+d/u/8O
vsSZNdJGfbKgrzcE7a3RrYsdnjJsYBuoR2QZOyfB3wPPrmwtR9s/CpepQ+hXFDaE
4gjUbQzgZarmUwNJvhFvDII1R56tesvQ19mhcHoflTAlmt6iyEjexRIBXFnLtZXo
DyzaocmR4dgmVMxVsqk6cIrv5XtusMt2Sf6geOVSXX3wUsHb2orWd8YAfTpuLbGE
MnwrS3G2qlyTGDgOeZPPXPBxxhvlFtZ7O6sK5UDtBN+1s8IxYwS6D7Z0RKOU7QNu
cTZeKAX4ncDg5e72DHhIqTGTs8YYdHnBagsmynbf+cl3ON9G6+apBC6AbOTopIor
/pDm0aIYAvVBuU/mpvRT/edFN9tHs3/3SC3pBra633DA+r8lQFmrm21g/k6Bfze6
W3242YuUs421z/mhsEVJF9XfYaiSh44ktxOA0PYFKlDHeV6Hu6yCm5E+K6JUyecx
FrBHgiIBLE8j9kaAMnPr+k0bgwIE3McCcnTck3gIlgnNkNUBw7/5faSdxb2eDseL
Ti6ORnc9XbijiNPlhr23eCsjSVh8EdQ4T/WZFHRQrfxPuelKDjdHyLRs+GcJMPlM
ekGwUsi4Hs4HiufgQeV22kjyhsL3uTV8gX4YWrR4UoBJESe0jJi71tPQWR4wET2f
moVTVwobRtdXBW1Za/1O9Q/NbiTLy/z6/BGuwNmFeaPhuCBG9q0PJwXpX1k291k1
SnSUBwSaAYvRH0R81DPBTyOxVt3X3fnrDA5S2oX3NQcm09hDnUeGfIRFvyr3jUik
vn2JDsSqCrkaSfWc0Gq31Mq2jIWHYOLgKqzQuhlm75RLZGwYy3S09eRfpQzOwd4e
F52mPIBDuEGgGwz1rzuDT1rgTACIPQScyE48YTfXt1CeqPs3aRgXFGaJZNwrl1HV
YSj2y1iZwrr8T60OEczdjusNiBedOjD8J90ZgkPyuaMVL9oqRp18W8qZd7OHKvL6
UHT4OZ5GQuHKCpYDp7NXMezsNN/ty6j7EKClvXoXGr86hMx5EzZgb4dYGWEq70Du
PYUI011hJgd2w818RWaFD5FONhAFWV9msCGE0Y8ZUdEoe84ujiHyQNkZOiGH48hD
hZKYMUcdhEce7HV7y7DHlK4BFrHj+SDJfEpJs4VUWoIIrz0nc2QW/0BbY0ZpoGV8
YjxPz7AOM4e+eKrCPABQT2nunCWSwngw8AzEbp+dUtQ9b/Oq3SAI7lrC20Rw2ZmT
JQB5G+8hM1gGrqspE5hesGdhBmhVNGX4VRuO1hOTIkSOPBMx5GZwpUUdeXK81Zig
qS4zDIsU23UE+JQEWu8crL8gZE6yXF/eUlVt5E+D09BPv+x3Z52yE3EdqPaXL8V2
W7qCFJp55cDManWq2ZyYjHQh8z2NTlT+cd62o3/h2yihJQct1maqyhdenjiYts+p
LAksFSvCwnPHIr1xLoKgxGqqu55d53KLEc2Y8K0gE65qervsP4JlZFtwf16Ap5c9
4CpGmuzgzm468Q46p8kKz+vqMlVYhJXpp7lr2sHSd50ovJDKckxCG5OYUq7umdhQ
ZwXUtj4ODoTCQtgWHUOOILfYbrIwsJHSd6Q30YOfsfpiEp+luuzPMEnS2C1R6hun
u1dbRfiFpV/+lVNEfVj4k50OMmKtdBfUvVkYt6IUxvCnm9QJbMnLOo5glN+BDqFJ
S97h6GGdgZ7njOl9UABzIQsOA/9ATH9ZSpoHQ51Bug64gUNTw5rtVURC7Q/Khnqe
at4WUKOS4cPXR3mp2WUVWYQrjoOq0m+5pnfYrpKTfTyvyE/ENcuAhMC9RrKDeNdD
n+F/9pZWlfq8qt4AuU1jV8gYiw98sSJsxthyjAbaiXH8C94CxzkUYfkE4a80XXql
kXSds2WqYSYc1xDmJ8Y3M2b9y3/JC4AP2PMAd3aojxwpRP63VJwZCZXBkXc2QBVf
AKfQ8IotgZzcSdTQyM/FvGEAJw9//dAoz5Zm7xec/WnVFvCKXVXRnHEJ+bFFvPSC
0OHWwQpOpuUCRKWil9mmsdjwpQglP7aobAoFgdfk9zYlH1RokbjDh0tzE4oB9sDd
BTZKtZwemrymJIx46ZfvnBN4TSE432HT6ooczT0FT297bY1tmWmvDbUnlGntA4Qf
3I3dMCG6pgXAJObdxj/UtFxC+lPilJNdYX4q4xPsKVzf8dHOYk1ok2LRGP8Jf4eo
jN4SPl6v8xlkpGJW3oZtxzd1sXd0YYZBCHF4bJnsobOXk4RdWEugPPBbhMXa7APg
Sj6cDfn2SkKFh58RnKp81zuZxmYhV7eAGG9Rz+gCv+XOKRq4zqD/ZnKMiJNMTA6I
vhRr3XVV5SdlG+aA+TTERR2kKYF+yYPY4s+bgLJe7RbdxaziGzFz40lTQYgkDmGT
wllOAZr2dZmw0t3pk13Zn6Iqnz2t9SsiehUfttsRa5PYjRrll7wYkvEmhss3h/X5
3VaKiFN0yU8DxI9/DuoA/jWoK0PhSF6Zz6O4wbGJOVhHuR7nWkFZL3BwUWvVQ2Vs
PP0U6kcReNDTNIlKjjOOuzBusmdXir87pHdy5EjmjdZb5owSpA5MSJZcCctO9/os
q8Gbv8hnDz6y9J+3smhAm2RzWqLu0sKCuU4ZTo0L9K4BwBlEpEc3ddA+s1UtfbJV
uQD2xCtU0JWXmJdY1AYBbWECCBS4bdFKwM7KhTmJqAFnEnnMpxkeYvSidu4y9u6h
MKR4B1ZOx5M/bfPKREp7fFixO8u7KoIjD3QvnHDvf5Uj8VWP6J2v+saU1G+zjrSk
XUp0NuDVFfCbWUFABGOHXDIxJEDv/Sy2yx1D03YgMARq2ip4ZKp1LDt+Phxzd64j
q0Yjb3ElqsdHwQUiMxWxdBLxGb7Iqecln4rin1Dq+t/bnaJA9Um7AGTMlmwOBE51
Te1fpKeWOnMmgP7f2WqXoBDU/eK2FLAEQsr8gt1FAm6nqSVfxqgykl0dWM3etNYr
6ZmAjejajoJfjbWIgzg8uZ2Vt9Fo/O0uQYe/FRqmHUYuiQmdj6GBXFjvuuWjPFp1
o4663aazYnF342Ea+3JKFxgHaVC5nvb5ytSYEhlriYMnT8/T4iyA0/tRKheL/+aB
02qntKO6wMbMR3ur7QOoSrLaR/1/yFj+XR22s5C+EJNMFJtPKwHJ+BJ14KrhuzkE
AriGme5JoLsNNqVJSJ0imO65TrsEQvzZoIIRNCqMj4fWj7aL4kBatuZ2XERFOzY4
QkPBDPI/F3MxgWwocL0DLAb/PMvxNAKCaz9EYjGwBLTHPnk4WppZvPbayTVGow9b
xTijEfWAMJHaqrsu+/qsni2hr2WCETerTaA6aBTFcCUyoWZ9WXz317cAk6DLJpS9
vIk+8Uxf8bnjriu/AyQdjbM2XrNJucakZw8JcXgJ7Ku7aIREO2DzvkWzcioR1R9K
lHxaNrz/JnzJfYeqKa9FQxbfLiJXxwNpjH4sQfcdTuqmXchMqACwswm136rM600b
Pvz+ztMqwG30VCRz4btgbKOTrsX0ldYc7LA/IsfzykVWVrl9qgAw9RJa5r7IFajB
TUfiAzjhJm4xJyrpJFLdVQ3umrAg28H2QVHFVWRj/91HAT8f+EvMIiP7IGfiuzg0
6qCIyd1jNCORAC4zN8MDuPvcGC0yHHZ9I+VO/xVF6CeOzbUCgy+EMs4Lqqc9M1sd
1k39cXNrVyG+/fHJCFnMQy8P9S0fDUaolg14CoHecRrd79fi8MRHLAoXB+MHZGci
6yFK/44H+VFx7DA+I95S5O9jXrOrRgbEJITHVe0vj0XOP02x4VTL4A7+TScfZCle
H7/ClX+vF9PWb2oBoqxcCnU+mCpIv5cbIYAdoUGeewj7ULWelDrFcBnSMdHlwcd7
SFM+ImypYg9dDP3fC2GFUlsZmZb6vj51AzkF9OH/PPPsKDpkvML2YsQsUpNYtVhW
rbbD2+JtArmjQv1r78ltikS9eVRj4iS2Ko0y3W/XGzt2rcI6Nv1VIr+syY6pxR0U
J127ZzLrz+HEbDBoT9cjVNe7Ep7caHfv+LqEKwDeC+kEqXkvZDqYQ7BZ+vSj7fqT
dSSn/e1pKOU50lC1rfus9Dta6C4CW3wXObPg/1wXqxdeOE9v/8F05PNuRG+m3m3R
XS1+EGVQRZjDBzntgISqooom1an1Dw5/MfN1t2lxhM8VMCdVwFwuOLWkFF7YlygT
mbbItBJYRfRveXOcQyFLeo98vKkGATUorPyCLldXUCDf/T13XLL8tvKih0NywGij
kI6/1UF1VfYGa4GAo61brRszNfM6tggKzRm+ZkEMspwvSV+Vd8A8oZTJUqA6zkdW
t208peNQMYM05F8zYPYaLBp5kUecVuWK0ggcEafPrH/QUHjFqMp/MlPeTzjpHRhY
fmfsqBAzokroe1JNXoQ9LPCL7rsBaJxjpll+dO2+8ok1suGuI9IxFmKLHMn73PN5
arxXOuKitAmnKmZaQQWQ4hgiF6wcmMc0nfukxXGVIaMYHheNOgUqRKNOT2CPVsDw
m1j1iekhyy5wytH1x8vS3IYba555UfMcZBsiWZtriSdxadke9nKU/B0B2x4haopF
6213DrVR9E+dZqB5/jkGQr1NMTB23lkn7BHOb4v4vViA04bIIRJ8955fX+pCqug2
0DC4Z/1oF6sV1TVT2AWSQ7TJ3D5WyfsjgxLcO++W2624uE1M/QLOa6ls2dgohW3w
ys9MpRzs9nuqUef1n1BOZfLJE51mGeoxvxm/wf3f2QRtd3zwYx7JeNqZYJeVebBY
TdNKSwvoNoQ5r9bbPZFg7fCHQI8c/Sp1WniHl2nJMEg/JyktW+3gQCFRrnBl+iyh
Ky5vdMrji3bynbU9rAZAY49XgLFKsUBpmxYp0tnzGzgvtgx5yy7d2Sc+wboDr7W/
qzaoYhXIFYRLStf4YOhTFDu34n7BqYaiHECFAdCb/+Z7Aw1LMyA+kIP9F4VfB2u7
TIWA/ENn7UDXA5e/2J4Ec/vu/JhzqkM6I47kbRzhClEXrteDXeYb9d3DnUdso0gn
1rr/oLnQMOWtuU/p7f5i8Pg7bq8CKfDtQ+rD4Ww570kl2jO789k7ZXKXx6epMoAy
3/gKqOV76OcGygk17bfFIAM6XwtkwfeD8Vv/xjvJgO9zawJNUXiw+O++d2ElCIpt
62VqYEUX0Mmv069Z/pJJSYrsxsWOiQrlJt1ptirmlqBG34BhQ3SoYpjoxzjnuQLB
EL8qqfwuM/ITceV3vp4zTlAEQcx3gSoT9j1g/0uEp69YjDUSwNKTOV4bIksQqxsG
Vlpk/XMhEDAHS83PHib9VYTwzMNftKNdCCU1aL7984FA3LRrapTLD16JCgmLNBO3
zr/OoE3+nsVZiCLZW0BizmkBQHpcDdKrP9X/fxqnrO7Axy0WbAxlqbub5FSp6OcU
fG2XETE1+iPZ0e4qsjlRneLkKVY33LcR5vUywCuAK9A3hGoXXbFoI22v8EVC5ulp
rmDZNp4Sib+T65iRfIcm4f4kVRL5XHyHAh0vAtsEsI54H6E5OAGLqkYynRC2lBhZ
hjqxWabY58rtDNeimjrrlL6qxoMxjfgaVXgxgCotwfcuf40vhE0byxINRYSgPg2G
ji+2Ebdf58QDNChGjpRmC4Ji/Rq5bPiKMUZv0SrVTic7LzDqoBcja0C0mYnfwVZV
g7fZJ/6ADKEr9zSZTCWK1EoHnydayn4ncgnWwVjz0Rrg19fgkQ3rFUmTMox1YaFz
r0KKCBl3mmiqshVNRy/9eGpUO/HDrO56FVSaP1MPiu7k3qIPJMwP0u3YH6woinzr
+rhJr42Mc/Uo8rE2sclpu/letglNqqGzekNO9PLnC/+ah5Oxzemnn/mXoVr7fJ7O
dHTwSFGtLdFsc/J+cssJU/elFMApr7zyn2ouzPhsIsvJSJt4F2kZCOeTy1loavwD
4iX949CuPeMOP/1hFCmiJy4Yo/OO8p/OTmc0ZjbshlYpVmpAUMv2mPpvcx8Ph3cu
UN7kUkF7Vg3UXgq0gRiOqrGfms1tcwWkPxXX9Yhjnu519BXhoYFGUZNruh4uWXzb
ewIxcci5gQgShi0lADcS1Sc6Z0QtSom7oHzfCZh7BJbRz0vCB7BMiAEEqjsEmvwZ
3YEKs7gkt+Ym2Q1u3nFgfz8OKnrLWCue3hgK8WaQlKAvac9PeswnXd2XnLzAmV1T
bnKYle9NRKj5LeLLVygrL7fn7x1xh1PiScC1xGrJOK0YYjAY1GvyrgHexx4rt6lQ
M0WZSoXH4m4nh2CcNEQarWCkQFRz2wGxcT0WfKq7BQkjTl5Dmin/p6gCBS45jks4
lW3QsBq1YYo/joPsnjFqN6DE13K78AJj24+mTBsvnvTdDqy8az8aajEN+fIflL78
Y5w4WTYWExILwdosgVxXqIc3Ue8gncjrpjhK8MBF/FsP7LLCAhUQ7cxi7bh64g/m
RhPuNgvJTIq8SFg3bpOpIDkeeJluA1ckJ0xw/Jqbj6KA3ysUHr0JrALI3JwYZGz9
XgLmdJRszbT629vYV/JlzLA/b64qD3cqaGVPwBZoPEDssXaAlCpIi8n28xeqaRc8
sbNgw/2m7bgsnC1llFoXDzPcOgqU6sK3rMcgWF1oZ//rJHMw6E/pey69EyMszQRY
EojYZTqYg0Cxm8vRlpN9IvS/QWoOdQbX0I4U+pPzn+AKNsTLMUUbmGn5Y4ipFzYz
QTVzPW+GVORTP/nEhGZ5CZQmk9USGQwy/vZdZxFsRrQtF52iOV5al0eRRsOPICaR
w2H9hhdjTUFMhqciqYn+e7UIFKEsVyYIP/lOhQnmtroahc0q4JpLLPIG8MgLqhDi
ZArFF9apXWof0CP8YLQcLdidcPuUZva9Ebue5J9TzP8fnpKnd7CxfuQUE0QtKJya
czL6AlV2SdaEN6FJ0Eu3wg6rAzirZjfdHkmm/DSk/v/8BC4nAuYkphUuZBUC/WtW
w4djvY77meQGKn0wLL5NdJEvGLTOKYn42bFr5y/u7u1SGIoZtRqTkWu4APEjEqnu
pBCK/K7FWVsSwZtRwNZ/jStdsgfK/03zRWv31SJoctbsORcxCzUzQoo5jkarj+AP
kB2QJ4TaGhaACwBZXuWnx3D91bp91ia69RUx/6wPKM61CXJBL18Uw0ladFi7wbfl
Lww377E/g1irqrvJtOkok+tApcWGO/p8u+YFWYkm0Aq+iPT1/fR9paD7NHLB9343
JttH8p/3TFLfzn6EbAZVaDFpIuq3kN5mVMhGap5wM+T6ydY47Wqs38V3CH0H7y/v
dp61P3he12b3cEJikeuaR7jPIKBA8hbP6dusnKzqy10zIviUZipRIr1YZ6JMzeb9
mKg2sk1ypn7uQsZZqGVBMTxA/NGpeBJaSILB75m55m1vCqhPraXrNF9RHoxVytbv
jyw4MxwyInrZReV5bfNYLmkOghMYImEWnOb6a4lEafWbxuw3F9Kp+r0OcArhFbMy
CE16ZfPdnxQl5UPYiuoGsf+YXpLkSGyQt+DnO0A0DOKUsE1mWxi2fpdQL5qkBrFo
lUT1tmWC2NcUdnUMY74uUG972Tv8dbosoBwat42LH8J7IAajKokbGa+1wQHdz8h7
jFjVYTT6G+9e/Qxwfqri6IjhT8hd4Z2tBaZ9AcUq1dfZGsy1B84ul5HeZS0cLrbs
Uf8PDHQFqlRbUqnbaqb/0wsBT+FQbUDhwGCQmqsGwmyN5EuXqa52TQaZS+nh+MGe
Ko1HWdbRM11ve/nX5Edmi+83EljXrKpmlyouO1iuoEWlhmphzXOXZthqSiXMHDwH
46TqIbvJ2mLDD5U07ZVrUkgNjgWw7mLKYxWisiQoN8NP66LWDOohVqfLVP6KnLTz
UWJqLzfxmJfx21jhFPDz+1AXonNUOK2jkU5Ev3zX1XaowimfMrc5Pm6XJ7sN+hU5
nP91FpiufWlVdqaAsHf8+KoYEkHHnq5m9fEFU1pXSa8KwQB1gahN1wHYo9b0AY4z
nUK7bx/F7QN9o64xsDi8p0JQ1pe3Q/CVm1QrkYlrCVFpsSU07r54teOgCnIA1HDx
BswNMKrZyrB3LX/i416MkIo1g858Lg6bVCQhsF9U7lGgpp4kk901OThSqdZ7ksrK
Q6MJzAgRLtyPHmxQBL5ivc5zkr+xt2Uey31IqAaBA4KKXDcUrllE1ruBBVTlouo8
T1QXHoPeklTkeEyR/N7MInrjo5R5INA0n+VgGp3tRts023gPOUbZ9dgP08XaK+dW
P/NbQxit7649WWxU1xqOkBqxorxP3O9C6vfUQB6XOoWOGzJidfVF+Zke7PldVr+V
Q9Tm3NTDFGbI1sTIHEpW/9drFOthBsOn6t6TqmfD3CnS7s67mvuJ3YKolHb7JK4L
B0JykHo/xKlNZ4xdLZ3KIr/X+EDr9ZqHH2XxAC8QIBPEg38WhiO32RI2QAP1TpGz
BGS54DNY2gBRl31UzcKFR/D+0nfWBH6xaoFRB79x0wausm6Z1hRVvEJSvmtMQwzk
vrXVL62WQoJWhDQc+qUiEHYwg5jPNP69/c9FyCCM/1IwLzpuP3pDWFNvEL5FJqmb
R2izvm3QLoJplwLeiuVgGLR6H+09Fh8+P8i8uxLXwr4VgnMF8UOGXQQg9QDEhsr0
zNPUf3mo3Kz/sz4hVbHurtKH7Iv+DRcSIWE4VwDnFmdYguXdg9GntTowmadMv6K7
7iNZWeEmHiB2OAQYWzlkW/I2shBSDCZguGD07JK3+FKaeXCCyFFUI0vpJYHdW8zS
fH3SSuxpCPh7qZhY3/4o4iMOhZlAy6uyBdm5lrkgg2xWFYwAakq+Gwps4zNiwEZm
OjBAoKZh/oXH3XzK2W3NGHv0TRheoV70Glr6YGevIhHumzjW8ie8raX7DisGMHl8
VBOhSQIr27o+WjVhqK9m247WI/cLTkL2M256r1ocTL7Yq7u0NQFk2Xe3rU1d8ODa
xXEAFE3uiqrchuE11wL6UNCdHkb1Vs2yaRbJ5dpkXJfDK9F6mbW04Jvh7MyWra1I
6ZeEMdkWxYcboJUnCCNwRM00jELgDrvusjp+bJsFUeWzPGH6WClRmYbVbWFJTsxh
kuXUAphcc38N5ua0nO3lEO7Z5yDgHRttqfPgwkX2ZW5fkt8cDs/Rd/kXnBDb63C0
sGPOrngfk3UodL7/Ifg5BSNKzVx8lkEyW4dfakx+5OQT+1X7Bx8qPjvwWDbZUQpn
E7beKFH3WdRx3UdFqvjCAoX9vjyvg5UqmqiuvgLvWA8kS9jPiM/yzblhNJQFa67k
5Mpu25ThWK67GjtVcCYvQckjgnYtknm8L0ML4fkqkLTnDP0mYCY3o94PZnRVecyU
Ku1eR/+kjtSzTnd/L9tNFEdxko4HZsQWzkfgMByfdXzIkRRZD3z+sRdxc7h4MUgD
o9VNFDf+M0MkJ3wcUCT1DNMI3Cl9WTC8O1VjbkTEDTJKi2l92pvoVrSVZNMQ2wgD
2i/pfzgcxVv+wDoqxgFz/QNdLvJGJ3ZFWMvxUi5pbgGOKB6BqF6aLcu6KMrMUcUa
+4mDPpCIbFwTtPYxAaBaNyn/bopaDmf7sm2s9wPMtKWq27LmhSj3YWN2D7sLpjGw
UkURezrf93y/9z/+Hn8DCZNQWDBZkU2Bjx2c2IsA2mGnFzj0m7lHqZ8GehRddj76
6vJqOO2JXJ3s2wKBCPd+ZOzySPAoS1YxXhOTbtN3KiKUKhsoEVbPhKgumAvub+4W
7nH6L9Hg76lZFawDFPB1Fu1kuV6H+jGVeWqRGulIzGjHA/g8/IqBGhTusqwaYAfm
PfECv47m+3qv7LheTyx9ePQTxZqnXMEbjC4+u2cYE09UWaA0jBNLgTx9yj83QS/v
Z5AVI1ZVYcVpYlBFXAnA3ez1V+E5r+4yYiy1aF4eDBIqsCkZeejsvv/xpGD6FDBR
c69sIjdz3JbAER9S2OuKbCyPrFkfGBuwKQywwkUVERxQzSMx+NJugpKpSRfsW+Tg
2mL6e5R00EGYdKhWIsX9NW8J+VEnLA6IURssTqF0LQwTwx/rdqG8TsJnEfW0VjWc
8tWaLw+V+ty8+mOjbM+sS9HcNJHGwLg/ynAxBkr0jZSkrduNcutj+TaHjXximwFp
0nWvaWZDIe7lgQcYX0BzMnwD8OGDAOqzmEN8BSUJzUUnBdj4ph3KZ8y5Tf0YWdWb
zbaesx0GY7FXBcgAfy+M3DeViwFHJVgWcr/dLMXkKkwzFI0Q6HDRjL65Y76yfZFJ
NMJX09j6lReuvF47tYa4MSTAPBKQWjnFmvgUfPxXLj5cow6usC9Vi+5G2QbUmr7E
+NC3krgPEyM3JJzlDY6oThu+CHBY9GufxVmo9JOeoRNvK6Q9yyxw3NHvWx7VbQ3m
ca3TmqmQ1Tb3YoLaaf2/Mbx2pDbgQXNKr3Ixqwz7os22CTxo6TbKvh1G9lG4sVTx
z9Jo7lZkpO6xnslMyCL/GvCTSdCMpyKtHFSNu9tZUBo4KHYS3mL84JK1srwnAdsS
rIS3SorzuwKjYaVQN6/QbXdU3pcy/cBNzo1+2gKgbRXlI2dG573EBMkDotg+9nij
6CD/aYvVHPe5lW8RIzw3e3/uIRvEdJlXD85GKrWolQFcu3nfisda6JQ878r5H6pr
RI2WImGDWJ7WcXRFxK+KJ7p5pwR85YI4lao3pIvfDJX/VsFIeApbl/rieB4SjoyF
S6Wk6D/r7y9V0OIrBNft0whveWXL1ZHQDNRgNWIbIj+5Z1RfIUGU7fTx3h+1T01e
L6jAxNK78ChSNZf7C3YSF6jHQSHeZY2AX7VtLmC2Y1d7SRgyWwyVYwdXc2ACe4AW
uYAoNfQK9Cbeb3HQps586mo/1KUTdw1Sc98HOxHbEpTIcrU4JtbMb2MB+LPR40iq
r+IT2U1qQ2w38X3kUZn5L42Bw/9iYXpBsBda2vkJAMgYZ7s9Cuud4ueYseWCkzLo
R32D/6A+Pv/1OHs03CeAqYfMTo+Txxq3SgEtVC7X8r4WGdVCZ5fV4m2fjG/UG9Wd
wIFdxxOuDyp9rAp4Pm/LWng3UETrgDBYKQ80Hz0NjEX8qLYKlZZX3/vdrqmRIpyE
VLbemq42NHJ4wfXUOZaAr7ey54mEFSXY0kdmDrVggXTy64+KOGTwqO16xLJaq+cC
O3oaz+DGm37rM6h5y1ZpI1XeD6JWq4nxefVP8darb5Rqw+cC8znKyepVlZDx0vpF
VqpKARzwPgp4Ow5LY9ns0j3rUhWRaDrtJQSmtR8ZvvFw9+by7O4+g4Eqh7aFvyu5
uM/+5N5ouQD0Mi8JnJJVHhf4V55HAOVzZ60iAyDGvrBqq4foVVy0GZ3NE3RbxA9F
6WvXh81LHsiZ/ClKXk+Yv8PNsvOj0+CBa8lhA29mj6xqxanK9KTRp+vpIOG8Pz2M
Vdm8PeW2IStA3tFFe/x1cFsfKZEUBP2T9Awrk905vmtwGyQEXOoiivA6JG5veYqU
c6jQAjhDCAvE/rSTqCcqJn5baI4Dl92/WNstrt7XRkH3z8e+NvhexhW5SnF+YpPs
AR94qfrZP2qmxDGkeN70w70Eze034+mtniXVIvB2j7G2sR67IEA4mUkVpgb66/nA
wtR4451OF1qCIRp6Y2zoo8/tW/AG/8AmuJz3G29wAGNfjbzoxNEXsA2SFVmieqNA
ytG5d8YtVBI/7b+NXYg7Y8kYJM6XfOpXohajzX+S4WmQbAxR2QRqpa2s+ysGwC5J
5DFJNSk32+br93C+MPM0s12Tqu9pFPacDC5Hvvz41otFA2ojFzF5O3T2DLMhRXhI
OPQUYFrIQZst11RPWk+DKwR7BGAqTLjHJpb35UvoP0qU21Lnyn3y6YFJjtRAZqO6
V1+Xt1lp3rBlEFdJjjPYQbnGQqhKcBxzdJNq8xjt1jKy3l56tvJGtHxJEtOx6o6G
1r4n/rnPytwPBgyAgKCoGIAJN167jQH51F6+tZpoCzDFNc1YtRKsLrYJb/MGxp7M
63j/G+bpiPS3D/mxaddylHR1B/AcACfgB5C0vcp4irqcdM6755MhIcSUMJ5DBS7l
fll4WoygSM2yVPxdiZ6Dofa8MbmmuSvF7OonV6GtzCO7mqh/oQ8f/5S6jqDpJSsJ
NuIFDDnL/IO+XRu+9zB3Ip/nN/Hp4ug2OE7HUpjECJGJB7n0J3zJGMemD/ks3tuf
bw80IgZ/blzY+hN+L4xmsseGjYjeaZdVRqF21s5ys1UiQynOQVJV3UPFrr+To5NO
RGRXeqQ7sv2iDATiuynhLKkq/7NMILJGHgSt/pi8NsZyacClsC7vswz0lU7BNlyl
hw20N00k2GPo7Kz8UGHd+byYXFH0T7CEjlE6aLNECYkH2jF6Dpltt0T+he2I/z/I
86LOSL5SRKF4EMvu7JN086RZFixvXzHacDqLC95pD3v4iSR93AEU7Yl5i+7zfjgS
1A0A1Cy2Ca4pUhHNgnD96vqse+LZ6tJ3MSLQaxDexFvs5UXlV32ki9ZHrNlpXgog
lwXPBJ8cjKIn8oHUst2AHHcTDdmf2woWEvpGlREau1C8Y5Iw+MUIHIBWOe7BEQgx
cryVKAMPzpOc0iShZUATLg/HUR0jvqstMM0x2dhxStYJT3KRCR5gplZ0pcvt9Tm9
Hd9ksrYB8ffqukTg3qXqe36Khx9DaSZYB+ZU2SHm6PoFzngducaGx1C/td2ikKfL
Ahg2sPdt3CNmyAZrqe498Vc/9JwBTFfjJXDJtlm39W0mQmqrcishl3PqIPy/ghMZ
RYRC02SCA5F2hIdfKkQt9V1p7rU5sBy4dnlrQqL8hLcqFLXu6w/ein/0fjIH7SQ4
1KP0wXZQFqgdGlV1tXw1IjQ1AiTolrCGg5oauA0o4jF10c2MWbFEYIoWcYOmN9eV
VTAaurrCDC/5XqsRGn8OrKazFNEH9SUEK3sWZBxCQoGBAGvRXB4i9F4NZUef5WB4
A0BJyWXM3C1ZqvmhTRLoT6/f41R/tMf7WwfnRT+zcTPcIhO05TsmhD10NA+T05bq
G8VTN59K9/HF26EOv2g87W6kLu56mEcFSt2xih4Qc8SUiyTRuPlfDmvsQHLLJSv0
nVlDI5PUf1Uyc1Gbos+85fp1rWhVvaGdj56rkiD1kCFKFCKdXMcE4j2xuyKKCHjt
nXZPM7DZDJ3jgbgqUEIjQgCoxG8wHNLBue4b2H31WfNOtms7na5De2BOm1ZNVYfb
N6exT2NqVOK8e+Pcrq3kIsv9dZ0YyCTfvVxxHjFQCKLn9y0QCIDSl75p0jbVsQsG
fjPkYiRyJsg5i8Tu6aad/+7+xLg0ACCRFCUEiYHY/YTQ6YYneCVrAaaTwRogJJE6
43/yMYVUZY13uuqNvPD1IlIYZHnSef/mb83j+g0AcOWsRv+EDQR5+PtAGiixIMqZ
eT1DHxmTSoJow3g6kGJ6tuLKQckUcQAmMoG79SfOrrakAavqH1Pcv7BMmnyo+WhV
m05XBPNFsKfALCG4IPdlTmwKM6qJPX0KEhuQ/E1FDow3vbw+K/yatiLVZ01fzRpx
CSLcAGXiPv15pOCEsaGTVViphvHokD8rywRMh1BUTGXADucYWGhSXPF2/uLWZaXK
0pKLwrK+pwx5i6DXXOuq88CQq4DO6RmguxmvIQFId5cD89DkesGed3p323yoqbOW
Ii8DMQnEudl8kV3A8gcpoyqc7H2mQ7gpOyFWKRKX+nL+LCK8ig8AIQ7ko8ni1oo2
UYm2W6E9Ix1CoqTRna6IjQdOhkNXFNF4iPg11q6Xzpmfx3f35ZvNQDzfeDWxwOX6
n0ee2y2MuN6OiCW47tddYIaIVQzwKoaC7Y2gpeE0G32ipGyuUKo6go/j0D2SQi0w
biegvybSUgO15esxKyQvO/rzd5kbl+Tzz8ucgy44S6niJ4iK7d+Py1Di7ThPLO3i
V4qA/dieII1oL7Hh2TPpBSFwHNKMnubYh0M8w/VvEy0o+g6dCEMYsgYQPepCzLyo
bwENuq0witwerSxCtQznJgI3vkvMMw6jgs1q/foREm5EhSg2gWJOH6b/O6VDePFe
3DxWQH2cl0zCQnPLlLgXsM2fLU8AHsC65HcZhS3Is3vQbLfywS42G53szuuylxC9
DpDW1gMDtEHobaHGbfg4TM2Acq9WsOeqWgTb9pVS88w153x8BA7pben3I2sUroxH
dgS+q5zBOZH7nQb91bc6F8zq4N74lo+7CwpZ9OYQTJS448PItqAh4d1HmjDT3ZQh
ugQIeSTzzGpE26AZw6FJTwXsfiQBEookxle9WQZPvC+SOr9Yr0DCqKooc1RqF4Mx
yij6TD2QVUEJr4UHcpndnbwJDTyAayVxvL/p5wYzzGf9cIaX0CkuuUIo+VzK/PIG
Jpf2FfsU+S5g24dO1YltS7lm1AQjF8iiNN8bvDWUOqKc2nCH5xNc6MYGypfeWzQV
NsojBiwOO91OzGWPH/FsQEeQ6CH8UrJCOQz16Ya7oRWR6n5Mn1meoZYtYV1vlVQq
CSfV9y5mguY7wjQp50hDmgChxk9kYXqFY88RlDOsdBIyYx5Bq3uprTC1kMFFWP6w
NUYcM3qbBtuT3Angf1yw0xFgkUAIX+eEtRCB+Uoyip5CtqO685nHSxD/p4Xev6AT
1qAifgss4RiRpcLPh1ESWflA0LUFfaWrE2OzHPGrzpEfm7CP1fJO1xA0idFy89Rw
mr4lShxXoHTU5NLhL45nJNzap33mGcwHD332lkSRR1a5GMTJWaQXGtkPM4sn5OMj
8HX38yFmlOrLJHaEXCvPS7EUoyWrijyMVa8zoG533EoasdnzUTx1HkeToZMIFyCe
y6cQesxCroyKtRXdtOB5TtfCrV26jI00zS5CwTQHOU5PWBn8YnmArpjggV/qbiP0
mcJCq+nV9FsE5O9wUX8mE43iFkBPB4LSkt9FknjTKyBtAWr2lEMBQ2GvSaagYYrR
J2rMzvEawZZaKog2Rgsefa5j6Ih5+U+N3j2LNEDqs+UP8jt4TFWRitfNE6lUD63z
wUuWH98gtBTvYIX+EmTuBXWeI/uuy88lgDSixXZM+VrdEHWoBrp0odeK4sc40m1q
cqaX1fIPXRcHu0zxFkp462kijY669MzTLPGJjrmR9CUFooZQmGrGUb7SVwn9kHnw
Xs/I3C1rzwkzJjIY1wb7rD1x+ofi+YsPq3Ng0P4SY5mKIYLzRLASPt+YCuOKS/rW
kdMsbBdIp0MsXJh00qCqsWRgCtgyh9lvKTw9ADMerGVY1GKjBlcVnVN8jH0VZxl+
i8+i5cqihNMmzCkIgNrGoVIwMX1oZUBpGDm5ofF5BeEDRnjtgdKwkiE1Zv6AHaDA
Ma5yUjnX/sZSsdo4P2oXjZ1163VYZPQ7MDI7IgF7KdSkUmbZRxIoMITKEtx35ECA
lhtP8hGmnmBLflmmXZG2SBly+wNTi4KS5hNqUuSoQNrwL5WTH6CeoBzmSdFiUhgI
2LF9hN9gBfI6OnHa5QbJP+4StY34nApeTxyOZ1zK/rcSXyyVD9wdyc0bCw/FVGGg
PYUjxCGUhIrmCL1Bqqk72RZDqNzPaM2AF0yjzv9dR+xEpxzydZlaYQ8ECTodJ3rx
6GSQjlIzKJx5dCBF7BDvXgPElMGkHDxF834QZnIsoeDNtt6R4jCkz5pz62gJuy3m
YuTC5EhK1ZNPvNZeuhRmH6ytpHgjxzl1+8zby5lkgpTXogBlS3W+9suvNQn8NxTv
WKY0EGuoJcHZ4f4EhHQ/ZJDeEOoryfcNkvDgH15ZuLdy7xme1bUjHkwkxLms/a7s
uFCbbnRDyXGuUM5DL1lLTR/zwMteIxgh/A3rxKXk824r+lVVTx1GIExeX0lYlItF
M9xdEw54DpDcymOCt5GwuhCmADrfgyUMfHRh+OsWcbZ8eMWkktBGBHFkDj0Ynwik
pB01hwOMKInwD3g4qomIghLNGehsj21NallJ7noCVuahriPa366k+y9VbVvm1xDe
+sC9tzzSpdWviMI81a+IhIqvdxDCQy/LukWLCv8OTFhUDYf/yo1v+VgCP46J7oaD
YTwO3FOD37qL/5P9/WZNzWDJY2y7Z5zvMXBfgMVvttKqIc6z6RSfJ3KnImKV7xrH
mhq7QrjguoJY/WT/A2a6W5yirxmb7t2epKPSuodGNpv6VHnz136hfRA0f4aD1fmw
JZWh6eT+sIkGgh9rZPz1Kclz2uw5tk0F1DFIQu5zqWgGYOWl/8C7MVGNBtzWrYA6
E9VcOrMcWH/bmC/1fwf0MRxjwz7r1m5eGxU538F6PwjSgFZhGOEZYdxn2CgpsuZV
PpZTs4UynzKKR0Ugmjfp558Vu/sD+VC79a5ndeupjploKAHtCoSqyYjxZcz2C7IL
De+ZN4g74Yt54TOP18NnSCl9YCV7WPeqUykVmsdFLGi5QhAeqP3VXaq3z5QZs/Nv
P6jeVzQcwNfRCT8FMNI+9zMgXP5w/i64oAD312HpdNrsRqmyjkZde3Q5Grcmdkt7
xjuxS8sTMHQCM5A4WIlmXqL/dbXcrNyKb/WYnTi06KZClM+eY++Be19Dr3aeBUtr
kj7wtFjN3LXRjh+nEjJe1mW3BS/7YACGneSYhBESN74SrlJ53DMlH4G9OGQb757o
eyaU54HoB6BtjHk8vKWI51nqOTDKwIxyTDhZRZfp+d+0KsE0NRBOEoNHWxduRGnn
yjKEo6dNFXmLA3P49Wpg8mvxXKDeFAd9uTAiS3+Gp2y134c7AzIzQCKiF10GF08J
v1DFYfN7hO6PXFmUCzeqt8e7j12D6yxigwKQrNO9NWzytiJr/2phoN5iW74fQYME
I9McDk5T7okCVtMMaNDD4dZz8bvb9vHn2iiZS6K/I+EFxJ7euJCa9o8rSwphTgJK
1ZBB2b8BQ7tw9BXfWSR0mZ1dxv5daR4uodaGtQ+X+02Vu0R6WHFLnJSqXHU/Mowx
qvla3FNKh/ky/rPlL6jBta8OI+659z4Xcz+W2ZWzNNWoNjykGwxxUe0UL40DH08Z
ZlEhET2LWgsVSWzbQ1f9iD54YqL23MD2vz8t29QfGdpdZ42XytQ3wilnWPQnc4bF
aPS+wh7Y7rmCIb4b8IRLPzHGGGVoBWTLI/ZDx58MwCny9lokzMAv6KqOdHrt1hAp
9NvN3mdx4w+Of8tfCUQV2n8znekM4Ruvhhc0xIYO36U6jEplnG7PlHCrFsiZdHql
ySUkmW77Twz4KZNnNCpIYK1cPXjkIy5b1vHj9I+CdIFYYvmgZLOVBh72s/0IHONy
Pp68QK5YjMB6S2c7+gvdK/rJyFjvzONIx4+lrRGvr89vyhat0aNfOomOiLH4+A/L
mng27Cfvb9TxMN6QHJ83cBFkpVFsARZHYAU1xUd9vX66xbUn8a/roDHpnNP3bVQj
slujurNsUkklPtv+9JnyJ9EvWiMYw735RIrevNbgUoSpPMfI7RaibiQZ8yznAXXg
MINVJL2A9mJaXJfhAcoPjhxG2L7tOY89rlnAOeytHCMe6fznIS8s8sDh/OAcG/S9
oGIOoSJ1sb09WAYafQUM+0gokUsC6iWqyKe+QLmHzwTtS5iCWR6TWQm2nQTh7+fV
nn2bpR/3iGRchfrSRWqMQmTeG8zJxwdu08xH0G5sIvSQgn9lFQOqMIafkhpxKxnM
OTNCTdyvjr2w0JMinE+ZCQRubxPxxaR40cBIkX3+UZf19Zbe6inoGJKNIb0uaCAd
ASjHXRT4Xtzp+0T28D0llLDkHVZXK0ycmKUBaVjmVs9SSlsPMM95GaohOJ4JUmcl
2LEnZEpJkJocvrT5OT5Qo4ByNtTDPqZy939GEnMpM7yZ+CI0qNKwVv8+Zqes9UmR
82Xpxb5Ac8f1Izwu8WD6grOgClDw1acNmPu7PSoyOfLWnYbxbcLDRCGnNJCTM77h
j0uZFrilf/3CL1hfl9jctQW0+puPpBsGcp7ewb20DNzZzCrorbS4MAiZbv6YRsli
2DYfNlqpyBK9YsOAmCvt/OXGj8pTiF4ohRJ0Dse4JGmGdV4u6BaWNIwf74gVm5iP
JNfXxgptrfR/gjEynIoeGoQjQrlituGnGCBQOohno9IPjckGRqFdWlmp4n44Z3AN
2H22LD9/FRx/dOh/sp1FP8XXUy39ztA73DIPeF9p+iMotaJ03Hn2eVXnABmxysOV
GW1Pb0SHR6ENZuLlqa08tk5JQaBehXiyvzaESfMMjk4U9WNEY69/R+1L6H8DXU7v
aZ1kVuUdgCQq6ME0LnAzyr+eBCRadC1EXcnktSNheCFEA5UYpCk+iskB4h5+o12j
KqQg6kdi0udb0P6+WitrRWPCLGX3ZA/X/2k6UO1NR3JqldFSDMCCYir4pEMVQCKD
cgAjYhGmzS/C2wvMGshieQ+YPdVpBB7P2PRc5y0od++O1gw43MFEnYcS2V659XMb
QvvZq4W6CEkPDDyDnsEVc0s4FhtS6Yv5OcUeiB4l1UTA961e8zZ2TnT2lORM5qhV
Cnh/tW775pCmqW8hSn/gkTXwPy0dJ+uudroTWTDwPEuMzKpRMWch2IExXoAttPBc
h6JFIR5nDI84/MlVdLzBxraEIWSyTeLz3tiVKZud2NJBBJ9uzEnATyqi0/UfCZfE
mNSGzISimyY/uBwH0+TQ7MhflW8O7R5ffpNGD+P3UblbL8/7+TMDd/j/6FLlmZMF
HKK75KcJBqSWe1oY3PTH4Ms9PvkpAeKJueKhEdr1yyA7AsKerSONTMqxOspWyjeG
Un1SvDFJZNv0xw2Pa6CdNGEbbyXZbTSjCL4uyt1ySTR5alXtnmX26EiYVOft2ou/
GRmqvhuK406u6Jl4Sdt/cNu7lavkzAPnfyT8dlFIBUczA6gqfZTShRi6neU2dAnG
9ZZpyJS0xZvoI56dTTmG2lHBeHZlmRuRfn1KG/nSeSNPTkXgyL6v2mHvVVSW0NgB
DtH4+uetFKUytQCnJTCMntBcSwvscPyfxMHE79Cc7Ji+uu18ALJL1hSowvTBDMW1
G4e3dt/uRs0eLFf3pZHi35ZNNuDrvJlWgQaCg1Imxn6h5pWMpiV968gQPY5COCfL
OiEEinI8myEKq3L4k/JBPPciLKDsDBVVbG+wONgzCo6Db58tbmnsgTvxD39BFhoD
1zQ8APAi+mrUswxS4EOYTYWvsHS+/WqtstkgO+bGj7plVlDa01hs6G7sOO1gnZLC
fS5102EFX/R7b6FvQab7fePgqrio7q4C3JCs0YSLDEHF2REJcSlPPgDzF2Fbv48W
xeExhyYogHZcwEFJE/HP7aLUox6cAQHzwcjOh1XSA7tAwT99pyYgcohH5W6NyOK3
WLg93+ekcwCSRIueOUveaLTgiX0f3QpaPLT7TUkty5GWnzwO9jab/R3+MSR6QQTF
qaBaV6mfSlpv5vQ7AyS6T2aTA43Xh2jrecyD37HXdw9fVADOUyivQF3CGS4T6l3k
W2IeKaIf+Iy4jktFyaAaISBcIgxQFZ4CjKlLB3NwamD6HZlkQN/P+DGhsokBhUnj
oIfwL+pcqNuzPYESydrwtzIPr1UX64qBHOkEXSj5NYRH6ehjX8fjRLaR4pWV6nY2
IsujPGcHPYQ6BBOK5fcpYK9Ll6UKbdLXaFefaUDOg6B8OTpXGA3Wjdkr5Lfwm3T2
woGPW/ZfxnebVBkoHbbjqPsq/nEfI0uh9bOOvYpxiOncoyi1FliX40eB0EY7sBJz
BDkA2JmhKQvDjZFOfdHO+Ey+BLzMzBVea5CLqFqt1ncBrGGjK0U1MK5tNyweTi8E
atGRQOmwKVm1i8z/U0kDXgf31i9pdQptJS2RrRYy3q1e6aamiFzQkyx97YSWMCa6
wrUlWC0tGwGVbL2EufZQK0JN+xuGP+FUa+p/XcHN+l6fqmQQsIxzZUu5ntTmECCx
HCLIj8bwEqtHwGJoK2cyCgdhiDK0uxU2fdE5le6SwOTrStLITXDseVqA+WQLdKOK
W8Vg7g7pUwoWTofKRYvFDHoLdzyXK6KL7r40TPFmxn3ndzY7ww7LfdzmPLl+IlMy
CuGZMlBM5BOlUqp1gSOQPXcmOaw1ull+VtBYNWi9/msFWr3nQqW9f6olp/liY+Kr
NkwVDvFO0PU2Adae9mAwbRbV/tipd/cUzdPGrBTJ9Vv6rsT4FXpL84nJQOh0ptRZ
bPe0aOFQ05bIfxpwkBXhVZZ1+kIa4RqyPHzM78cVsCV2C9H8Ev466gcTKUvbcnA1
UI1nSiDNJ9uAbRlJbi94Hr3ZtIo8cq35O8ORQPVX6ARt9XY5Aq0SQxQsCtZ4x22x
GeLXsQ3/tfeCMnzGOdbXGnGOmiKW7Y2r2sXXPaxedN0TNlHSODzW9oKN9oAYgC1b
wlgkPFPzM+NZPV5Rb+BIoGp5r2msmA2yittIw8+IJnwrguPMGMHaSHaRc+gcNlF5
vG8TA+Ahw5jh2nn3N+wjSnT2Q40WHYl6LK3+NAfUw61jXBOFfp9xGjbrJ+H/iMUx
8sQfVxvHOX1GxDSr20nXf76LhcNh2vAb93MqerbF1D4Z7UH3PJKdyBOFJFRQs+l2
SxUm1MpWzrsaXvMGmB4e0zyV/ghOQuC8cJX20kzdRkK6c4ug+Gflh2ZFqIxfFhCn
EYpXa20iVnV/yRXHMvKmGG+zdLjAEQM+khKbMB1zfsPuxB17DLFT3hgWuFmyNXfL
AGmNc+KOLrGHjYt0qcEnJ9AqA2+1uHKHwZrH4/bfjhdwtGXtE+OdyhRVCk8EtdgO
oFGaLgIBEX+JHUvou/qq5nnvno5hYFOekiKkj+XEF+A2xWCC+02YJQyfafgSFzuS
8JVX480Vsep4V9n4ZsoEhtQqCypy23NoU5s51GDMkGpGrc3fpF1WpFsqvGVwg/0D
pJoIMJr7WI154SeSpAx2DoTLKMh3bW/bMexGIsbQqrnKtkw9hzCM0kJDsit4PEWq
Ud+jOZKuR6j7T5tjhT/TNabsNSeFEVo+yLORn1Z6Wh2mEiiFtmrW/SgT8kvwRYrq
T8j8bNXmserrNaFo3OUvgVYxcVqsHeZuZVdlwvu9caVw69z9I6o6jFka5kRtEnAK
wSh0yzWpsR35gjznL+8lpSMNFc1mLobRxtUYOX4oEwXDBAq4+Erh09cimavN1CVB
YwPR6JD+SC3SqzY+L309TCYgehQJi35J6TapQjoI01T7JVGmpKbF44sFfYwH8Dhb
zn5ho3PCD6Fp7am8vhwASw7XDwjpbbX3ybsJEAvLfaC20CBvIRUTyUbO+IOFk2ZU
peJeNAM9e8k6NbKvyGqNXVpt1AMpa6Jmuq+VdFRUKNy9fx1nbugOPYmLooToDj/s
A8BFZaIgAWZUJVm44ZchLFaDrXTJaXIXC4Qe4LbXYUVuVbfaqcv6EKuoLqniKvpG
mib9dfxQf0W7I+NAPpXtWu1Ib8ouh1/dosiy9AXgqLswBbBfLQtA/xdi6d3HJwfT
mJT0cWOxp75DGhIKl+ATtEN9mkDlnGWIINFDQrvPeucbdZlFhm8JEkWjx4phkv7N
D5vKikMftKXBlpt465LEoAY65xDDKL8bHkDJY8ueysYr2wVzmftZWZykx5CTQPNP
IIy7GlflC6zTcf1ne3Cq3tOeeNH744Gx8HrLT2ct3Zxc6zNIwJzhjfVSy+Q6NEeS
n6sYDsQ/z22SLDcm/AGtfTKvWHRu/W6t9sF7Hk9EXBV/e8Q4Oalk3obD3Q5oxyVF
WzaVCUmvvQVvs8VvXNurdtRQB/vXWNrpN2xH//aFTOKlUWhkTfLp/Slt5HFPUnOo
yWeu+7bKn27dvWrftwJil9HASefa7pAP2nDkQ2ZyJi2rByePCAStgkUkdVcQNEfD
d1cocJGsMPnXBhZzU/yoo5/HNRrg2nHGr1JcgiGWOWzltQYuTCprN44CjfETf0Xs
hTsDlziJ2WPmBQQa8vwg8SZIU0s2xDYbmxxGMYW18e3TsWtHTSJSjFCupjsM3yNY
iLMwsKs6bhq5k6sxOQMhU0zdChisc4ARF5mxoxd+K2/sqHyQcKNVmhXIACCpbIRL
hjUOdvjd5PPmQOyZiwG80riFJXmBJDORZxjnwuLmKT0znM5PU0XMDN6oYswDWiIr
Cohcc/cDgV4k9hthZEbHK4QsJdCJ9N8rzJIg7aluM9aq774JyNv71HElmVeKDBqv
qBeTFccfgvOvvCG9xeoebKbu+dpzkaOijoZ8gAj9lgyz04R6yW7dnNVDbCs5t+JF
0Y91IpxCbMIGSp8ucgYLUDRUIrVoIVKNkOFYUYDGxLXC8AkhvFS7NUOS7mtVsChV
UykfDKWglXqO7hAvvaIQJ9+XZxebOCM1h5rOcQGVsOuSzOGCKr/kiY5h8aRjJRLH
R2nA2/HcRH2RARlIaebcSzvJuVbBtZ4KVJSzb5vBOpeopddNc1SJC8JsKaKAs4P5
Vtb6gSbzstg5snh+nHNbbIjY3ZH5bdBPVtQTJYvT5LJ+/ZmjlRWcN3KZPjDPDQEH
oFNh6S7I8P5AS3cS8Q0rTTADkQA5kV2Nu9zFO+ZFoh+D6Ve1C9ObM+4lBaMsjVgP
/NYZfSvfIjGjwWu8Vmph1c3Nf7NQx3KQ0GPKPloDY39jrB4bRAcYFEVRcUldjBGY
HId8fZWalcuml1iYHLPbquRgv3TNzH8UOAcCumVmWam3ln6NtLnAbjfh6hsgiY+I
MvKagfBPrPxkm+Ueke3R1zvDECavBbpd8UWCFRTQxar5tg1SgT0GaJ9vK7pu0AUr
WXdQEmTv6NiTHYjPruSf8VzGzd3GeMbnJA4uyOarvmLctMClMervtOIJnFmfzZBT
vGmvn1jIhOhpPZKWVFOjWCtneukFpDynfSJerXC60HAITZgDdZ7VaqtmyF/ierPW
d5qpOXTTvQ/+kg/EC7jv1gmi0VcPiT/DLqG6DEjEnYSx/yvRuW5TaRzD+KFThsbG
3L1WElzyx5wHvWtwPD0xPm6HZFBwAJSOMdx8txr2AoSHXsLvxA9afqgPyv0yQcO+
0zoOI16FlR03uyv0g1rNJAwNkCvz/nBbGb+XiTNYkG/2Ws/bJPYmZRs6I05rkTSF
YSK1iuQGeivsfe0dF7mTI2uhzeR6wfdNUs9hCY8AKScLWDbX3Ms5J8hQiLRHafi/
m78HAfyuAU9MithTe5iT57iw3CzQtmCJH9oWI43FM4y8Xe+tleYJbFrIr+VHUJmz
APw8ZupJTFEJZTRyyNECFi20+AQyc5dUKiCO+f/NPWtOxxG3y0CLOl4pnYq94hZA
LLbrLwvMlOqxEP6pfFrtWGjmAM5GtJnNzGuVfs4B1gshoV10ov9dcXBqINSMPhYl
rV/5eFxsNc4TUWMhtO/1lYhql+10OfMwYXl9nEm6ITjk+mR6v3WE19XJTzcM1Rc0
Ta8OZwqrSiDTC3gj6s0o2HV4zF0Hh3OvScnUynhfmNIaFhnxpc5extfJ7Rg+k4X4
bsSURwlefhLNd1cCSDFfu0GQmHhPv51XB60Q4tzxfgUJVnlP9TERJY1yDKH7OGUz
WpVVl3k4jHMPSGmqy9/rC5L+H6BbQGIhbkoC8OTt+hrf0UqI10KV8K2n8dHKdaoQ
diYe2HFh1ctBfMZwEZzDr/DBbARXvmPPL7H3mQ2POdAhUZqMVefHfXLU0cVmtALK
voLlGKtaNPWLg/ruRQULdFGqZaD7Cxxg7rhaT81hkvw68edoivOheEQDX2/JKSB4
Kmqni3RiyQpofUEYKW3YjwGk6JkYSnfY3jpo+mX4joyVTQx1zkdu8MSFcVASzky9
imrP5xlHoc401XR151IFBdKZ88ggBZG/DJt4QYmiPFttXxmHlzDLVCA2iu8a/XEJ
HFbVXb0HogftkqdN9dspzMf2KKmNLwiQUgiFTVYNRA/prIy6BkqY7eESF8rExiwy
pTGfE5w502aXot2D2PVSwBzP1YKSQgvP2QTnQDjyiLPgttS2yKQQ/PpwnGtQrWTL
RIDoX+fZhbDmeXN/gVva7Dt3n4I9sDNKoH2LbKtL4Kycgqv8R17RXCwAFMfW7A9z
4cuWaovbL2f4GLOCHuJURGPvuqDAgX8p6SzM2lEpUTWFKxnWwLj1Tq652/yghbl2
lKX3hVd6SMvm1N8t972Q2UaHjbF05twa0mZLP3S9i4hmWuDYqcHWj64pyrGMB04L
q8cRw1wO/TvB5o7qcthZO7s9DopX9HFo1h5I+Nn1PXnAY+3DOxB0j19Onq7bqKZB
5rt8hZpSvgBQEE6lrENGdgxf26enSZWIKEV5tndraHyvE0mr7Bo61xtnXI10hKy4
ChAVOPL4BsBsO5KvQqU7O4DHq4hr3uLjRV47D8cy4EBqhhc+zQPgheW6Trj2IgP+
vH+ZEQWTvAYAhygRr0w/9fns5yXbzIKS2yW79q6TdotSYC/j965RrcPqQgSyj2qF
3+CXOaSGvCmyKzE28SlwcXTPONwVF+jsXZjOH986xZLci9w+dU11QLc/QcSnaZtQ
utsnRQ4M3L7XV4vqLVAX0JTX+RMx2Uc0qcogxZ7cQazCKPVlZjZjpv555EfGPPVc
lbpRs7CXPeAiKR7VdXj1CeYvpf01R3c43Mja3mLFhS1Ji1ti8SQHQTUh1ZLhaQLA
KQgoUfOgoCNWxpJIhPBS47zAxZhsPFUGQJElwPq595bYzSrPuskYjSrV196wMyyQ
AnLKv+a2Uf4UGVCsalq9sc/fOynrDrzpuF/zXsuCEgETWSblOf0Q8EsjT6r6x6yD
aM0ZLX+o6M1/woyb8A7oZxgRcOQ5i4pwkW1ifxE1HBaCwrWOXGqWBBwMbKIV2pdY
8h6KIare04QzjoFGKVyC5X0ZX2JHruzCzq/AG/BFnYBv82vWkzbnbpFLpyoKEv9O
JAlHq+Eheg8YoWLCO0gHo67CJU8GYKOUTGCmfDNlMmF5vQlyGQ9WTDgmgHb7sUNs
KJlhDselITu2Efxfyg8i6CXJfkS6h7jJ1v1FBaYA9WhWW/ElMkkaYHO9i/PYq89O
Na3M+N77dfBKVacBjfUq5sncT6TiUic5rlZCi7Zmv+TbzMOwnAkRcD43/YQFk18g
3BZb479MywHdq+dzbXIXpeADvHgKSQGj3KaKSu9iDySmrGkoFPWCrmFS2L5Bo36u
iXEn2SdEF0HdKWqqtEb6HeHUUTNjBG4l3P/688DAgz1JjU+DrgINd+f5GXqF24pn
IGr6xnwwctMeIeiYTtoRYcGcEMbqCF1F1UbD1AnCneVmZADD+lR1Pb4H7Y4xiQ+G
6VPpl7VO3r5D6aGtHh6UwrNvuJax+ObDcY0HFKUpMfxgLmT12u2eXZ1MtK9ovseO
AjuVk/X0Dh146+Ny41GGLrPN3PdLnt+ryQrMtu/QDuP4wcubuxzVW+VokMs+TdNQ
erbTh6B9yj0iuU95Vn6U4GgXYe3KUdkxaEOdgTw5LHFU4DdiCqs+4NPTFAxrLhP6
xisbOatjBEo1x1nV27FnGOZ2hMgqcMNuTOitMRF2OQjU0A1au7UlHhvz1yRhTXal
nMhQ0p19I6Ego/nMpAh8xU7CFrC0mQekIloDctZ7mHIJRTM3qZBjQ7EDFm+dxdqb
C6iISVwLW7k9rWBHHVawEP9bspU/e6u+YTVdXv01dHUkvDNYceO6HVZqxOa416+i
R2LSUmDcuUNJofDKMmnNt56q4de/aszB5nF56OibS8DbIgYmse08xg6tDypyYH8n
e/WtkvFeBXHipgwnReNGfI9VfTkTVg7RJpowT7EuONTqmMtT5MhH61n+6/0osHwl
ZGZslWhLTF4AWN3ICM+LgnLL0VuYa77WyELmk2pRdybc39i/mpYXbRT7vphtWsNu
QoN1xxNymZtzr7++wYUIeKiJAhd2r+OxeK9f3PTv/o7BYd7zptT5OHxKr9GYfdTG
6UAuesGtRzg1qq4tP/WaC1r2LiI9DYljrYM34YZeEiiuY5fg/I0R/0Oa4OQuxjSa
L0Ep7kGbVUAIsS3YlZfUY5kRV/HkfPmXMMVnny0k7rUW34cn9EVZ7oHJdkcMTh+i
Q9ipt2rpUyvKLnqKKLyEk81oTCL8JvRtuh9tChwovowVMNQHQaHy16owvwxuqZbr
8iCneXY5QztVKKYcEjrgSZWzMWbwFuH6WMS+IqkVHcegRhr8+CKrTQnmkb1M96PP
j+m6h2zKet3+FT6LZXSlPIfjouoeiMLPVltIwVkhy6kTdSGz4B8tLlwY2fAYndb/
iwNc+gqOE0QGC77g/etBl9zhJoeagmRYRS4RGUZz6cuXsgz1TVZ6+YFb51vp1GBU
aJFwMWepg099IgilGA+wZ9nAeZzbMRImjjsG5uD0jy8v2Jlen6LnPuPz5rYvHZZZ
icPz0zEwl5DNcsqeeQvzI89v67wSqDA0L1aVg26RljuFeObIfvBjDQHpte1tNAz0
zlywRW1ql02aG49VGic8F2uKIKgOSHBvVVe3khcT1Bjdd0MkqlvyPJp7dw9LIink
3gMON9KIf/sb8MIVHLVJiEep+I3+qhSJ1AA22f0pI9EdE4x21Jjrlp5x3pfHoeFP
6nigDjfoV6P97XuPPMW82hXX1VcvYX+5oPDQ+Y/gYuoyfifCZVk8XNl2RMKAMXV3
/9cDyfvOygm8GLVbKz46scHC7LXqzZgttDrzXSKgFncqA7dv0X6UgOoxdkH7SxpN
AiWnRJUl//Swt9tqNhV53HKCRos3K7SiwmnNZOMaH5h/LynOLpUZGPeqCnKzHFOO
B81JK7pXe6o+fvaC0ZtvUEG4RHUmjR5BWgNZHHVMZTV212SymtUSKEJek0yX3HAn
TuyjAXTVDarhBkfwyA5Gp7MePtFpnPLMR9dTfWsL6UGMQ5OU+60iUN/9iFkPUNan
BfF+TfVo5A1mjfHXuaz38NkuTIrykQccSiwD7AU+LLQD6iHJkUqQUg/faIWrKboA
ngTSWuCrspf+Mj2f8hrYpoSqdoatMItYLqIHHaz2cLs+5bX1muRMFbfgcm+Y2ip8
+u6cD6RuvACnnYYZr/zxl782EnsZYiGn5agnyb+yLZKVkT0BzrN1ZuH9a3tpdUq1
9dEFweEmWe33vnUQqaUBbFQNveY/RZW/V3N1RsEH5iPflnKmALND91qJ8dOyABPf
vWS64AZmmk3CGAyo8Fg3RcXGPNyxhaJz4G93s2iGE6nuYazVv3QIIKnbvGsc/g1t
9DAeHcsY7lkd2zdgOIuvjV4Q9FvwORonmzVAV/vfStghhvFb9tR7M9COaSS+cMeN
uQFRyA6Fsmrsaev3mtv+qA/DFzoBcDNz1MSTpdFGqWRW5jJXeibwnkRhrVuxcs8d
4bXkF5V5+xZw84onGuLms9tdaKyILglSZdcJ9JP+hAoqEgImXZG5SXcw7zHMR2J6
HUU2JtpH3wbGP6lDzWeubKBCxaxEEt37+WaKfGm5uuji1c24s/e3B2vBrg632F81
FwDRwLScOR9M7Z45vpoEDb0DbxKGCv1Oa7AM/Y8AMZYmbMrDaET2pGL3V6t1P5jg
xhN7/8Q09gr/n2Ut6P8pi22iXZzWlR72z9lWPTWOmdh4elKmFZCFq3WrnYYTJS+6
22XqXrnrm094TJeLKrZYHdUylKmqs41pCwnHOvhVB7PhsrMR11OUKwTCeqZGPMRi
4KD4FEzlowlV9v51nMZXs/l8ntUKNE16VP00R3KtWC5L/LNcpaXreqSnQwg0gdnt
raGliBi8Sf/fi+bYd6GBUd51Cgf4VFwGxX7/4CEgI7zbWwT/Tm5SPnrQca9kSdI4
72o2OwHWYSNfHVXnO+QTT35jhneHXP6msCqsYGqPe0r9vqcuf2vOLLNGMy4xTwW6
/5ifZk8GkJrWcaW7IXeT6NG8e5bcdieVVCbhThIoHH2XGeiUQhAZjebMIatBCGZB
m58Zs2WugTmhDyuIuhGRuxpR5NlLEcdRkJukBrj6aAjny5Vrqe6OslNMxpooJvf3
SJM5FaK447A96XwAJWWzwtKILuyKYeseOXlyjIgxK5xeTIrO36+FDfTiJYMpL403
pM5mjWoD8EtWXP4T0UwflPU886AEe8S0K2MnTDa/rbS7MQ5zQnv+zRHljgUfhHam
xnBTjK5DkRt6mN+a3Plk7XdfQdDKifPEjuRgBpJ++pwkizMLw72qR/zCuvbhH9S6
ZQpTtz5NNiHpMn0J1ed/2YKKYkOh/fbmbqf7pQ27Jc/4YU8/x6eS7BG4ZD9xmm3J
AVlkvIM7Rytkg+fgSYrdHdo7rY7HI4OaZAJAIFOp7tdvHryqfOE237Vbosyv8ryc
ExChC1AqEd0goz5ira0O+FpfdIG4wN+hbIjZyItsiY8BaSHvuxqPiuFoPtYqCrj3
LwsoWt3Tw5xImGEUO9On16lhH71J2NwZ1+krSWGLv78kAbuS2cxNELNcV4AZZxl/
ldGkqpJTH7r1t7wzHYedIwJ1lEPGVsXzk9xjyj+14ybtHy49p0dHo4Hl6MyJtGdo
hDe/gSKH3M8jpUf/nAeH1wV+90RVpIJ8Hbu/0NqySVfUmxPFBhAAvjLeBWPN8q8q
FoX7B9fftU07XQz4i2tZ88D5tLAbBiZmfW0ZSJU883MYuukUbMY7UOd6RLAcQWQk
YQGoIJIjGNXdUcwRllJgXSpQJUbJoi34l19Y5MeAVq0NA6s17GSRzKIwKwnFXcum
MXZLM/RNfVd0OBJn9iklxMmFL4Bu/dVwC2HDmBZvJG68QNuWzSXV8pk1cUnoRvAy
YHAXVnHZEHhnp3gPeWQsRdYVgbmrxC8bOTzIu87Jc9qVvyPGoVSXvBOEq76H+5yH
OUJEEZsxWXJhxNZlJunxVR1dZQhWjiZzQ42Zz1r5AqFw0cz7XaQzYFnYp4kiY8Ah
1P78AqTlYpfwlQGKaBr08+avs+O5pUacjFqv1u/VyRxoEkN9WAoS6Vyb/4IOrIkY
SzQDR4Y2EVO7fTrc0su0NT9VkcaJjTVL2UcHk1rIReWZtn4KPODKHA59DoRNllpf
qpzmO+nMySwB88OHykg/bXDTnzL8SwK5J7rgi7L94e7Py0MRQYKeK3aqhze/ZURs
0okQVYgjKqZu7J0Y5usOUmItPvUoOlGuehgAzc+xaUXeEi74C5VOhkbD5DUKTEZQ
2yRgNgPlhrdTWpTcNiQGJxgomH+k8ak4V3pocS7bzNmwlIpa/ZrqxrIp6j7ehsaA
F6QF9TH2EvvDZ2hWs1YPbZqeZNwVLQ0kKjIYz4OBVrMSmuywWCKcI6L+KmubjvFs
PPxfZnI8npNaCQvosGLt+aANtBXwIH7G6MRaJq4wpl5WxKwhuKg0mVpz6XLIo6B+
WG8bNecanA/BYjTKG112UQf87fdqx2K8Ik3EovpBuQMR4pd5rfLdfj6O+fCpSmKm
1nMEumT/YPzJlVQwe2uEIOoPHU4EMhgAp1866ilFusq+DUxwEI594rcKvudC6IBS
Bfv16Wt6e8cMTuNoLkJKunyWvuhlT5liQqFnY3D8qYIgERGvAoOo9l0Epn2Jbec5
NR4hSnfQjdgvSsU3TapU9KYbFR4c2SwQp2SUun2rqfEQPUQb7ITIAawa2bL0qcbv
dI0nxLmteyC0M5qZF1JJgyh6FlCzXFvHrYmkTy2lPfdXBaawKKyrU/iSzYKeg2OE
P7D+ANeBrBsprJ5Zqos8su36i1ZTRopdsUtgON+PoG/lbSRZnDlSwHFr0saDd2Oi
52RSwhTMxWYP/lzaeUpVO4/tR5ms3hrwzkKnUxPTPayoRUsuCAcnyN/04XS8OSOv
g1fi6S7TH64REcUS8YMa6FBM7btBWWVMrBQm+nNfmhin3xYxb6TWoXQqcH3Q4HYj
3rw0IUtbzo2HVidwYHfnEVsQPLE0fsNOrhi3HiT67bY+qdSZt1/fFecrHQft+8OS
n31RQqS/jWJ8s1Kh88mzycM6r4pbrLJte9wpn6NU2MGRwcpK9Lo0Ajsi7meXWgqq
f/D16GGZcGSOnLwLbMOncC2tjwSekmsdWizb2CL6VvQnVejnaiDEhOrr5URcFkSX
zoZpKuBMSBy3/Al8JqXwIebWIH7mKDl5q9svtlmRDbrM1SyOBYLeQIrQRCAfsA2o
fsV6tzZLGgGa0CwudyPI/4eunhj5UDgmxSzly1ddHf9SCgC2bWYVPOslyBQUABFw
R73oCSSVemYNYoGJnbSjstdOm3MFiu4cuTiJmtcuerx1Lyd+Cm6g5f36CzwcESHm
kEKV7kaFD01Byq54K+hgZhxL5C1O7oSqqKtyAOOMuz+U71ZG1NErw+K8y6TpdLgp
IybAo32OTPqNJdH5FZlVfwb2uAK33cM/Qrzp3V3/OKNjUDytPQq7zB+6yE9w07yI
TqhALaYjt0RfTVZd8z7bDx+6zi1Oi2d7tJDtKxwQqSMFz8i8kTqgPueIBx6Daq3w
bwek1JPw6noy+u3A0+UMkuL3e+4PeM3Srt8Nt9oxE6n4aDBxKp7e/W94bIZIK8XQ
vAb275lZKKklqt2KT3V6eJhK2yhTqFC6KEIcp92dsXcYcXLUKqgGHja9KD4M2CEc
3KvkINXg3KtBlI4c67qZW46g4KuL6c+ddUgvh39CI4lddffcFEPAggkT2rkxx6SK
F8/trCwvXqX2ahXMUmqe4U4IMngPXLwv0Dsr7YXnuRluA5qlGrIQJ4h5HBnd8GTm
KOrdnhgsDN1Z9EBogIyTQl99/2nz+lJROL5AWpDsZMbxoFmwdN0S1Br6cLLhNUI6
CdgfsapPSFezV//SdLPGOu0GuclNQDVMAXI+gh+q6l/3qtQgU4dU9TT1qUzFKG2j
v2KNoffZRarlCMEzC1Io8RGGQT2sQwonDorb5S4YFbtOUSIsGkPijuAMu1dcx8Uq
Y0QI/lHnMNBk69V0cO7Djz5zzOfAF3sHHGvnIxKR+NosWri6QOE7D+iDwjFiBcrr
Ua6i6B/L+x+PwH8tYtVPp1UVVPGGXU6zFymggox/9ivbrunahsuUzyX4ei3jg8or
jJWo1EAwjlD2LVNReg2BnYQXoSkJ1O0hnlNouPLGOPZmgMsihigJmq5yu09TFWR2
xcPMWrwX1nVbfJifisG5KfEvHuqZk8wGY+HU5yOmVTnW25lxSww/ohFnLTjH04d2
AGa2ZpGAZGTszLAb5WAb3B2XvmJTiGJGh7xo++8GCvTeKTveb6j5oLxMsLg/n0io
faZlW1hBdQczP/4gQdAP349Mk/0sGBGq9jFkOQkoYKEcFsOFgjbZiwndXcQxAKRv
ACHeeDHBTm/ke6toVdbQ/+qczrL3cY9GShAg/ZPL7QxYE2fsLwr3Jml08MuU4oD3
w4RhdpZ3rC+zrKF+5CAsB3wgVfD4UREjWPj8qmslRnWYLY+kj+A7RvlxrIwZJph+
pel1sxJbU/uHfBTMgfhHuZje29Z8DD3BZZDN4TAEJCDV6VefDzUFtF4NQrQGeP+P
X3WvFOBxelpHaYnSLUlBFiLTLxH1OXPjFH9SVXfslOGYmajNraXjkG5VVI9REIKI
ExB+rOZtbDnTgju7iNAtcbni9H6N06ZUeDJYDcCDE901SZRvlzhy6IjEgr1Y5pmB
Qbo2XTmcqhYdA224zpQqdi0cO/nqL8OgSUJ9UPkXeocUFhxlOsgZ3u76r/pZaV0H
4vlwhJMltsHhbPEmuA1ZtFAx8HSXjYOIiCQ99z7iQO8PDWcajB32qKuMinc2QxkA
64WPouL4Q/3mprOO3S2ErBiQnu7TR3pfNEOryQM1EoxCUlAi0gRdZOw32id6ftta
vffuZe3uPicdsaoj9UHZkw+ljXvyIknCX2NwKwkYpoybLDXg2YzasCtIDVts1Kox
FEk8UoAQA/bWnnp+Nv9Y2G7QkNcPA8pgATIP8ggEnbrGaboKMapST9RTxebu34OI
4PD6LFpJROKRCOepoRBi+0PhO6VyHVBTGL8sZlK4Iq1WC06OPMPALTVD3SVGuxl3
6UxP3QcdH7llVzOYVR2LpODEXxq9MyY2KT+eeiw5K7WFE7arvJwC8FoUFxAFUWDz
HeK4j0uelf2lx/oNAtz10St5DPFycnyec+JKm+rnSZ+wlcZtRaPWpiASp7/rFcPp
sRStb82ly71WfF3mNtQb7baLXKlB+HypVyp8EzQuPJCphDJcjATf5VWv7mzQ6fgl
U8Q0xyLYeQwN1rrjanvhPQdfOHL0Eaz0safky/DnG6HBThxJYk5EUfqkoiHoGxfh
GZ86npgff2nnaioWoy77LM10Aej8tnoux0kkn/H5JOZT5Bk9lKRvJziEE1am+lSD
9ioTDLZ1kAzwUF4vU3QNzIxqLF0gM8r6/JrjYrYPxM2+Sjt3LAI9P6pxUjNZuLqs
LPSQpXndrFA3cRj2BXIfArqZ6eQ9mmJGqlOYYAaAzj4g7Z/uT4a1Xao9SlAH/Ky4
yGMIl2tbG5B2ysSPPhrtkNqPb/5+q/jzto5t/YNmpsqKRVpcljjn826U/8j90iZG
Sy+dUL9U1ytYppBlRWT5X3L2cSz3GLWc6ErbV8V6HUAFMIS/405cMdHYwAPc1PFL
neqWPi9X8LImT06NLAwHjukJ9upexeUVReCKixwfNLmCVFUmjndDeEyYYTxyIPma
FSfUJYukottpGaUqG+3vX5IpIaP811suDDWX8tqcVmCOU1UbFTk1O+2A4liJ8kWd
wP8y+yHi1V2AoBiZRFDdb9Bn9ErLcPEE6xMPQI+33B+2B7+dXOekDlyzRFuyB3YW
5HbVp4vlD4nR3BEEzauDoZSTHb1VMiFRe5G+9d9GQtOjFNIUD2HClM298ulbohJi
KWYTWFyWi1wVQyyPmNX4NB8qsB8gFIKxWWDdfJ94lp3m5sBukpTnvqWrcmdVqJHL
NYtWKVW63KsB2JPi1RBsb4lxlmrkq/IJeJSb93cMeSce9vqgQaDa0PutMgYys4zs
41eY0i0JoZlgmfSwog40QOriLgbjUQcYq8eAXYryLF8Zasq47WUxaUKlroci+dRO
ySXIfUyknBD7JbP5vIwJSHmQhHrFaOyO5jhuELEMXbm1Qsd1yCM/IlmRIME2ypGa
ILT3py84iSkisFE3VNN5NklOV/JsBMPkugmiubyBjUmnjpG9SbGfTfltvcsFotaW
tYQsnr5kBPTRE6WDj3gvu1qUOf0m9InR6VEE1LNS2YC8Mnl+e6DUSEI/ep3fa4nM
EoiO0NXzCzg+RVxjncB3XyDanuUdLZLx7MchjSqy0aderApjx/S5sWdWSFtmoD2c
Y9wTLjG+2wnvwh1augr+UhUrU8rt+nyP07jCCS/QJ1tLRySFUPwRobDLrWGfCPyX
CNg1pfTrHWG0DZ2m7ylJzoqhcm3x98Q6qjFVQ9u84aWj3LETr3DnNeZcANKwHLzI
7FoebgR14OODFDKZ7nCuewdBWnz+yOnoQ9R6oep2Us4073a36/YiKKaeWSXiu8Cj
RqUFIOdMkYyAMngzweH6JRJuEWrXAZZ3EzK3drr0HpTmpnKlLz6YlNy+ybfpJrHk
vw9LrfzAdrEvJ45amOAFk0zd3E54EJq+8F33iOGXs/bSjHUaKP6jWWAl2jZnVp9C
PXOzFZhLK4KvPFdi6wTWiLGZkvH/5K9L6K5NdXxa0JopFMWMbIYrJgPqBv2Blz1O
noJa4hcJS7SbHUGutRDjwHkz35Bs8zRdOgPV3gKCU7v5Vu74r7gk0CfQLazvGyCR
Gv2U71vC1z5cM9lTc/kL0YuHhJ1oILFmRAqDDlK0L0UK5dkT6U/Bg0Z5uYE8DVwr
ZMMURYrD7l/gCudpAZotMbAK9P7xW0qbI5SaJFH8alaGyVqBnuWwEARr6M6lxGzH
hM9lOEoHu8HpoO38vGWdQqWMRtqeDsx2EP5Y3y4S4ysmd0wgI0I7xfi0sC1MYd81
CsiATFI74PLBeQF4TpORZ2k+VvpNnWS32a2GDMwJce69IErI9RyPQH5uCc3KIHQd
6AsZR7K41fk0hmbzZN1rLEfosY07AO5JubXnfZvknJvV943o13NCLprfdlhA5ORY
/Ccg33mgJSDECc4lBgX0Z8fem+K2WcUukxfOVRJfYaNQpgTI9V4K/5aR2ksg6rIp
SPEAyqvCnkpcvVMglYuPZNfNaW5R7VUBPKDBwwsIx/2UYoCgwLd3AsJmRIKMZUKh
exg6uPgVcVNW6+mw0DMlN9DXdXTxHZndwYz/DPXQDiuUsw/LQYPi1p+1qicpd53n
p5kzm0kz0GVyYOILeEQIZXGxf+VG8ShRUJCL1bp9eoM6DSxXo/F+YnOWBD/5iZu+
inSI+dltpbFcGzrG93k/sfC2X9h5v7ays39ndg9MaWTJ9Qbp/GDkC7xKAEps9TSP
9fH9PugUA9A9VyY7PV6JmNr/a8gmF/1YkIVgeV+ytPoKeyHEKP7uTDVuBXavwdlE
foEwBe/Qmiox64zGD3+NUs8l4kwdjn0UHqqXVAdyJ5VA2ATq5niyFyBTAqkYDEap
fLkXbCil3waHr0lQK4AN9fchs0+Lpg9VsfZMDiW+BUMmIfmErMQW0jZy1rMqsREq
da2fHNRRJHN5RZO8Lf/BGQhs+GgPj8DWCh1BVpxGqf8DZlwQT3eB772bvOwZuwD6
7AXCAng6lvuCOgICryQRT5o9iu8LAGMPPxe711sdMisP9rc7BzOwbl1qNAcofhIl
g4SXYsne4sTpu0gCNXzLP+96J4k2wqCHQZCcqBqg5ozxdoG9G/ea9kWGo6Vztb3+
TAVUb+w/qj2mPswsbDqX7q8r9+jKAFElzjn2GWJeJW3DiHR1iBTbZzV3dv8IBZ2P
MMP5K+t5JElPc+FUVvKBHyy7mrE9R3PKhnxW7XO5yWJqBoNz2eapO5KFe4LtMc0J
Jm9o09MNMaSb/BLgcOfjP2K1DOhNHmbRfCUGx8vl5CJ+D476RJ2OJ+cUkQfDR7zN
yYTpCOpfM9mOABcGFGEd23AgQdqAbPbnqM/t0+mk7qH6j6HZPkzJkx5FabnrJTrK
F8w6dluDA9FNYW/8o/u/N7je3YpP0vozpiEpieamqewy3T/l/e+f5ZGjbivnsUip
YAR23AOd0IYvahz7s5JWlNJQLiyLGslNOBlJAq4V8KKXmEzpV0EGRQPailwFp8FI
O+sUf58FUH/5wqW3pK4Qd5BzajY7rUBaRGwTuzo8X7p8t5sZWpiAjDIXzyEbWx8c
SzzYMhHrwdWDo+vb4BitP3e23YBzzSwOLfwsmA6rekH/HwpA7uPOIaqGC9HkcZqa
RP3D6DAxCVKKVc3CwF03vI6GGtFmozLwPTYak1uxWMWEdzCfclF/Teb2bqPtKTQ3
5/pxS2yKRbQMZQYx9xEX5utIrQPe0iQ90gj1OO/lGOejQC0F5FOr38jEO2+96moE
4EFpQNpSaMqGTVvCOBM4tB3O1RBvKxUmf1GRCYy+x5B29dQAfW6sw6Ra/mb2jZdQ
ZUPmI8UqEbM/VL8X8JbROUIhenRiY38g4UEGuXQfkJEF/9ihMw05/kweJkKMBv8i
74FofIkXWgOququSJsYDdS9DESy/ODKO8JvJJv9Xb5kcZWKZAf3YoOMAlKObszuh
7Dk7z/hKRW53/Tkl2LeH8xurQw/FXPALtpzs7sVF+38gA6J+UKwgIMPgjv0hzgl6
Zr5EZM/WlTLvnZ3AIq+ZewcK97HjaFGYK3I9JyIF5Wm+Wap++v6CQl0xIkpMKqAd
u7v70Tb0MWdiyx1CGGgcZghrBeGOGB6yhKWLgzD+mQ9NGg67OtlQ+IbyckDup/8W
8jK1OuUoACblBA/M8sUPEE5siLnM49GYSRpW//wf7aklmVSnjvpALO0HLf+lO/+c
bDIwFShjrgU/yZoEF2QZ4MSPUxI59VsmHl0YoSIcgna4nCaqQSBk1o1cgJqnb/Yg
cIltBa2d2hSZft9M4xv2aIJK1gw3OwCLV6Y9nellJ0/TotUSvjfyxYaYA22x8oVY
F1ZDZljN3S+OBCLDo5dIDD1b/6ZtmK3N04Nj6gfAgO8yONz7J2flkzN3iOQxBCdl
tqZOMcnktri1UrEFr1dU+AYl8mxPL2PTWjMVLwCZYXLnoukuscCtCOyFilrbDRmU
wF1vJOH4xd78zri30JyXV+Jm59mQJqnf71NJPtywhXjKnZBjpyOWK6lAn6+X5sgU
fB0UnCHrEIHxMKulmUfPDvRDa8VK74mhXAoh7/q48VQqYvf4Lg8IBGNNddkY8IeU
bycHmud0cqpJw+crZaA88tPUviTk5kr8nQArlKyruyymQmDgbWun4VhJCNPB6eny
3oo8Ix50GmT/JXre8J+VlvrpmhuJRu7QHI0xHjmOJk1tWM2w+DzfGFYxvrPejodz
H1e3+53LTxRrvd1YxXNpTwVRiXSHWM0FKtaUgRzEaWdhGUhhq32NcRTneLbbmGEz
F80EBhh6t1exCBNBo0DciOBAB+hQ4UlKQcLOe2qa7Cp3v8AOeRra7XOnxmYBE4xN
0X4834qwIh9E4Kzp+3DZnQY2eC7s+tWc+FpaUvY2+OcUk94wLcvZ8/lxoIGwrZc0
3fpviQ/VxYH81dejaruPk5RicjXwJcbXScN5pu0GNr1MayNaQIjBjpVO7GUAQ438
Icb+Bz9VsekysMKbHd/MJpZizuQNJiDEdgAF0sbW6n9/MQYvovjiQFKWrTcM1M9d
Q4CBGJaiF2hiC5aFglJ/g5zsGZtxGdiDoeJOhTJeHPOYXYT0iA21qWTdhu5HnWiK
foXZY7f0l63Tl0YG0UWSxtN9oRjh+J+WYtdr06Omc9suweNxMs44TtaVRuhkOJyn
Zbbrx6uN7ptuYZKd2b/rdr2RwGbuOdhS0edv/AnDG2pzR4O7dE4oHNWpPAV5tC3y
XZQkFexv5PaFY0u7G2iYcYMbOANOvzC8tq9wLWn93Jym/N/R9p+acOzhWlPIVOLk
Zh8uwca4TOvXaCrVxxtj2vrGSYGVCHaDwZ7jCZmcCoZJ1HDUIxZqjNsdyQ8kODy2
sME8g8LEsSeor1Ph5UaXMsXSuS96ctFM5sQgAG/EKogmGay0K6Um0cj8dHLXCzWw
EQ1XHygxOBPdTj9bVh6MeAroogtU1/ftgIPdaudOOLjGEpZ1ayYapbDTFkHwdW+s
WVu0w2vxR8lOCqFiwGWsiT9RwLMShXRH883nx2jl/RCYHWLhXCxSAAnYc2glsIOX
y1Yn6cNMk0en5vYndxf2SFXtFluOsaXvMzahdUxi1+pitnw5cF/OjKrLbdEm3wJ6
zPjfrVdf35PCtIqEsqNpvGgRGF3drh4Ez/VIjL4ALP1XENLX+SDknyzamac6H7+A
0Vf+6F1jKSLT1Bwk7ozmC+hPr7GJx4fsNTYAI5QkTh5Isi9HDxaubiYjCn9XePrj
xqonAXzndjSEpt7BVz7waONtt9BZKsEcz/Jki65nV40N+wOVz9CBbR1oVJ2aY3qj
kpXAw9a6CzcPNZpHKQVj89Grwi/KEUR3FAA1Wmz3bhm59qJPLlSraOCDeOz8QEFQ
9uR+1L52GGtkEhdYczbQhVVbJA+kZZMAzSlwVudMOhAPuZMy3jKKylqbMNqagjqj
IVC5Ezn2BzLFMddV2wCvUOlg/RciAUvx6eB655FfwzYXQkKQ0SziRZmn9rokZ0J2
6qynp4XCO6IJ/tBXxHso5HUHbpe3AI3bwwc7oq9jY7hEc33nd+gPCzs+xRR4ZCbB
BwrTMGZI7xAkRvsYRY1Lu9cPndpIfpkbDQMPlVwhp2J4bkM0vZ5SOzsm+8+M1D07
InqTUeSPfiVkJsNwy/tUCm+CIZNf+OkDQbX4tHya/izx+wIx938PnTOi02DpmKIk
o2xD9D9nD+svjh/IZSxwypA/l5EbpYAVTeZ2hyOIPPP0IxFbmG2C5CuKsvqTBN5j
VbgS3MEMuidV8y116rTeNNsDx4FX+V7R/qOxVs4vRcG90X+8ZlVPzFl1nKyjpmXG
0efEEahLyyV8qicFcMb6xmn2g5ne0zp2ITyUq0QuutLHZ72mOsyR8B/al7Jm9zUL
2sbeQ8tftfTeds/LBt2bMlZbbmhePlpxLfiPmdIWNDgMLM9T1GkFcRLpqB2q2BIh
i7qa8U8QCLxMCTtXFPlkjhkONFS+d9+0bQMtUwTTq24P4CXxcWIGX2wWs1mqPp5r
XpMj/nHGqDZXNgI+O9xZ7+QLE7GnhzIfr/vHRv/ZE8yanb4edUU5lo/K8O7YdncN
sn5AqG9IArpyHWCAPyw4WE7p1dCBEqE0voyzA8dBJ2wmZ7eyosPbe4S0E0RQRIUw
kOO+E/mH7saYGO9E4fqyC9iZBd0IxBAPgXtnEzkkX2He4bZaR8mW6GbQ0tPMHqvW
lEQJsuVhEZA7ARl2DCRDAU7TQQ6NWwKH73aOUgVa9NNUsiJC8B+6QWr1GqAgXNNF
d4g7to39tEobHoY/1ySDdmSa/8h7MPZthDkPAeETenQM0t5TarnWDyABa1xhRL6D
m3x5b3OzFs058o2FmGfnzaPKpbbNyIBBXXyX8UOcq/x3SbxMXLqWXXvlAGXKZMlK
iYc1Z19YyBLzJ4AmF8zoIJXDwlD3jQ5I2H8Njn7slFLC28PUYOe0qYPIhIOmsrab
MjOpl/1pbS6RIQCcAz914EDNCjyHQj9ckjLgQrYAd1GiCP6J0lVN/3lbjdHHq+5V
GOh1NWbmTmBXNrnXLMg0/sX+3ruVe+mMJjuFlCt28qjFKCljFcB4B4J0m6f6mDr9
B3InGcCuJPHm7hhzzBJBfiyNVHj85YMsTz4/F5DH/DhHPM02mCEpNjtiKxSAi+g8
9oOuKaDoavtL9jkyTpR/5iomBKrE+G6u3XaI8Eea0EJu4vDnyK3SXUIy4vV6Xfxt
xJe2NZpm5+p91p1ZPcPxn2NwLfJIU4eeioOFx9LduuUhX0/kzvnWaQ3ZCLBAKOwG
5tWdwpEGZAEAt8R2kTZlM245duBfGMVOx4e6pGmJ41P6WHtn6KaHBL2YcLCQrJ8F
2GBe3wZoVmklqn2gG+rXGIMgNnU3YlqnxP7KalCM1ot3ZQpsEQS1mq5KBgJqvhNB
Rn5NiQpePLBq0GWGyBx29b2atAhCDLMbqkHivE1RkwuitTnFkwGIIbYR1ngFExwa
vSu4nIeLlGq/ys4BMIo8AkUXXzDz0xHzgp9Bgf0B7/I4zV7Qy/U7EGvlkDSh2UIt
1jA6Z2ngao++35ICb6/7Pa1OZdOO4roauWbEt3gXP+2aoUHLSUOygqHqd6ZB+Luv
ZUnXoMKNxVKsdv0d1pQV1k3gDZJ5TyN15bp66MRPePDd168NH72g300OvhINBZD9
j0FdtvADYEHUGGGTWaKCTl5WwSzEHPq9EJEDZ/ThH6nYTZmtwyUi5sNWbk2ZpAks
fdAV7BaHZAW+az1sofbo0YowVhFSkOs7Zw9KjX9UTNA0C/9XJL/c9wjfHS7h4N1V
OD+OYWPJVD8s6YK7442H5S8ARWoIW3OEhHp0GT41cnixip/AUl2cSA91mty46dEE
6n+1Q/j6QOH/wTOrZvazDH1VhyEVpPY++u9m8dQb75skxnwbieNIkD7BJDK46LYS
nV7eZXFGk60O/7CW1PShu2XQJHtyS4gZNTSHrcA9iar5vWXpqN95tRFsah3L2tJF
gn5Yn/YC/CAG9RAA4CrGPesuBmCVAz+nAwLoPgKtllrOOaTipoXVG8e0VvuZ6fCM
1xjEjBKFtoyMiOIzI59+FdtOogUi+rVt/1XM9vTbZWxkF+sAmeHJbkDwOMrPn193
I2DFkRvt97KQVM23bWxwKAfCvcvxyhiHztVkLiPZCPlWFwfkZE84ERhu6k3R6cbC
dsoA9DvIbw2UF86J7JpThuXuvH0Bfe2uTYwbmtEnw7799+lSKxito0asSjWg1e20
ymBVzw8N3P0d/K7Y6dGXIHYgbsCxeqjr0FfkTeORC2fNbTWhZ3XO4VFmw5voPKkL
IkGHn7L9m3Sdilr3LnBPEGAsz0mKnIjPd13QZCnJJD9zb/1cqug7Qmng/VCsxK/7
ewOOJ77sVRcquOLNj6JisFVI2QytI9KBLe71pukbfi9d54jKCAI9w9N8E4X5NkUl
jPy/y7v1JXMyeJmpj2KbNYXRTPdB1bn2VKBOl+42LR46ub/Jpk/wCGPE0uw9+fh4
bqG46CBdU43GTqRm2v8mPTzQGOIMmwFpgF7o2wS0ljmQq/2UeWG48br3zlE/ImPf
AGHgg/qsKQtv+KRHTC44YKyj3i/HjBfYO/qInm+7ckWwS3mZpKJj1GYnd3vI0JzW
0g9q/63eO8VyXFp+uaiFr+GPrIg7lBMBmwDwKgtX048iLejVR3n2/sIjBp6Kp+qN
3YjTcHuLD8uih2yB3PPHOiH1NV+lvU0+rjgvXctoEYjJv5IkOaEagg2IlMLf94Fu
nhUE7K/VvkLhK6YD4/nXaPMfcLE4vo/2GLC9FG4efkyxNf3PdZXPsGehIiV8AurM
l9fau0lCeGscpWW8C3qIJZjlbx/kx/UDX8Jla01hs4S0AT9JWmTxab9zNBa2SQD6
DNJTG/f9DDkfLhip3KOD/0c4c78Jojs0APjg37UfC//fGhgHb7UOWgtm4LE3zYU7
HOqno6dH18V7/UyMTslNIFZ46z54W7G8gEP+ombveHTXvrCYviEiQVCKh3Nw/lSH
z3rjWUxplGYlyhpzHGeC+rd73laMaZuZQe+ugsB4tlLHzkzLlVif5D/WauhO22U1
hUY4XSPyzm/TF5B57sxDSkWdJ7VweBOVT5EKLhioRCCYVd3miSFG60PgGjElTMMV
fzwyhsd7E4zIcd1TaYYhvGypLA2BKXN9Kzs1NvVJwBB/81T66nINGK516HrHJnq2
/FTTCj1h2ZZ+jwffSDGInOu8lVgSPcWu+Ww/R5j/3+9g2Hu7Su1WwUtyyO2q0UM/
MTDXUWZ3OnNwPpx72zFVrO+mRUGIUdxb9Du4jTzZ7hC07s2BrbyojjinXvTHISoy
yVyouAWl+pU6DdVjjV0OiDWlfD9Gth+MlXs4TLUKNsJHCwzWoYdc/CyzsqehXyt5
X0wkpsM7SmNutiMZIb/0DEUEKjOcMUwYq44qdC4kN7PmRmASq0SfDTkPXjqIGDDI
5u2isFv5L9zJpU4f6QyzviQUmjeqfL+yRzkcPVo75+SgwABvfWHFUmkdv9turOj0
9rNhaPgxMzlM1d0jxnWYaX6/75TLZgtJUYO1eR7z9UdaWKXC4gWHsGIG5q0/i7lt
n7UtxfDmni6u8zKuwDWk0EMjmCpNrzAstoFJw8hL3+eyH9XFX0bhkcNDytKtXERe
h2RaQnyD+TI8jhly3C5AyoS8kiHER3W18DBXtWMQaGj+1i4wd2kgBnyT5a3JNyOB
9x8foWxTxd+jQl5sIZqfHK2JiBIM2qD3zI8KEsk3TM+fJ73DSddHnh+oIb2hlZcA
fu2krSZpiESRSaB2oJ3iRpWi2fX5fSz89wzSkPVGDePrAznUqsSSaVF6e1uftl0t
DuSmeqCQd0B88ZZo7ArqUEp1Zap5v07tEQ58Rpp9bTDr1oeWr+3Tryc4Dvj+QPDc
U1gCUACLE84rrH95V8KlLXDIKjLEznPVTac/rqoLT3nU2WIJxssANhpaF2Kn4w8o
d8uVBR6nrmtvYFcQLPYSH08ZP3iyZa74iu0mv56OsmYsG+eWt2bo89Un2GguHGMV
aApAUdvszkZuDtXRVOLJEIorNMLESVNiOxuaMnlgxuSThtWehKZthB9AbQkyJkZk
teF1HnGpRNf2jdW7oVGAkDawMTSs0nOvFjJP5quqKz+WjAUZthbEjy/6OK1rIQNy
FFnyCd8RmcPvVogLHsSouDYGARALkn0xAoROrt3nZoXu50N7bfLcFqVd+BbZsnkg
LARun8h+1DIWTRncuylolcR53vA2DllH9icaNDTcjY0nLMIRqXYQHorDqL8UOD3s
Qg13SUJBHi1LyxeSuq/AwiTKOHhRW/nPPL19LjUg+JbUrj+a2sbKotOidE2+bQ5d
mlil/Zr4ndKpxYzLtKTBPcwaY5R09ZpUcboAiIZpVL6bTyLHVcUW585qZkOmIPpw
Prtdlb2RiW8Fi9idbhXo8PgX8Qo8xqs0pNBGQHscHBXzInmno5kTUSQOPsZC6Gc4
SHcJHky3s/349kk6FWl2S4U/jo42dNlSO4w9NGvQheqghDsUPyVQMExJC+XR9gjN
n8UiLZASlHFuhjGdmyDN0pvzWtIT01HR2OLzh5w+AX2hrePRJVk0jjATxhu5Z0aW
iP9pyduhMYRC5dwqH10GMubCN4P/LVox8u4fvqUHMi05WNAKRBX8LXW8JnENseMF
FtqNENlSgP+mv2fGYwPH4i8WVHv/wMnap4EmnxRNkZr50IhgFDdFGOyCmJsqXWoM
TRr3IM4eikAnr/MHpNnHpvhU5mEsPzIuZwYK9kAAn4rK3nPol14X2ytNLb3UxUtp
PflF/1qz4oDebkAoYWIycEJzt2TAJ7n1Z8gyYFEJvaFrRVshw2ZONpR1IFPgmiJU
Yxa+oLiniSSepioZYx5p8uPaLHh8UJDBPUDrd7qOs5rF1Tq12BRm4uZh8SSncsyS
O2BDweXd32jW6bCpHTo2FQxOHvYspIDW1vWvI9lD2wDOYAquvKtbVtO9PFM0VBSI
QWcruHFYZr02RumdBhfnM7TEcMXHpYra/OCacTl2pMaZgXq845c7q3OL8hkGlBcD
DXqodk6MYmWjCmaFTtK8JbgCMoErUHSYWh1ttHhAwV14Z1hv4Up5n/IiIRjSn23a
oPZy15EJ6KvGemyyg0lPlYAf8PlJkvs1zL77MjZfWzP3rLnIisOzzmDLMM5IIpkP
AejSG1KEK/ZdYyWU054+0vx2bW2a59Bbek0TXdvy5xNDGANFEUe+aOS7snYZKG6h
/Zx+MuxhfaiLvRwsJNENG0IjX7nTlmxSdYSqWpnPHAfzqyKn1L6FsTAE40uBmRK0
ai1D8r3ao0/FxKPXWyfQqYTkxhiBjNOoaGmkEIr3RkqryYSEI9Wxk9xrwCARcIYt
ixdXifdUcW1/qrTBpVAiOjqDVcBCsKylTGSDwA7QJ1zCYBl9WzWb3tlwbh+USbuu
EkZUX7KN6DiH5h1l0mUX2CHDpacPG42hsPsg35o+SHibNJWI8jKYg+5uwbQyy/L8
+rTsZrp9gxM4fAjP/qYTi8knIbnE4TX/pZpKhUjpe7NduXW/GEhMU1RdeRzf8i/h
11PI+xiEDCGufW+hLhx/CtxpV2gGRjBGNvni3XLaEtj3sQLvD90dBpaFiwWcDp9i
iPUbAaLE5wCtdAnRuX+HrI8j2LNjlL10SNlJxsTTILXneeXqHFWOIzxX7+wxqJv9
ZgjTULkd3yhrW9BFTBIXOTxM2BzmwcgDZ2DfK7t1nWoM0Mn6/F7hCfE60jeTvrJl
CBmf6p7HKIqqZbFvEZ71apw0oVwioD44nT+BZcOS1YrWRP9IMehQcIOIglA6tSSa
WZ7yf5LQdoKWEqnJ+vceBOaWcbSPCOw9Lqee66Mk0S6johoLvo9NYPUTpDepEonT
lD+n7e5s9e5hU4hNBKSj5WhpxzAi0ajazk+B+fazB/jEDhJLc+J98wf5Ozmvda/c
4OEZ8+8xPLoOyLzvlgel5vs5Mb06s9EBIc/u84J6aVJbT72GBxQsUH+Q9qv8LJd0
hxHQFBdU6NWxyITnS9yAjWbxOW7+kRjLd+lHkarBkm8F0nR6OS75qeuwFTJixyNE
vYz3DeQ4SKK5XfdtgBbt3V7r6nJOFTW2MC0CgElANF93+5wsbitIobYMonMpMwjN
yj2pnFhVZuNdQJzPvSYVg7e6iz7UeYPLDdmkDNe9tCcOvdOjVyfMy9J8rQwRsLe5
E8VzwPaiPh0z12lekmsUfL3p4MiJUcvgCBJe25J69e5PLjMGUfnBwTfsQnhAYW93
nuTBA4CpxNgRX9tVt3J08v7JdBkQBRG0W9BZ99SnqcF0dRdIWrE/68deNBqd2BgE
vc1LtAb+BKVrJ1e9B497IVZ96rXwafP1IJL4BefJZKPJG2Do18ZqzWUH7VwyTX/N
h0GoTSTAnLYPoXC/IoJs+gYyxBVk3wP0po3+94xcBX026o61uEwbXIyQitov5PMh
AtpGwXYl8lLIBMIx9Rw8VdimVaCsKxH9YQ4TTETALfUPXrCUs/fWMqnPT2Or0cqd
2D/SJSwKaTMIBRrjxQAG98yLpTx8S3RQf9051wNPRIS+PGz40paEac2Sd/6bMNko
2diYD7uEDm+2Zbdoeta2dcAQcALlxLtEkNzJhu/Tt6CaehCw466vUNp5+Z3/ZZFR
3Lg1F2CZnS+8H6ekvA1s3nbI14yRtoneEpTvjShYp26qV2YlKFA7LVgoZWmVPMwK
t+laAm9JaUY4NCT5dKIWtxv0uKRAm8tw9yFBhnkmfR2L+/mmN6dl/Bfuo/d1Ktz7
6Fqk7Ga/bCS4eveI9gfDYCW0IkLxLMhkteSJQSOSd8ZruNqdxMRpzYH1bFsjqJy3
IKB1NH4Y5r95TC6ZUpr5LeHfqlqlA1HQYFpuW4Td6Ryw27FV8Bcmi3dk4wvciPab
qQz9xeBWWtdHPHg/iv5q3oyypE4P3oWsI6EeV74LJ+xLUmBueGjUkWt5iKYs7B11
59sQN6faF69+IOqHdLBtVLjGPIKtF4RNIO4JMCuaujAbWYwUB+ognm3khqU5RrLe
la/nxEGnJukdfUUVnA2CRnfk/YdBF7NTTuQjDHYPJxiaBAITykqoduYt/VoSKKU1
V4VC17hUeN8nO7cjesahhl3MNqOI7DWFhlftBdFKwO4uMayfzU/H+NlDcgiy8Pp2
E5BmRLSnV2U38ryKzjXGZ7mCUOce/hOy7fmg2qbpel3Fz9Qrrin5/RMBsM8rdU8h
Jnj4+qh0rUB+sZ3NR8wmjc16I61gEda6xsGCqcACaRLXvazT0HJe5bGknkfqZupS
ph3Orbk4nSRYWWMbuOreMap75lXzuXhvcpVVS0UAaqFH9P5Hyj5/S8oLyXZyGZOj
04zujBPP2zE3Pu/qVJclMIyQ/c8LngpN7gsvvXgMssg2pscJ75SRYaJ3eFjoFXyP
JxWwZGmcE8eEiU+/yqvKhvjQKt4R8Scj7AHKVnaL8t21Ilr06dznGi+XMpylUSyW
aCqb7NjpCTgu/z+H5gr9GsidzZzKmEIWfY8iRrWEvSLGQhBJi94hTDxgiIh44drI
CAbV3/zmivXW59nkqJBxLJerfZopcqhrc4ydAYoQL2shhy+utw5wkgVCCUGhOSUN
XHMAfxGu/WQyIWOEdr4ptDzV0NyNc80LnqSMUNs9VU1Li3FuTwnBiqdkHi5wB7Xj
DGyDzUvW85nxm2N/GMZjU02DfIwOy6PeBXsGk0QBer0aDtKyS5gnIRNFmguGJKlV
3chl+rNHo2A3g+4HGZPrzcBCYPrWzfQwSor70NDhZJqs2cYx1YKtrZIDEr+J+ocj
UphmiThCFG+squzE8RjUtjV5FKybwqepZZ8OgsrxnZVXSz+hPNU/Id6T/hEqSrqb
UtBJECRsheOaeSeXCIXN+P4up2cOgBP3r5FWNeTFNuD9imhc3zNtDQkb0OqEoblQ
aRPr1qslIvxqyngONcClk/5vwB7s/kSrA9Kt73L6OUufq4aQq4z4jLnFfZTXmaLA
N5b4qUfuroVWn1ZX3FTBdDHIATmVaLjAqHzE2hZhn00W0K76iX8mwK3lCtnsUJgy
7ri/SRFf8dx50AiJ8GZh43zYupciOpHbkKggi9SJn6dRYFZUYhN3XcYajpHJJKgb
r1cwRKNPsLAt8UHeYRfbDJ3gHMssVbaBEQ4M4WHGhfy4Ry3G+6inL9EmJmYrchx2
toyMYUCIUW2exiaPSBm6nhGVWTVzmhPORNDQ9JAa98gqd293CxE2UAYtRAZm/As6
6gKUvSpEJwu1/9KrzJ3d/Aim4kUNUzeO8RkOtWPuC26xpuM6b3xKxOoZiPBP7NC7
lomEiBij3GUT464WAkkIEZSa+GhCWV4ObXWme6mqNCsRBaDP8EpA/xL5eOp4FHyk
YWlbuCFEgOx9YM32PVqWKH3XBUoJ7XqfzQdrTIevxrVBElU8Ud4y4hGkfbD61qwl
3vsmkXO/66WlDW2T6tblY01oBPo/ANXfuuvQOo40Dasj/AWoKPXK9WMrVZ7IpEye
LAJaVnl5CPKk2xEDOKTOpgr3dfeomtwxxW+HKj26twKlJvhmgUeYX+LsJj/2zhgZ
R7+UGXLIAd2MEnTTpyr5y+CiT2vZmWoP8saTSZnLSeVZ1/7VbsjSMYbg2uosLdP2
eUGWshUAVi9cwT4dSsRvnznT2cgLZ1+pXcvqYQoGX7MIrgkPmHD9xEV1EwMheyzt
NOqSll7y6I5ICGQiu6XJEyJoAqeGGyRgnKX42mtPUQBpLrudImKJzZLCe5Z2OwkL
BxSY9OyqZT/2avxuetWW7g+fKE2f/CvEQWHjhem59X6qscL6pB4C+3icKZsRsVw6
SErAhf+8f0qpLAO+pAS3QWM+V/OnHP7uKpDJbijUEusPxNfqdnJ+0JNapPqDq6cj
ZeKispCYKx1v6Sqn36BYE98vUlnSbNVVsdH9QHIWKNFtq5fqKpctibQ7zSZAK0IU
f2zrGwPth4T+e0uNV/gjCSxhiHGINMjKM7pVQYBnhPZHNF/sfmc7gNsorlsG70rt
fpNWHLV+ys17nqO6VprdnL+dqAdXGVPS8n+R8TnAhVq2ld2lQmmxPOYo1+ZZ80X0
QU5d5Gs/e5Jh7wjIApjVziDC/NGe7OU19EjjJvgqKR82yt5ozQZ6IC8QZ143eIg7
bdfdRlzOybFidv1rVfB7xbFNRZrvirHy2PTDHYNI0K1CdB5bCjewktmU3gvNKn7s
6xThtNveGnEFjVlZlR98cJX0DTXrMp1aHZyb18Rbb9H6ECKI9N3/SMAuyW3+SJFu
NmzJ23XXUvvF2QerRW2P5C2IP9vyqWLWNZM5u+QVuUZJ1/zPUBYNgS8W9dbY0FVg
U3lplvOsnynKLYvSpUpxoHNqkslJP2PTHmXgk4L/gTt6MeaRVhN4S/7DEB/cv/6k
ke1CVnPfkl+q6fw3T52qwTiQ/Y5iqs2oqDnukcQzA43cOPT08/LRd/m7LxNNnstp
hZT3PFKc6mAZyf/GTCO3bK+kgpMYTx2QRqKAjcq7In8JI1ukDu9xLK7Rw7Eh8DN2
9Q35RI3/DFjFEdx1ozmtlprNMjrfBT+NJiObRKpmLCE2BYStDN8hlWkl0m6p+VWp
sVBdcGtvK9Zw3vPu21Vz/bTg2P+XManErTlTa1MaUBYI91UILDJXniQlSrX7fwc/
3JQnrvaSCyzIOGlyYic88DgwfOpao3fwqc3pnNL5qTv0YHybZoximrETNQyCcYzf
0rMc05UECsJjvpz9PdUUM3qrOQPWqp3Xp2vu1L0qHftpDM9KNMew2wN63ZkdYSR6
JHwh4aKt6SwEWXdpNrOGj/POilkPJNReCl95MhEGEocNTQURRSaPMRa1BLRnpKdB
BKhaN2BrEncZ4k1xYMnqOaUEA3ilTVjgFIlXYD8sk0EdV3RDfPWvztwfpWp7M/gX
Z53x7VuHDTZCN6P04QP2c5FbwPf1m0AfqeZcXZ+cPp/4VBERV7Q9GqIAPeAyovqD
Hv6RmL1DRQzln1h2faa166WM0XrfcKRUEGb/RfSmU2RZ2NQnW4AcKmreqPXSlTSf
XGQ8uv1gkvseruq6clxeGgpsNOyLAUQpRwQe701IbhOJyQM1FvQix6CnohFT1ikm
I6YIaMIlXrWHRn/u38soxIIS9QLp9pDTRuKAZr43VNwwItoDRiKq/vG6azbrjm0A
Ps2SL9k754GA07UCqplz1gu8IKxJzNeeeUi6POmLhhS1ifJZZvUlsOtFU7pVQ4WU
kHxbftOxG4vgiHja8pF6+51mhH09crEE122j8SFnTO94Ba+LwslfANVuP9zXkxFl
+kD0QFYwzms56kRxu+3i9VSXqRMWXK0SO9WcAB/bdKk2YHgB/kTWj35M7BNcHEGq
R2kR9R8eyCt5YNvHuR1RwqUKgvmGTzLoZXzJWol0TB/ZXSAVaLe1Og5ZMgDm6rt3
JVmOpdAfyizHU27NmInrfmKj2/aKEWcFgVu3FbYkbAS+s+d4gewoB6QWllw2ub0K
CfD3oiKGxVXOB3+HM64w2xkMqERO5FW1pvUa4VK0eiGnFaEr3J2UkFqtXyu7TwjS
G846wRMiWgMdg0rzNZUQRfBEoE+CR2flDSyawl8NU+bW+gSyuxoB6J5XPYQJhCOK
IJWWicSXj+EUZEXDXUF4nnmrWoXbkerWN0idRhtRtw3ojKsPcLnqNGNFD4bOapu0
1EezWsAap8sLvrncYvPV8CWt9nMETUyMKAkjOQ3QL15AWA52vsbI5HQRRVm8T2gX
iKpO9EAQgMsF/f9dEgPeKYJHaYn+i39NcgwVDCZ6dswhUhhV5kOlk+G3/3ammjQO
PeiFo1Jo70lq9RssdLFtm6TuMZak1VJCfdPH76wUklG8lBAvQXh7Z7uoqeWn9FH+
ScAyWtcuVXepz8lBasKUKFYEb3hUmU3m+6l/puZllLduh/CmYtuL3eoMSWDHfaZk
ynQUsMWvNmKownSYo09dAEObfHZaIxio9QAGxRYx9S22J5ofhjmm+bLJbPUoBSpo
6AZB61dU8ZhgIw0PkcDf3O27FS+U+goFW8Y8fyBYPN+Q/qE57yZJy0bKjhBCfrBD
Ng4w/ahF1/lSiLG1rb2lD6/POwslp7qT8a0RLieUd2Idwur/btK7W06RvlKCpYNZ
/QriOjw3vkjgPKybSFnkGmMh8pGGEezqJSfTM/7p8FlTCxiZ+SOEZR9K8bf5pO2m
Re3J32IhQxRJl9fn62MCuLQYdfKA+JslUP75xPMhU/hV6GV+8cHZVbkeofudLwBH
4g9B67dmjr1fS7im+UJhV2B+r43F6odEKbJWzOwlvHyxXImPKoQKXMQ6diYmEJ59
G61C4qp/NbEes4I24IRq9i+zgYRVeo9vnbg7QC+o5W1Z62+kQlii+CCyIBcfpjQK
ClGSFmylUOWwHRJWpHBa2qcspEtmsZPgXJ8MeW/VZFt87BSgHE4CTceMLr9S/H96
YAg3PJAHE0pRGmaJB+Bvztx3QfumkM79B5vzlKzFICdHjAVlGNfeWVN2gW3YyRRs
7clAksIzU2C9/RGKp+Et1/hLyvCyocjfj/CDaWqtaGhB2RwEpymXq8EevxurK420
KCperL99Y1RNoG8wvts4iwA7agUMRCJM+K6Pj4qVB8nYJCrhy8DruHAOI/a2O7Ly
wfsOEE+lMfHqUK3Cgpqli6/6vbotCo1v52QGZHvhy0XFEo3SbWzOJQphZtjKMwan
JSM8Tq0l0ILSMHewOJ1aqDxDG7a7PXq61E1ag8FbUAXiGnNsWJrltmhQYi9WLTXU
U/XU/UhKRkd73lOS6Ms1xdWHVGZAQMYHloqlXWD3GNKPLOJf6LxVLmIkKm50TNQD
hYaCP4DDtpvl2rLuOi43Jt6YJzwRhrmkdetsGYrLq15QwJr8qwAXZ4QWoYrqnisF
WmiBbPTJr6XqjMyIvv6OvY5YW/XZjJ1IyK4Z+PfNJui8KktHdT4eN0EFea8/OsmO
h4DlB5cg+/iJozv+3jGo2FQrkSPNUowaThPe6QfsUpFFx7ez0O9ZFxUIWbYC6V69
foef7FfhIiHqofNRNmwT2awmSD1yB/Zkd8oRZMbYJ+Km2MG8TitSifeb3y1IOJsA
CRdd7TLqy3My2INdhqWTn1+eJIaTfthpSghj8x/A6cnt8MizyWzb9C6vsJSDxzZo
tUG2nPTHHVq/swIaukaoRMNd73CgL5JnOBEwgPLTo1QwQkzKMhOChwnL2SWWrRA2
jgRyQsXy7EQOeDk90yVelZr8cdnnB0KpGC6OMmoFHbz1UTzQhZTfs6Rys1wgV7Jr
oGLFlBXjh046xeDfynGKIFo/YpGb6pt7Mc655g56MniXjViNBTnMjijdnsSK2flf
aJe5G4XtFKV89ZlAY7SpmF+vu6M305kiDTKSrzUNl0zCxUATKcH0/O9jGNmopgya
3y6qhzI/uPWi7/3CGki7FijPAYTfcVaEdVId1EHX4ZYh+S3h9TMWgidaD/etBaYL
yMh7itN70Q9zD0LYA87ZvCEtD2TtTmyG5iBy1gzl2zxVUU6/PfrzXuCAh1UPHvqz
i9Q/fC3j0NU6qLMaaIGy2pBJh4a3mXC8wvnppQ5RsRVSEICMdrCcBB2wZVLvdaXr
d76rHgJWNoDNyt1bfaQU5W+15GAN2ZWa3fbzqCBK+o5NPHad+hmtJCN+sQcKMZMI
6RN/pVSF6mIPHbgtpdezZ7vZ7gbmx/OqO7Fl1JhOxfRUnXm/VGNyRRZYri7GSryZ
cDU270Toffq0yPABGeEoK63R4w9LNAp9I1w33egq1l21UlG8xVt3AtV3Vgepy6IN
GhBwkRYhrdCiMjW8jNOBwXcuK6t3fmojCQqeTL2wIIMp2JErTcG5g83+dWun1g/p
g1Lzs/koVGn6dnz3mbnC7cTIlNa+AsbZEQIo2DGjF+APnCAEtezj37xs6YhkoKRt
TQT9xgwFpg4/DUdJmBZ3y/pqnghlgohctaOCRmccOQ4j5thf+nqQy41jv34DfqSU
ImqkTcyzZjmLEfmJHJJbhsF6Ku9Gkwy/QnghU43+pqj0JM0/BWrShLUFJA30LFpR
sy/u1z21A/b/bA5WkjFCvSdJsHWbcwa232s0r/QOsq7mCJlhtchdqtRs0FAGQSLJ
yCB/YUZ/2h84b4JjHLhZ9uQo85tooaaALJ33ASR4EmmiVE+ZnzihTlSVQdHvr9u9
jETO20ryWGnLcMl/lJLfz4otaVY7yZx2HJGqf6NWn4V/Ht+II9xxuWGf2d6SZ8vm
DuOvNR606teBO3wYKasT26dwLqgUcQz9NgeMabI5bNLhTPicK0e46KYIea1Uyjq8
2JeFK/pJrqeGemJU8uIdusI294XH4ayvmR6e6cE7/R9A0fW6vV2gzSqigsDeKgOQ
6+ZA1mm4yoEyQA8XrsBFDjAGXb6X5ZfA3X0DOeWfAf9vxbKFIi3GJvHey2BrVf+6
z+Jl6H9F0SBuzcoAcIaITBiu+UGcTvrtvnrzuhQ8Yg+0M+TpTjtfYWj8G7U9ZN8Q
8FoTdD4s34JgnkFF9Kqb2NEco10OftwIXxQGLppOS4Apajun69Eu8jZydM9IMP6I
rk/zNsEapJsMlm1x9lkXWNneA0KBaKbGZt+qykol0Q3NYkPbPr0dXusCn0UmU/CU
SPiQh6PY0oHqAAQsmKDAZUFT7asb/gbDM20NseQH0+SRX7eRDkjZ0G5tY3HmiJf7
fY2pEFBqxSihOsbPkplJUCDo1s9M3hG8BXKgEFEA7M29tSM8+bTP327H8bWbqvbF
M/207vFHCTco7zVPvjZpDb1tY3CpnzjJtbuyzelmt6qN54yVuiW94HhocVVWpPBW
RVMzWvUppj+BEICKnZhegb8F0ZUhqVz/qjeevxejJrWHmKt4pP7rhTf9u5jgtGnz
/RkMrrzXN0TJKT22Icr/MpW3Ouo5J/suVln5xem0IFj7dkzJajB09rOtcWlf2LQr
th/ll9kicaGXHPDAfsKatOcSa5O0ssmWN2OWqd7AmrS7p0H0p64EhGjZYD+Y475Q
dIx7h5aYZl/16h1CsaZp+ZAdcNLqQV16G7eF0G/yL5hC8vu9uGpLc12C8QE83mqX
fHjRBs0gTSWp+p8yl/br3ogLNRIYfxkn97o3Ob5fyKgzodjvSFXvbrMA47zSnpg6
ItN0F7DC/kUUHlfoHe51yDh/xJohB/v8R2p0Zp1RNxIU7/003v6C3ThL0rOfzXkL
VaWqeW+WPdZ+0Yl3n34I2LMIfJgdtmTNyXv92JjHLxLB2C2ePLMe4Eo/54hCYvDj
QegZ0Cdrye6ck5sIL7wOokhp3GsYj144SNJ35+4/UrinbHzIdPHLQIa+yWWulbU/
pai6afib8ZJgyHA3CaaqwR0dbQB6jx5pKaPeM/8WToDMA50YYUKKfd1175X7tpAB
vKjj9JUO7bZLwDCbEBKhR7ak6Ry1TEa24ia7ZncEK6az1EBN2nkJwTv//INxAwol
hLPT7GKSwGtxEBhJiDgLFaLUAkwqFwf+dldwZH0frjxU8HjeddReOSemxrR25mYL
9KmeadhL3Dcv7botsnarKrbEVJFfVcEUtB31aHf+77UQe4a+qfDw+gI6w+fKTzZk
1RqAZsY6wYm5fqcuL/BT5tZcBFho9eQnjSNQ25yl5ems6C91GAZRHYSxrK5GEJfR
DNDqoA2/CeDsBa223f4hk1apABem6EfV4p7kl7tWnmCv1ansTDyJ51e9NfD4SCA2
rZ2cyprj7QshPRNxhwsdYHeWAo1SVSyoNlo5qQ1fWupuUcooyYzt2zdpfAoyIrxF
zF6sY2UtbKXFXh1TS2x48TnNxFZoRWfF/Ta7I3R1HrSQKgLSmy+Ojj3m38uGrzMR
ZAgqMW2gDcGcAYwjYZvo2ZSm75PRzRy4KdQh52jmIaXD8ZrXyJ/XqjiqCw9Me0LC
uRd3Jl6Gg2iu3SJrWBrooAsHeTswMo1IEP5ahxPYNy/kKZ7ymGZ1usMWzN6b7K/w
9WGbJhstnfQJGZSiOjeFl4wVizSp5oZR8Up38lcKsbnj3x259aIGH2hNR0Rgl+nL
7cssKvczvvuODvBiZfHPjIZ7ZIpfRP9feSa4G8HUOVOT55fsa1LITns7LucVUtA9
MeiAIaw2htu2v4MlbbernaLwo56vNfdZbbIaCgvuwKcdzSlvtpnoYQz/+whBskRF
To6uFmL2PARI01bVudgmXOLOf29OsxxoQsQMX3WPVEXe96d2zQXKt9yitY95ZSiV
00sNqf3TBGmN2tCtsnWIGSDKIAmwCiygy8mMrRLXrMK4LqDaQKY7YXvWo9kcF9K2
af2ieVSGLkhY8t2rECrMPSnufYLt8YPtvdrZYqMVv2LMjCzf3ro/zGVjB89tIVmU
I58QSk4rg4SGL8JsAM+4yUOfSmRs+LS6SBfCGn6OpBtHl0rsdBJNWtCrB30qx3Qm
zt9FDuedMdJXz3Nzp9RF1qEdmxWul0vDG+5oBRCNlkZJG8iVH3UUGz6zgZcpSj/F
Gu/o64+NwKdUr7Hiesx3G/uV7t7PTZRiFN1HNImaE0+Af2MRehjCx6XjrOyjLwW6
wKrZicKzELgtHPMVM1LbxVJK5UQFGBHZdHAv/VzgXcuV6sSTeouJWteo98abATjM
PHXvwDJwx0fny0yXZvJWwdEtLap/1xtBMtmBENcqc2HZaWJ1ZEOESlgNdRYk5ybi
dQbXuRqc49b7Ofam7fyuNrXfZS03dAOIF1NAfMXEwUGfZA4EondFHExlqYWS/fpF
6VQKdvmCVaZKH9Yv9MyfD+f2M8nI0N4OdNRbE3cFNI2p7DY8hXqEn/1vrTp4ath8
pnbI7YILr4v/bNDViK4qW2vAw6oeV+AxsjOkvEaTAB97/eVQZ+bx6p2KTpgzdPJT
uZQv+zliRVvMwFl3XmgN4pDepiJ6TSDqWBwv/ULU+SjSPc+EX1A+f1meNs0wrLua
KkLAJcnh+KTbE2YOkzwpW7CvaGokvii7Fki7U5GdsgbG8LhnYPLjhpi11QOlkH4N
wAD1VHH2vGznmDzKV40hB84WncIP+qnu1WMXeoBjNxUYyQSQSzxbIdOOjQSLbFKY
VfajEHBU3ANgRKazSur/DXbaCbyS3YfBy30XTfAP/rpo+phya0rUKPmty10Vp8QF
HGdpMM9AMU0xGbCa7PVQ2qn48rUUoM0eSdBAABCt1N5Ztld+EWoIXYavD15x1KCU
ow4nTIcXEIxGNW3+V5G9YbyDNKdz+ui1FIre78viN3EE9dwpaU/38LeYOFz7b01A
285wT4wTnXdMLUZZnZCn9GsCP/faWDjthsabKRTiAhYkb91ktuYr0CicQ0eQL5Gi
8KN6TMgg60W/xXfG5mb+G2DUT1auVVIn62MDdMtzFwTz9fNt2KFnfzIlzK1VWiJw
yPD4ihSAIyyJOH+VFsFE7NC/JkMxxcrWpF5iH3Cqfpb/RaGXN+YTy6e+wbPfFUry
m8ymgaM8s7E10ZGD6IH8sByhVJiyRAmYWebmoXirU9djusPjT4pLQJlpZBMciwMT
kHMRlVY18buHFEKb5z6DzfNscsP+PdFtGEVF7ZtYnXjISPVl7l22saxXlVZ+pZDu
LkG0zXxQghOt26am01ruF1TCw56mXlVnLh5Z2hAiZGTXjpbd4fgu7sSvkC1VH1yX
pBK5D+cc0Fq9guZa0GQToxel0fGQAzAoyG62JzTYghUha39bchOx79IUHRMDaWCO
nZpeMbge+6PskwJFm9CClBlEMfo0joVQIc7hfjVZOSWIh9rYufI720zFkRs8ZJkU
d0ajmdRGz4nd3h5oFCwkxwxLhTpI+3yfQJcqqdqeX2nGCXIaiATc746PLjnhNCkk
j4FohbTvAZdMKG+ewZuEKLeGN/VRyjDSP6uIAfJzadibSew9/qTiUGeH4CepDAX3
PgVNqC0RhymSHzLQ+73L73XIiHJOzdln2yZhMjbYbLKQunaQ9PGShRHy2re1oryS
OM2iAk36J+5XGxkt4Vj8CkjES7v0p3epsPNDN41gPjQ6sq1BSI81ktTIRdgIqwD8
NVAEtCKKbz4VWm5daug6w9vbOoOLOkNtbwe5yYTKf6q6sh0qUUJINENoZfForN66
ioEDJiYjgbxESmRenHRqUyY88u6K1MGW6CmLnDQRKmB3VAAcoDCr1qrDs0Ok+o2v
fWhegLnVOEswOjyIskme7L8Eh3f93inD08/VFJEYvB1Y3auMneaZAz8nUCVAlGx1
5ByCH44yRmPg3ZRdyRrMpsxbbFxKcr61eSKKB66LiW3oq8Bbvr5Qlzb5Lonk7/hU
z/1bBNu08XuK0cIctPfg4t+otkW2cte20FzE5g6x79v396LYV0yWYYTyha1uMA06
7Qx8dS6/N9ExkVHfAK3T2A56iJ7cY/tavyteR3DfSGoweyNCGQdy8Fts2hDTCuNm
s9kWb7WUpiPQRJqEZGeZVzGFDKYmfbCAeg68+UYlrNPA8Hao5JpycQpsQ93+8FUX
XhTUwN5HpRzIBoKwz4PuH1yyUunT32As2ynnNwY5twRD9utcosKQplnM3HA8ZIpi
ttBVZ+UTQz+ydzQjs83sSceVOh+yoLMnUBWt85Yl/5CsLO7HwUfmc4T4QTOUmvqK
jzsWgg/bbJvOdJqUo0Ry+5YJ6MxQpNlomfH+jp+q38tbyjGeZl3jojD8fLJsLgNr
B/BliIBqVs3rNJFeb5Zb+tAhcQaW/7LSSTZE5CyMCOz4CSnQvUgyX+OAzSTn3cAs
Ux/p81fB1xx7TDzqsKvQncE5PaHbP7fjGviJVIolxwzzmEXftzZvHUt9Opka33MB
rw6oCR2kPvp316/rvI914soSYvXn2CWUvc5/fhiZ7iSQb15xXEDBB02jiLll/I1c
bOY7ZYDZLUG5vAH3bYkgxBxxpJWXL/e2IU29qp5lfTE1a5DWlxqjucOwNlIDDp0g
605oFgymlEHFJo0TicUYkIh66iJJWOoLFCq6JKLmBdl2cqScvrld+gA3oTpXE6fP
W4RKomkCUGaSOQqN87um0RHd6gWxbdisE8daD4NTdxjSVp6HT+ThEn5x267CSNvp
Xdg/DdECZBtOo2sMXMxwUktl35SjIrS3iu5bjlGzJlhtflVaBWcjJKX0XMAzJenw
LGO6GfUCsdpbkOhifZokIaz8151sUqGfnUQ/r5pIAI0Fptx3DX1TeyZ9fkI2OLeD
4OOu9qAo7BjVWR0EnEAIqGftQhHGg17vK3PR+7Juva2YiyozvJSXXpP93qf60mST
SXOVpXegO8LUobfjJFVyQgL10CeMnJ668H5ur1nKYD5h0ewF0WK/pA8NCplQMNqD
xmez540hLsxTwtstf4tJtPmoNBnE3vkbQOu2nb/kH64dPnwcO2kKv/H2kRWRlg6L
FrzthdnjTSTgVKSclFM+C4Uh5VITpF/jcYnI7AjepUIzAm1aNHqGkDWRk5UM2f47
0j+X2udeoiRXEpajpKJpcvdQN4EJ/81+61aSFMNisyVOjz1Ym9lWqYqBskleFhKC
yUpvKW/VzZQtPGWRJZgIkkW0V0lUKitZpBi1w2duvV+wUD0T8o3ZeS69rnyRHnTn
ORJchg+gzEcXJ0GmFtajaO6e+RNuRZyqoMtvBEvqlCZlQ6aKRkQ7uO5QDvnbdtM3
423irN7defMZpItRWYihy4V08ffOjAj4wfFqbGzL/a/9iWr6dd+i7g0cusLwt+FA
BjE6cFdM6m2kryGqfQiPwGHYTOdSJkdV17wLc+RdujYaVcrywhG6700kWtlQBfhj
ftcQY5NsbUEr9IrSevuktLfyFiP5LHvM/wVw2UqunW/KDtlYZ3KegCoTtePL08nO
bQIH5IARh1MPiDZPFAYzYAU1dvU/sTeJV3c3Pg6BcoiFOLiZloDa4znQuqAUB1+j
UsWtxZ4y/vfCDlSVXRt+OEgl8nxkxJDfBIxkm/YXUcn+x3V+9W8/pUonHnR8CPIe
XPDQnQYcqjW8+ku5ummWfZXE54/vLCZZ0n3pTZ8/oDMFfiHt2oA40qoRTKWzReBA
qSGN3vyMqzKXxjm/eNfPpzQoCtkjroHa4Xg+0sFhdB3ZIhu7dgjxcO+U8AXPnPKS
dsfDpbd7UGTsKSLo2h9yW/bmdYe8RoCf9rZCiQFBzh3HOO5dArCg3nTNzIL4Npl4
IdqGs8xHF4zBptcaqZHfxTbo6/X29F44kNEPk5IygpSmCCbXTOyANBY7S4c2oRCn
CWli3MRDj9RONVFx8oqDjsLNVDqF/VAUKWLYhajfRoNG9sE+Q/nWvyz5p9yUiUFV
VMhbCDzqMY5kPxfwRspqWoVKLVCOIk89+h5tcIyQ0wWJtJeMvl1gsa+EHJaMn1vr
1brkjvGJ3nhxKfbyqzCT7rTNiFAG7MsgGyS3Au7WUaW93uA7xblh+LNJvxZnFXe/
A3BCOr1McZFoEOfREQOj589nMyy/wu5gUU0O2pIWuZt1eWl8lnQNIj+BzujBsiqI
YBnZFuOs62nvQyA95bu0f0vdP1Iv7Dd7BIiVykXDV0qQ1oVD/jvW4fMO6W5G5Cq4
55jH0aGUb/MS+t9ENSEg5RdrTY9JJwXMeOAvilMo6xGOgL+OajfUt2TaBYP0hffj
CO5VO5F/GeUvlP1hpi+v4wdJdbu2fEvoyaLsJ9DBAwoNAbdCU9pavDgH0Nk5xuwy
8tReZ3fUgqDEXr7p4bicyK0lqXAI2n7O6TOV2EX+aAlcC0Z554sQurPiBeRMRtaS
y4P20WrqvrSfbEiML3krVBSmOoD4lSLJTIvDMgf1qEfO0Quai+jAGAAzO/i0Mpoz
UfRsMU/AJHY4QZ4hZLlVw0YakuRUStSdkaomn/nptdRhrk1Eul8Ly2OGp2J40p3X
xcWWAsycXXhuVHZIznd9oLMPeDSdSXZgzFalUAbljIQu2BeYYeGrhQYa3BgWSdzR
BljbvbrNaO3vhmmVzsBAM9hhKY0pL3/s7CFSic9AOJJQiX/dVVRXVBHrJocF9paW
cRHJpvg0nLbFrbqmQkvluqekGTehmPqJ/bgrJgq7usgYbDppll65AmiTcTP7zfma
KuujFG512jnEWg0IujaoQQVwd3MpiHN2lsKpyiX3VxA0U5C03vDN8VxQSEmUf0KF
uoZOeXsi1CIkulxYvG5GPN4m8Aq/Nt2ErGbTobb9MnwoekyggmgJO3FsYOeM5kgg
f8mIErtJxdnqN9Cp+gzKO/dO9sLwKed4ndMTu3bnVuMnh/jdO6AmIsDf2raw2Lwt
NRkg4/xUsERnDG7kcckWt+rFeRR2yWu1p3fElYh6Ro0QDRnX4RdMNqvHih63B/ls
GjZziiV3vIAvIYeKCPh8ByWeey7M6edzPZK5kVxA+vVda4dDPnVANaj0/aq+rWTg
+ZtMiVz0uX8cnhtSv3aL2rznC+j6nCg7BrSGxUwYQ7fGtfXVPw1usNtF+vgQ59z8
g2IS1XwQdPMeDcLc98qbDCyJHg/XdElLtgbu0dqHCeUMNsjm75iSvLHRtU44BqDU
SiKuMeVsOoUxgzewyAkP2fmFeJVxKcRykYyfXv3TtykjVMSooHEkEiSAM/v3bDpc
9S6O0zqr47urDEJGnMPCbSVujQdOwLKo6meaOBj/XsuAIPWaWdgdWW57UFL3K2pk
qF2GsyD3vhJBi/QlEpYlB6FKFpDIL8OzhoZepwruo1jOrBTV5GMmKUx/IRObLpEC
v9BzswWjnv3A5NZLidRsgXSegqS9sigeucaMv95TmHsIgigaEtLRz/A3pOHpvtGm
XHrlJvZTHlXjE/IL2vY72hN1PEhdfyy7bDB+NQlrecrIg+r2oDIzoG0yCFgxGHDB
/+MNhDbnkKBFvrJcQCKwhE5FLG65EbZSXl7oukvjKuwDYA2BStB+kPv96TFJAdxt
iBrka8l3ZQn08m+Ge+lvlVWbwDlw0+1d3RZbbhUV/nXjP3pNdifsknq1FWmInT3C
DKQJd/mATOPJefdTl8DJLLavaaVo9/b3jHcfUvO0hsjmFLvhr1iu5lYnEjhVOBLW
M+mlrfHeIeyf/IPS9dUNAWwRzc92JtktO1A4aU0Da0dVKHYfP3/16u8r9hBtR1h8
mqtHv5AFWK78TV1zswFz+AxcFE0hbdwUjEWv/a46Bcj7lThD25DbMdrmtDDEcqmY
w2o3SY5zkz6/gZ4OPnRnLj8acUDphNKVtGjzGavkOxFPO961aHb5Az9QiuPEakPa
vRSOTJkvtXv4qUlFfr/KFvDF+Vqdobf4ZV1sDmQiSVpAmxo6C9XRvm4Mz3bduCHi
EG9VV6PndIyHCMKqMURNi9bByySDbkP8Fk0Lox3A2d7T441K1Xa5BFZE47ZsSYcw
bS/00+w8fryInSb/qFMZrerd7HUXiH7DpbabW+HO0xmBTE7KL+s9vJYKjGn33xNc
ziVdRqtGkTPUOZ7sum9oIIZ/K7eNU+nihjqcVeLm01oYL3uI9bHnfqLwYxYCIPwh
KkH3uj/P57FxG3YzRRXiWiSPpJMpPGamBkXS9fkUnlL5K358naAhf5wMt5eVxtVD
OBrxrj4DuOYRVyE2lmzpR7hKfnPfxxBiMIhS6IaTKDqrRe9yObhZFVVFmGykUk/S
FYmZEwOTDV5lkx/OIqEuOf+WF7O03JLpNGE+Mnx4vVF6WYsK0WS4d4zwJNwte+Ae
af/wzrM/x3yspYLqP3NPz52PK1YVKJgjyFjEPA6GSNWDPJ5pIYQetrnvdkvWh0e9
pbyu6SSOSfCe6/fWMQcFeAww4NLqkPyXa382TpF2SprR3lAxzRRnyv53QN2LBYIO
BBDaC5qvKToN3aW5XJ/Quaw+Uhv6nZXqNUxQ7NafZCL2LqBDzv0IJPoJ824tHZoy
D8jZVAP+1kpREzqTKdNxX292E5AYSZ7jT+aAQwTvY9hhz6KXdXzawry4CZo0WKWs
+WD70aqmd/GRv61H+HHTEHOF0BtEOIbHqB5DW1ZuViG3TPEqH8bGw4L3m3T+h3pP
Bj6DfUvYtC/LA4SNSL1JhMA19mIlkeek4RX/hqewYI0J942UkrKgagkgS29HS8OY
1jW8fPhao3yWCDf/OTKe19CgvQawlZynGrgjbN0BHi/49JzUW4vlCRp0s0gomaxE
PuqAolFJmpLoIeB7LB9TyLOH45ZuDF6DqZ206Y78IRkw90oQ4zL/xKeI3Qd/ee5O
bAG2IjsB7xV0OwGsKmrmbK9H3W7cKBE14vGF+63VV9cxyWuWnxjkfGeH5qRp4y5N
hh6uD9VbfaPyR5YfyfvnIRfybPbWTwC6yBRWdNmlLiJPU7Te+DfdtG2LesOn3sUb
TgwT/dKbbMPisRm9uIzbkj+Cuqx4n3pBN3QV05oU7Vj6pOCqPGq9Ui3y1fSNk2A8
qrJ+pY2SHnwj82x7UD63HuRQ90i2gNmzSdhDJ+nHBpn/96znpXfWtKdrvqEcoSbW
VoSZFZx296LGPEA1n3qM+oz0lypoHBRAQqZARqTS03cAH7WjLzPKtRtyh6WhqYGb
UJ9igdLEqNkU+mFsqR0XsOjFuwT3sEdIdOER4FDCCzX7Svtch7WMRQTzYLTxLiDT
B5KOVh2UflNqZJq1WbJl9FskF7CNbxQ/KmZGX76Xy+oyEpuYuO0ySnMlNzahKXFv
KXEGTfeu3vMXVbsaL9U0kaEf/zSiYXi353qFhE7MQLZ0MR+Dl0hLA/pcd2i9Ks2m
kXq5MNkw+QrupQovw7L3Hu/vPsMLNU8uAzYTI699TulTeZIa7s0bV06gr1zTj43U
soKehuU6i57Gxd81lkshYBTP8almt4spNfDPajKZAYfP0yUUI5hn18oGH6SO2n+D
Jdn6xO0R4ieI7ZXy4zqA//sqdJWsbkqwlZyAMZM/zEHSacWKL14x4LNsqDRqPK3d
XX8YySfwkmyuyYSF7j0jteQg59LboExgpmW8NDtTwBd++9aKEn2cx/bIfd/G577j
B8vj/1yv9qkuv/dv4qJ9BB5KMgR7W2ocxlLnsJmOsIl2Yb6sJnVIpAclJq5aAtTv
VP2sy78mzKx++5BzK+Dn1X2Z1f4ZSIMGD6GCDoiUvZdNreMNqY2XvHCFnCEPMpXr
eu97H989uYI3PHhX+jB7JZRcclcpE3DiSthrHfvJpPKI9GXiRGAx0R88XOuM82CS
KZWI9gNROBbjNk/W9D7FZxEPSS7thA7SC142HZhTXniYZRlYy5dqQ3aNpYuI08to
5amAdpzvsueKxnVg2yIXWYsQ94vxJCJq1wqG2Z4gklMjNMwMPctEXtdRjihMjSHT
858aP0mj1Fpf4vh/EiSENoGiP/xVSTPfP8SeHmipjPOJB6OJtDjprz7BHBxQPc3V
Ief8DrqFCWzpa3eZ032W3U0nmGYSdec0wsvIXdbPrcbyANT3zOBFwN1H0+rl7QRw
Dm/a0dtfEYCQmF69ubJWZINK8I23++Edc60vNV+8YlPX+QZy8OsN3XMDFsMwrJtq
7B3SOo+1xdxY2/TEf4o3s05z40QfEA8Z2A5Voxd+71jFGOP49ie3lC804mQFvK4e
kKD4rI3QhKdTn0llgeWibn7GjnadQgtAZIGb2qVDPXa6mIIIyM4EGIuZM+xEiGO7
4nBVC2B2o2q4J/k3mTQo7ioel9YCvCRpuGRiAQ/pWvsbCR+nUjNe41DSIIjSECkw
C4loYj1is9u0HFsoawrfPFPNaiplQQcwUbNVy84oG5CbUZkdykU+kMQvEhjbTm0j
yAtue1OhKZKpnISZ7UfplBiQpze4W4NVqISja5aLwlpIOwXVaZ6HyG1Prjna5T+F
7swYpylI9/I57Fgnu8TCY2F6lPUxfv5GykqJ537Bqh8VvRGdO2FODz9fkrZ/V0Td
WJt/Y05Tqgwh3wZpm0bNiqmvdtbQMxGHch3XkGJbpuxO+cLepLj7z86/A+mUemIU
Q+0t9AToWnI0Xls7aJpaKzhwIdXYhkXgO0VSn8yqLCRJelDUyoIkz/SXzmbjq/E5
z6jlPUUsV4bvpl9Ns05mAmOtjBexrFJML2uQVxYO6u+0IAyhWGQpz+TUhsmg1H55
YUyAzrrrsuCtRs25kMi51z6TMoxMNC2hstqZLOobCIHMu7X4M8Wndw8ndjOWMs5q
zmBk66IqpXbro6YPNBpcYZji2NZItWyCGdlb3G5LW6lKY9ZrzGLKXQtVRmao+jfN
WuRgGH5Yyi4zamE37m4ALWM17f3XslDqIO6P3cjSKmRpwfEI2DyqOo4BhUfQPJCY
DILyLrmo5ls9r1gfwYHnUok1esBiyHf8PR+R/7FZpaxEGcXaVYBKeroUImqW0W+D
KbzSfelkVcrMrup3nXvtif0Qgq4pjpRTALKFbCK5xoHGH2cLxPEMkI6231zA9wK7
mRMqULF610a9IEWHyrmeCYIdE8SxwH8ZW24+v+SoXRtjgB8AgOhYiFZCYV8P2OpJ
6oElfo0ijDpRWoUPRu/A1u//RsNE7wnWG4JDAncrp0jmz3kmsaKpxajeqFJKH7tz
X9gjw7ats5Se3JCIVo2PdgVjiUokl1BROSm83+9KrJPRRSANIvaQxOpADdVLamgf
HGg1zNbHDFFjKnmhJJ7xPP38RkljH5bG3AlSCet3tIkpekh9A8MhmJpET3esVpMy
bOz2qDa06L42ekgZppWTk61A2riqRoEi8U3i9BvyXTLmXNdD8ec1OBjYCyFm3xX0
xPlgeOkiLH9/20Wd/EcDCst/0M1kT251/C2/+1iMhf1mCBH9TxoOKbCC56rvwJMK
9Gl62tGnfbY5gL6JKak81h+qfPGC47U1Dw2N3Ujg/KqeQ45djKfy/DUx6KN9rgsu
essrGzpNxirYaE3kEWU24vbD2ANUJvKLVCAFg6Az+f1KrDJ/V319Wyv7MziW/sHv
AwXH4yu6SS8j6I+RiEv4N6aVByhJmv46Ha33uhJNqgkFmtgZqojdXn1eOc/ZkP15
FiNc0xjdZIPahRRb+2+3lkZYwrWYo/d3UyxvOEKp6YtyhULBoCsi1jC9I7t6m7o1
QkpafK8L1FFHnatPPKuDY3D8Svowxr8a7IDL3H4+JtNUlpHXcJPMnUQqhX5awF/m
VPV+U26Cc8oP1cwqf/Ma4K3uL/m2CXmtUpzlcd8whNqqeaChqG+B8xHsR4ISZCmN
m+3+0Sdl+tc+ufxUTMKrZg1xRzY/hqKrz1PDMufSfyYZuYwtr+vgS3C7oDzov0TZ
lzeIEjRAhCuK6dhuIMSv65kbzTtwUfaljLD+JWn3cLScsaSsEdji2z/Q3SMiYe0V
gCassN6Fg70PDKakirbKgLTT08FWkIMu3zIiJN+qJ9V0gIdWczXLwGHSuN4+50Kb
eQnu2AyGcyGKf2sRRs1oSUgDsLjSVoRGjZkNxvqeGLI2D7/O+gOqT1qODWCfeS/y
PeFjVn6qfqS4YA8bOCo6liC6UohXWvwRZm1nkTcNft+7nmWaSowOrvjYEtJpNzCA
t+VB6Kd+oXdGfNXUR6OpZ41Fc2d7kQToKsym6/cC9b5+iblix6cuGUlnXnJRHfDo
YRShxVPfVG/yyu9o8mRyUnj4iF1HXOYpP+b7OhA8v0v/sFIwrZzfgcTnjMM/1hqP
+iCyCROWJTBoZYN8Rvw43LeBFUf76jTRoXCtPUdsrL5AWI2NChrViYOyE1m1vkAd
s3bmz/TZgBx6YBmZwohG3BnloU5Ad3tnZwk1jI81vIndpL7i8Mu/2i+t/DahGF2w
feLhBvttQhKEcra/l1EMNkrnD66Vykl0iJk5dj4xyPZ2kM1yKlE5hhwOSX+ASGPI
t/AOt4xf0OZipQR9pg0B6J5SCQQUtWhA+lSyqZJkagk5GY/OoHRWkZVuoiS7HbUP
cP7aGfiUhNsKrNPOMqYoDqejmWZS+O3sC5RfOrA+dgk9rH8FCbu0kzo3+k+ngEwg
oZGBFAICCTDcOT+34Yyg968CJNcUlHK+8tsV78Lv7vtMiAUbuxWqXvNknwVoV4UG
qh/TiGLVHqR2MCXUk7bkABOac4EeEzZlOxFQdlhyYS5FtVsDcxcdFo/stLKnkRqN
EW8KEN8yM5QDyzn+vlYn4JoVxVvpcV8fKcMhQSQJTpDZ8PGeKUIn7b/Ikz8w0ZAa
NqKjci/MO5g+SySAwApZDtqKwIxMO81L9Hl5cPJwgS2TTCgoH2Hap/P2gSjNHY+h
VQktf3OAvPn09/elBEJCOcCzEnKCTCLkbcTHm/4ufu23JFCoco92CD03k72g4gnS
H20qmukHHayqoWw4qgMf8cQOXIQXUGD2GdRT2SOHyzaT+FUk6CJw4d1Wm/YUYUtB
3bL6YMMBetZdOWjNPfFcX3OYfuyQFliqQ963k+2p70e40wudIwl/6vza7L1RlAzz
RFYV1PlMVlsWrjKrRt9EH86qiWeCXBaPJUmGB1UTAE6IikSUMKJPb62G1ygUWsZL
hfXpS1Fjh4iw8c7xyd3UOtUPNjvBRcsqBrsmks2KeKm7uhBC55HzSP0oM8oaZvsy
+3ylcjS9B+q8M+ihYvOW3zgyUEWK1OVqYMMHW0gcnPcxkb7LrGMy+xFJ4WTuDU2w
0Vsw0a509P3Wq9hMMQA3YdpPYtR6mtVHabWkMaArfXfwyd+jzvQtubQh81yK5G0C
o8JOAvwVKL+VyEvz/NwRmxz9Mb/MHhEiDSpUsuey4Xzb/mAzi2O1MPdKq1XPPRCu
7MQVTLLHRCLiyeVj81BCQ1i1z4kEd1GdE8EHG9fuOdXjRxrAX8u9+zc8jpaEkqGr
75zBh1foQiVCpZ4AOvtPhM2W7tcxkWU8iNRm11Bjalo+aauYsGI77Q7jA1n8fwce
qXs7nVlAHqS+vpO+t6O/Jgo8V+HhabZVI944jPAsZI7e2xtsG6xKyMnYwqb/kaYU
+mwboO6FMKXDvGDWnOKUSkWFyRD6Ne9sXMIoqEN2IadZZHIjvxTOzYdFXSY6Lyvl
1fd/Sq9W50J6LUsLH1HkD7HDyhrIuFa7oZxtCwTDyfGt34rd0RZ8y8IgvTcvvMjL
kCptTB8+4Hc4kKMR3btb8jz5ho7nyJBenLNIZ6eff27UqHWy1HAfmKjR57tzNy/5
FTNR5gUfcyBbn0vk7v0EjbcbEk17WuM7SCeoMzCO4c6uBJSJiM5e6/H8Gst2+NvR
V2cIoL+AeM4M387AgLIGdlJtOgqB9QTjSTWO5KeRb/Nj++XpPZmgBhgtqvtYdqZk
Z44uxICd51mmfIv4Ywn6Xd6kQaLor2VK7p7m2vStKS5kc42vzgc4a5/L1Wy2Ax2I
MtvuPZraXMWvhMewGU7Qqnd38QGowjjzDQE90cMqgypglrJEBLLpWP98mW+eh37M
AAE3XHbPVRKmdWfISkoQh7ypf/IUmGMp3tAGTC6nUz6JB3/Mn4ecPvQmLej9rK1d
0PYFCmR/3ALs6mX21zNZwWqTxfu5k/0ZnIo4N2n48fqQi2VGy17QPaeEgdM6AQd8
65BtihS7k6H+1AG79INSSfRvLs4e3rpEdzep1SuHYkDEcImPKjA+eYwx96aeYFdr
Yv2JsFNPkxI9tuXoUESw4X9BYL+Q0Aj2rolHbCm6ra3ZzXb/CDP47XTVUrnpCqGP
R7InTcdUUhVVqfIU6/9ZMQXhEewu0b9hh8CcHu0d05xIpx+hN737EKeyx11RwAXC
ggQKh0qSbBZ+qMjU6RBMUSjLRbqMc57DYEiIjwg80H0oKyi2O4qjKHD7qfQHuOvQ
pSoCeFiVH+DqP6fjuCX1tNdF1X2ybXDX+PaMDbhXM3BpyoUooj/YNhn9ys4AEqBr
rEldJtEebcuoLJLeVi3Ro5I2xSTfvYiP7vfo6gzIkj0Aug0XCetidU28VOH+hF9W
TFfX/aRZHYmPu0y268vo3sC9n2YvAfrb6XwId0HzpFdE+G3MmvkmeR4p4bCetHcQ
IY25lJmqKaXGIPLrVd+nCnZ3Y6upB+4zyXjLb/cHCq9vajE1MBwKKyOzPox1Dpxw
1ezLtEjyM/9zwhigf/kSJt/bF4kpIJ6oEaF3vjBhDDdc2sCf/isKrBvjSn0/5KNB
gBtKGSkBTB/FItdcPNvQ3g2dk76zoJjn2n23YbbianNi+wmgW0koJcu5QlbNlc+0
Guvd2hZvihaXPsGeBqjrZNoD4Jj7BuFu+nt++YX4uHpdBzc7taI/h1F+Ror78JW6
1O1WrcjaP07n9uJgGDKom1JPLfnUyiu6H6WgyA03PitNBM2V+L6pxbdMUO3shYOF
vlGQYKA5n7hK/oCocJ/kjB+Uy62aUHUKeoF8Qpnb2ZJJ52sIktElrHYhAy3xBF3E
ocz3vx4oAf+kuVrgsGfXu/U1aMUkHOKXsRUHeSs3zk/YQpzQCsLWg9V4XUkurvjD
hqMTjHiZx5NwrTLGIioAYETIqxoywtGi4Bcr8nirdhd9DIDjJxGvB8tBB/E3jlwM
UhC+sGVx9Aa3wxOpNeaGG+Z0QLdYF5gMNa99Svlff7NErivNKdh9l6rGHeHj5jTj
aWE1z3cGvjTReuEXgE5ap1WPRMzragewi9gJMaAGPoDuO/NmwSYVrLiQw9xBOSBc
WZ+DpSjJZExsBZ2gnIDN163OppbVA8skBznL7Ok2Dbqig3B2pyDzQPxJdj4v61zW
Ykv8SmimO9HIm3wfnKQUSnhYtPUSrhKlV/ETkdVfUSlL42tn7QHdbBzfXJenKzAw
xhSgqT2TrKyNuBUd7Qa5TSbZZSc6Hp+1FDJMdRFpisE2y7B4unVP4FIcgXNrnffG
c16J4HVWR4ap/GXe4yk5ZTB1p/vvGH8QwDJ5eMAKlSd4uCsDkUDLXK0CfcbnyQNc
MGIOQBD2AWh8v1KYa0Mz5C4JtVqii73jXHx+ip9XumoN9HnByT6Ok1XDpjvQzsM0
EQXgkzB9Uryfhxb/5fH0X6vwsN2EVC19KJZ19ScmpSusGErnjrXeY0TLvKmeIb3X
v6WnB7bIjr1opskSrpPkezavC28ePDCrNGD1s4KqPeQU93F6IuRGznunMaptB6jS
jxQymYRzCmqYsSnp5r5eGfC0yvIXrePC/iJRU2fbYYGl9vYjn17va+Nau665b2tD
KPLGY0ULYB2R6pRQ92Nf6hEs+axE4yO1ezYDKzFfJMT75JOwcapGh2LFEWaPOL3N
yTSaGZdC/MKHjdBredZOqbLTiAZX7A5xjdt6fIuEq//xNcM04yNjIhh9TCDbm8z1
ODXvkpbDWjr6aNauyy0SLC11OwJ8qPxFBxDHPDaGsCZMHlHPmLw69OwXmbbwh3Fn
/OhgVk8/8n/q5jyLkRqlgHOn5XiPAmG86pOrQMqFKNjFfj7WDyGuiJPdqMjBKnG/
vcnX5p+1jzUe0rH++cKnwsnxeI3DjZ/kTr6al3d9OfeJDdERSSVNcH/QHZ6GL0GJ
Fbad+ZYi79j0DPv9xBuznAGvi1j3ZIxBivoGTMd1jtwAkQTqTB3HDoTSusZOUt8c
KYuTxUlwGWf+mcjZl/MPOVuUcnSmOHqD2GI+krL45rrKALkNoxFIR75uhZ2mQ2xK
8qDrhKbuJtH/ilRkVSzDYS/cXU8pgRo9LTc8igEU0c1F591aBOSiVQ9jXmUofb0C
3faMZTJZto2Vwytv+OwtNmfVcToII8sTAWenSspFLYFcnEiciRyRvZuD+WX4afXH
kM+b8VNM7ZJpFu5b3+XiUr5VapX0uViTJaJ2zgTB3lofAdFpHGajMa8NgVohvPKt
HJsf3ABCThxd11UAcofUPEXdvZM+q06B/N8HKeA7662m2fI66tullaXcrRyTCN+f
5Q58/FaIslb4nBrJTkV37Fa4hBy2xxZHEfOf+J9cL9tmwTo7qXiUelGrO3u49HE2
J9PqCLOh3QbOfC2GEMMvr6t11bQDKb5Flhl1OVArXZ1Xg1V2j0Z43CrGqiIBm3cI
S7ZfnAQyel8O1Hrd3VFlNOG9tzoi6UjXA0KPqDwE8ODRILcvIoKLq2pDtA2CEnO1
xikAcnSQXwVGHDdRbX40kXxrIx0jUYyHG/jECg/0QDBhIKGVO9hpJeJ7PfPYx67r
c6w+YZ5wvBumT7ca69gN6ixqTOCbg94cYXVxJ+pfGUBgMvYMlmvBFmvdlDzrQWzr
5BMsXO7vf8PST1XWDG+OGT5ZlNVT46IttndZQ+O4oKqO3mXlufXK0fXls1bsmD/7
RCAF/d1Tn6/lDtpw8WWaye5LpPEwrTW9M4B2731CeMskJyn+o9nTGsDBhRisk9oq
kLVOjYmL/fQzOyoWrRRRM6zuDIMwhsa2pjlAgTmFsbuKD4NWP0egXujRv+vAug0C
2K0gdNl1o1ZOz9Z4Ac86sS5Ol9l2yRbMUOUAwxKb6i+7xata+/VFmxqF5jDBiUE7
9QKrW1QdxW+yBvqktAztdekB4Qs1ZBDa0xpZsm4jDNX3RJPaq22lWMNKvS42M5Lc
mHpJlswxJ2aV6qdbRYu3EVq0ZALr4b1YI7tbQgURt1X+IzRU5cWJa5hOh5bbeLmv
JCtIazjbAxXcuewbsDKkT3GSGRAQJXpRGcoyIxgbFn1F+kI4AgQq55lvmx4MzHrg
g3W41WmtjvrXS1vq2Zrt7z+AEsSeBr01IEapPdOfbBXWchmpC2WAbOMC9TQqhnTM
G/t62rc2Ewd0wPL3yKh/GT/s+fOCs8rjNzuPbjMMlDkIMyusWtcLGomU5fqDgSWu
zwNOR2nzR5dwzGpwWADJ7nYBMm2TCKNMxHPweNsKQ7Mkp7Z3lpMutXgkULCqccFX
ORLHNi4jVrCEjychthTh1Tm3Id3QF09VfgZUV3RQNH94NibmnBMFZxI7moaGqqE5
1FOUpQ6LS3s/97IHr70mppqjfkTocBUnaYcU1An52XVA1bhX9Wsc9yQQGxNVCKOv
SzTjlNl2dvkZM3pTYXgqJKaST3VDKlY1bqX3ivDJ/3VQfHP+5/Hv/Aco5rlcirp+
3PWLz4GOn96BvQvfhjs7ZKaNsqlfFJlvoMPDFcDSMW/omVW7ZybfvYxUzwrn1n2B
lnUSOoRyCLkizS7oHv96JzqKZFZ8iv2z2C1azvQBhMzCxax7tLvV41sFgz8D5K5w
jIU0cxWkyykCwKf4JVzbjfmSxArwWBy6WSEruY0VVu4t0lT/xATnx3rDJvSjcM8e
GyYTRHX04s9pFYIV6Ih6Ny527h136SBaWDj3o38xuhQvn7vrQHKwQsOaWq7D+g2i
LDkGAcSgNIuxnTZHyNGKjHPOoo5Sj+4TyakniOyRD5sNmO6OiNwxs6pJOiEJwSLP
5Zo1G1L3wuv+CN9z9Z1Ut77yGacT6IW1m1+QkXJoD8T886Zb7CeOU9olH9lMdf4T
IJNZ4RMQbFapSJKeQssxggDnHMEbRTDXYznMZXZD2VDaLoDR2t0eGPaboIk4oKLW
OwkzrOygD2+/gjT9RuYvgzcrod36FH9rxLfGLn8IqfAFVoBMmcTybbHWKNDH/aCt
NGvx/GdZAnJNsfmds4NoeLEW3SCzkePvw0HN7M2Xrmy4xbYrGcmEG5MLBE02MyOh
3ujqOLEPenJIWyL9TVqP7wtWLAnnefyswiEvQQQbqmoJXMddUUH3zHjt7SLXU/yc
jjlZnGU+iza6NCy1sgPymh2YPbDKeoQ/nwcWFcUgIEy9sMadnCbCHe8MRJs5Vjum
uwCK4nufVpFHcXdJdyqH9wqjC3+cgcujCxDkbGDwTjDs2xljYE2udzTIZdr+xYQQ
0lGyb1Ops+5fkBg98mbQaMQ23YUFlRpPSjbknMa9/5huKJRY5erU5KyRlGU4ck5/
fcK3L/Bgj/IjS7Vj0823ZO3RNEGal+V83EqfO440/vsFk++rJmxEdPZk3S68qPAU
Dz34lj0YBfxRypEjFPEnEDJlAErJaEklpNBUg2JM6Kq/U7SY3zfi5chLmlg3mQ+4
TsLBa6QV/WFomuR0116sgrj9+xbmYMpFmPZhr3TyUWH1WhUt33oBYag5YOw0WdkB
L01Z/iqX4I2jhcCfbI8W/eSKeHNvv6xxqvVIFwbSnerGrK4hGpWgtGDvsyTJk448
NmZegyF8LxMwgpXqd9tv+wpDuY3H1seSeAK2QEtJC7sPDOgxAhDPJsjD4ZAILcoe
YmfEIjWQAAqmM9UC8DrGV6cbPQIjWvPM3uI/HtbLCQyHqqAetN7pinJs+rjSEkhv
5EQqsVliACU3wxxqswG6gB1j8Q/rHLHTmdILNNmncqz5Bp2tMjUVGm3VxMTllMii
N/KDJfYMTdIfc3EMM8u8mDmghqoQMJGAXCoOm4vylhmuTifcA5cykfvtpylcNYDH
nHvH8tBrChdXJX40Z7x5gFlZw3vnnhISVrfXKjA6tnLNqMe0EybBIjL09DV+V8R2
qMnYgevejgpRfwioUR/LUZPWmhX0qAjl1g/RiL5xkhtsh1rwGH+DTvV3pktm2d9i
puMAdYmvNBiUwET6kkULru3HZu5shSjgnBPI5+3x5z059EGNrxLjXzJC3srlhRLz
Mu1fWVQ0MsOKypnQIVf1bfok5HftlDWRzQR1u07oB1WEr8vrF2yJmPRlETlbn9zA
Bbo1P8vOwNDfbB0mH2vbWI+ZwZ8Qks/gaipOt+iw1J2U4YmKBz0qUzaoTLEhzolw
pBTUSjrMkwPDWhJ4k4Yut4B/sE8EJNWOKFql3Q49GErwmmjvEiYX6tmEWaycT5QI
/Yli7kPdiSNGkK63MQsf6sAAYfnUElVA0hsVdAuNc24ym4lQ93EVlOd61KG5G4c+
dc9eTIu8sauVTV8Zkg+9mLbDJYDWwAfb1DAimaw+MvrN6POU59bBGJIFzea+L6UC
Lj5tmwW4jXU0e5NxIq77nTALS82WIARXTdA3t4FeOnnxAxet1K/xOudOPBbBTb/j
U5T6nrulQYV/afUfEXSYshXnZO1kw8HntGWQort/Yr5nbx9F/2E19Lehvmn0S+Z9
c1pjyDvpiVLYHNM5Eoe6sUbG9KQfDGMOcBB2hon6ikKBiJ81R7KJhA8MhE9YN/8d
ioYSjga7x9dTP4jG87s/OcCYpGxmoRvnu4gjSIQL0RpcjpqUHZYoESRokbpiw+94
p2jzuCrUMJy3SPKPZzZP/z+iFC/fSDDC4YqOrDZ5uyPBPsUPiYZKaOjNf2f3WkVI
pF87cOCENi98OAIY8E0KTNgJByhhpiS0h6Oq0cIvchKiZp1PRYXiFN4UjO3/QCF6
oBzzo+yo6iJeYOIGeKFJLHQRQuATGfa5ZSBxwBmMn4VSsWimS+XSoPFksAnbNcxk
RarOv690tPAD2x/Gz8OFvX1LmC607+LmluxIxPAOSYHi/fgMTbNLvvRA6Hbpyh0l
mHmJvuXKChwQquIvTssRZa0cG0TaWwf7lYylqo6Mn+ZouQXkb6F6GaqGrQf2XFRb
7frPLpsNsOC0Pbe/eRLb99Eb9SiXM0teb7iy7E69eS3y5zSUzXOOqNP4WyeoX3FO
tfRYcMZTRwArDVldyML11FEngTmBOIpCaan2z6Bsh2rL+EMVlqlLr5kfTanvybzh
C0KWU+glvlWcHDF3eJ7NZcwWxlm1r04MzjyRt+ZaRnX721k3WpFnypWwE0+gXewK
eMwtp4S4QoWRg1kBgWO2CAghTgjYrBlqTlzVbIn5XtdTKOI2NE+a54XItlhsUqSQ
9NziqkvMMcnQXPbe8EZZzYXe0r3w479TDU97tFKOAnVemtVe6W+uXNfXTYeAuitp
W28jXw6V33an/c/Ny5ABNlMmNLy0bFBTXoe0PHhQh+SyCfe4c7vAqCLPS2rw4dm4
UMwuSOaEr7F62O6upesLr4PKCvt2b+yscLquz3kBwVtCsmiRP1A4XjaUqc6bN+06
TFCnDgbg+QcteoyLJw25saFtVKlqKIISMoaXVHlnKFAOlQkrohmnfB9NRPf7bxPZ
6aH7Wb67KEGp46RhKRfE2PQj4+F1NHV1Kbo7tGFBC14ws7zF4/aFJN36DQcPDywr
tM1J9lcRzVIPO0FRWEkUjaoM+IxDl9ekwp+Snw49pUhrLZZSzfCyPh4lSIGEfhlg
rTSgh+6GvQAf/zHQbGbxmxdduHxDaILy7eNgB/MhgRBboCZXl/hA7xBfu3PZoMR0
vOmFelxJrroqISZ34//Oa9eLBILR9jejmr6kssU4dmqs+YhJgUcNguHMrJf1LRqq
NDfw/gkE2HyFBG+PT18Rj0/Kq87WiTGE0ATOZqaA6vNX9neZ65fxkqQPFz7ZybgS
tA+prcmRH8phXNgrPq3nhlykj5t0oPlQugpm8xU1Jj/CnseQNUq1bYsqYpmDm1gp
jc3AZ4sMqLgbKw2gjkmkPp5jn9CAl0mpkCTKZBp5K6PNG1TwrLJkquPYoLSSnCSN
UztYMIE003Dvhux6/ZcDFDPb8BUUWCFAHK4//gApZOeFmd1SZIpjInSitkwG2c1N
Kdi2YITtXqwYYqnGB+jNWWB9KHwelRhO/7skdgRq2baoqsotg3PLi3E9xVd7laTB
bb/toqsNnDCo7sjKi/Mv+hWq6e8bGOkLp3FxfdZh0A9yKXFNsjJUj+RWhm/TgziE
1mIBf34uNMZQjAcbt2pWAikDL0Iy8egU2ny9F7kj9bI7ZXXbVxeDuqaaoQX0CQNW
ooLeQZxhsXsbeVMfEeIMmOgVkqlzu/WQXk7dIEv6IujEWzyWhhdI8ZgIkGMjp3DQ
ctFY3HNeN0vPUWrjdeVcvLVaRUusrVr8Xe4aPv4yQzPgqaSTqQRTrYgVSIKYyP4S
BWn7CyG5FHAv4XyWjw+v532RSAGZt0SNg95XJJ5Ingv40ubyuxIEHkR9/Biyk12e
cQ7s1/1BGzxriRhTdVZogePOskgdQ9tLUwQ3T1LpFQRqvF6wa2AanudmxcRrgmit
2f8v1ZIqf7zgvX1kHa7yM3y+/cSwE0wpLN13Eihpj2tm9TCg4LctdwmR6CwKRUWH
AG3WRwKLX5ep3oOuqfitM2OPKgXQzYcg5lWeXW207VhMeBwZ11uF7fSqMKrUcgWm
8TQbz19GWX2ZeyqA9x3VW60uridqmvw7AmL/4MTB4CTPUjMQvbp+zCD/K3yzh6zA
GkcbxPTEnZqH5jTtba1ldws94j0vYVo9W3AWT60v/+xgOO+pmaFOFDi/8dMB51C8
G1wfYrrvggw/wbO4ebGslppXqC+ueRdtgWNvp22E6rT9TF3hqPm76U46b5OQCDJm
GE++3a6UBMdG8rQlOoDC0HqhCCcc6v0vgEovOz7eNv78WJOjUdNdoAkQM+h2LSI2
8po8QK6W43LYz7WhOzc15KOTMlcyfVJ+jiH6i6QGADvVy5tdJUMAerkEaRwyhpcF
AJlav2p3tk0ue9zwhlyOftTFt3xoYgTsxlY4i2x+xUq8b0OfKi/3C1jn28hbzYly
jCDexEyRzsPVk4z02vMwkpS17G+xGR4OmtnfroL9SVc0aFFuuH5HNcCWdOvzYa0K
BhX1jl7x6ChNYT+dcxrGqGjK48AwRIPASU1pmClmlqRY6mmBuo7j7dWXDIUuyPwn
q0ZdBAPl0uAy43sYNMnhY7iefLatBgQW8pOq7ZRpPdeBhYSJMBq/FQ121M2hXOMX
FOt0BmFIQTvvCBghIBWLF9Go5DHUcoLyWM9IMrt0tAJXPGdqteFQqtxMdJx28Ahc
nPz5APk64CLurF3i8LiRZkwFLBT6cA9Nw1bCSan8OydKU0BrWNhUuEDvbO5maOtb
uo2pcaXkNye3nfOG+Wnf6P5Ujql8tqbA45B6VP76MjazOl2aN50XwoYN5zWVMW3u
QuJsYQORLi/4ZtyxBUSvjUxRxRqsaAC7QyemYPgoO0Mugy+xl3AM2882wKiamJQk
aB7Ndg3PP6vCladcnYVAmvSl53a8a3kHGwSfujTmLCTvoeK4ERPdNVQqdUs1qj74
KBOMzxphx60nC1stzdg/iasvEL9ZK3RHLVb7FCJ2Qinf3GNOjyNrCfi5fH4qSdjT
Lo8Mq+51LhEOOz1ZXvQpID8F0JySxHdQtXi/DaPrJO9fa6e39ObO/qbuo0Ua587W
AXVM7Y8ajazpDhBk3SwxQMQ20P3n0eQ/uQTvUYwgjhjlPkdhVbg4Toml94/SQDFj
KI6iTeWt6svW1EXAVE+YxyfExMa2d5J5OPDzM/n662NKaVNeqDAfRmEvXLBv4bH9
zT6MkhVDMBUKHMWbCWGVbQQV/er526JrlhIjPb7ZnXpzvOXJ7OBvNUIUdMu8kAmp
DjxBvdRTYXM43BO+yQ3jNip5imKue1NhbANO8dhV2ToAg0BFTR3FBJmXf4glvk7f
nRTjAqTWcZO7g6xzeWDBdlbj0ORogDQ3dyE9xedBkPkYByvZrrzy1bPY4798o2qf
XctpMSrU5cDVwoXLdGPtlP0MKODfXOyhULEMK/glwLkmscd34PSVnlZ9jMuaMV+1
gaKYQMiK/tOpF7ghgxqDX9Af5HSoT+r2KhrumcgX0vubABFiNoxIj1m4N8soOArX
2ZV3o7Hvf039UiwlV3UiaNOFJby6XdSkMswQC0Mw7vyTKhEhSYRkMVckAxlIhNZE
mCx21pDNPgO3SSK/TkbyyCiP8muqWFSdz4n02S17oKiZAe+bpx0bePgtY4Xmd050
Q8d4ceN+ID3Xw9zW+1kELqpDCYLmzlCTlm8ygnpmrd1UmDoktxan2QHm09zq/r5T
bi4VVSPNi6ZThiz23fO3TqhpHxMqYOzweZhZyse6LZbF6yp0P23WiTaNJjiGWHxX
b7ZYI7Rdh0g2WNr25qG50OT1iPICEpG+Vz+q5fcN4+P8yRK5WFGR6Gx8aXxjwfmy
z4x36kA3AIhKLsBFLSwRURNwOofa6XG9GMyPhZ5pvqGstJWKzStkEhojhYvwfjp7
PA1dziN9baQGfVp/PfhcRPz0H9cN9GKXU95x+qHR94c3Mho1v3S1OGIHNhnUYkWH
tzwD+HBcXa2fQ2r0rco2fDx7fP38MSEltoZhxa3G7pncaAzOoNHCfcbkZcMny1Qu
WDkXJGs1hfLIzZJ18kbfaSx6vPQOrWlZbkIhsWGHtfB5v51LRHYKnXb++V4n+Q4z
+S5bOWRa0zGKl2XCLNXqGHCh8KccvqIHU6XM0NqvwLJ4uf+qPTv60emgTV3v3Dou
5dwD746u3NU9fKT+qAzzsziWolaBjPGknKkFl0i0L/cF0kXEwUnvfuJnwICtqr6w
Zjf63EFPZM7607LqsCeZ4ecaZi1sGLqNPih1/ynjezFX8M9gpL03dnAdb21IautV
i2ObxhS1eEu1bqJcSH84IEqwyJtQqHpX7+eDCPeOSORXbNP2VKVAaksli6UWsHUd
P8V3QE0WlNco2IIMm9IwnH7Ti1fuAyAcZs2Da4K37CQWGjGjjAmBv6iiWMLbJq9e
QfW9GdNPW/58K/21dpEZhPRVDYMNqZeAmskx06DYkSkuhky9EwjXXVQsH2F0e+tN
lvleu66EAm/jnW7WL6PcBWqNVUtS1jsz6btbQATbUxL2GynJHU/ID6CAqTk5Cc6F
qdj97jjK2v9LsJCK7+SZIUedS6xZVdSHAm3aVlplOAJKVFXJQ8dlCqTzpoVV8sSK
q1ciTi3CLY3Tv7dgWuAM6TQb3HLoHh564GtejPcBA5ZTVpwdhahxX8RwLi11XGo0
dpIY9BEJ340HTMHSbuMKQi+cXmR63UVloxvE8Ig0OapJUXEMgk1VuuZcG7tkUBO6
kaIVIjwcqMuRLBVShkuCqltwqfTGlOdQk1SaZ8pFactriBtTBGjtnpD1hhSO4QNO
kFkYY3GGkX/kuTNhTuR0kj+uFuj0jBSK8VclNjYoeW3oOzjSZg7ezCN1TVxDN/yx
gV+tbEsCJhFW6B6P67kW9+y7bUFuyotcMvxG/PgAL3MRFHtONhm5Zu6hvyP49ilE
trjjw2RZ0cY7l2i4crjBI7Cti8d5qRbeDHrrJtQ+OB5Z7EX2qT6GFsq6ouQobCZ6
E1XSxhmtih2Gf4LywdpwQKnFPthzw0sm8wtxjzlXYvpZcpLB14WngH7M4CXPn6RF
wFje9mOuAxWHsSQ3/uOCj5zYvAyD3lQ9NHMjgavIviYjJLr7GB1stNoMqyfNqVQF
C1VBnSDaydCOB6wcbIlulQqljBxMC8efWzSURGyC7R95rBhlTw7BODEQad6hJ04V
RSfU3xbow0uti/N5x4d7BIGs7+kHaEV0YAmp/9xX0aJUOwjb5IwXwnmAZYnWNc0w
kH3J3nQqUZ3k3BZLbJsZAWZmNpUkSZonVKNILMZDEvKUSVIcGe8Ph7Zk8iw9vs82
sr53/nJFQbt4qoxY7PGqt+5ceH19I2/wEBHyb5eEb/fD1DRNIMmbmD8yJzwkkvIZ
LWyuNUUSoijtonjChcoC2qNvLl33PRn3+MfIPEITS9UOmUFvBGfLPYqjy6zqWu+H
CHdlbZhP0YmoV0NHwRKUUIlAxOL19aYIfsJzWIBC+BWrSDdqrU2ckQ1Vwes7EfXa
vhM9J8J2ZDjw8tB+/cf5mex9lZGDvGn/wBTQ9uTKwujh3WgunJNWhxScYC9OaIjq
fvceGHg6CgwHe0BY7sSk7Kfr5hYO5ZXcQMn3/VC2BsJzOnpa6r/DgHeUzcnxglgw
fPrGIlZ4KmVethnugRlQc6ejUcUTsFmn6uVl4hqeCf31sXkpLPaKgd2BBi65tZ1L
KxXHVpQaYEdi6vZpyyrLCAfgkVdCz8AjdLjrpk2sqfNa/UU3+tJVRatVM1WyM25y
o4SljZrEX7252lWLdLjX6k71aPN2j1joFOf4AzvYzM1uvT8j2DKPeWUGbDUxDM3U
ody81t/CvwqA06nXaRtA3JS0h3I+GXrwwsHCt04rufQmobVsnwinPlHQY1RGEqc2
96mpewTQVXAflyjcDkPLR1NY2RJjS56LOEiCox4SBiCitIlmAD+HOxcPaPaoiDYW
+3onJk1fxnGOwG3sN3cF0i8GEBJCdXH5WVvuRzWyd0D77iyUtJf8Cap7JM//6Ed4
oDU1esCnen8rNSNHymPY5kUPBuEOMCvj86NPLE8cV0tDGW0sYdLftGXXTne23a8s
5LjNQRAGNNLidUYdWycGP6Tmqp5Kti9ptU1QYXJVZ+yJFQlDz8zeVeVc9F2J6a5/
Z2L7bfcvnbqmKQC1GlfY/dGnKKQusA2Ra0MPsJCp4OppgiIfn3kwBM0AJ17aAFM2
Gy6E1r+saAfNL1Ite5lrMtwOFVOPrFxoEt0Q4m+goJuU/zOzG0Un2sbLEVHYZoY2
p89OIeLjdt0LxS+95c7Vo6uqWSmGh5anZOq7Pbny6yfHb7PrimC4/zovJ1QT0g8T
yW8BymCJxMlXYMZnyvhE0hcQllTHIa6dpvgULJlIEi3/FPrAxpZvTs8zqbzcvzB6
6I9MGTITeWsxzFej50vJOqUQhvQBi4bBWPbwzKuSI6ondt9/XeFvS1mZorNy9/ks
dT1LZV1ymG5+cSWeS38SzR2yKsIpIFmOtAAbASMxzRQ2Pq6V2AFhXF4lR6SC0PkK
c8FcBwuLr4jLxh82/sIwZqPOYB/UZOgpw0ojGYmNqijElV+DWwdNbYTBCAmV7hIX
O71bk4ft1DWJMERvqvwASsge3oRCWdj0EgIN2Z4LzseakfuIcVQMXdGJ+L9DC4JI
Vn6yyUNyFejRJiZdbM+OojH4hTPeDvVrcQW1Nj3N0O33/9YNFnACZD7AACV/HfXH
qgfFqYoe7j0x8OtliuLt4IqSySmF70/pHyEKbipxSVjvMmqF7v32PZVG7GttHMY4
aPhBwaoOr+gKB4jdepd2z12lVV8ZjczbGBzmZKENvfhorlwaTgdMtxYruxoq6uje
SCs12xBredzUG4QdklaSzITbYub0W7IPLY0exS1WNHZOvjs3KIeaUR3Eo+HsgWR+
0YyTVYRbEL6/4SQ5R+iH7aLIOebzeWpr182/2wmUuUJTc/k+1lhA6V3BetdEBey7
Qpoj9tzCynapap38HAU6CcItjz+EBuPoLCtoVKIFlrcRnbK32i3wRvjel/m/bbK1
IfuuVPPdgjfkGZMxkQ/BBFueFDSazGaklzXaaS++l2Y60+dHlqNBMCuUR1Qk8qCK
CJ+WzQrGT5uBGNXmvEvf5Fb3/XFPnzaAFyc+YNW4dAyP36UnVqYwiW5ipZ/2Frgg
NeyRHJkdGPAv6rZdSW9z1jYMQJjnuDyOM6KfCaHbFBY13kd9tpc6nFL/LrESSJc2
n5nP098aREahzMY6ZxBWxfPdfZ1WisX3KBiSJLKvwHTcexXd/Th4Iph/niZ4Xlae
Gvo2vXtOXUrHAOV/XzxcBx6Z3FuGzfgujbpnlLJq+NCJ5oDBqepnSj3EvUjQ+oAG
Wz2SyGg0gjTRJ35PKfOwDyWt87WrN6glRTx6J8ZLFyJKL1phCFt1E2YUb9iLIGjN
bdqw/Bx90U40t8zi/zAnczf+C22gqbB0yvZQj0wB94LnaE4GhYB1buVdxYDuZjPy
skpLJQ3XaKSNoii41c9cUALntEGm9wLKadDrceZNqrkMOTBIHPMQxtblGUD77NMr
GHvV7Lz5M+8gBvcaES2bCQ/e5YDGd2yIavc6w15t7DyZtcUzvHHZSDQiecdJFjVU
oauxCgLdRxzwcncDk9ua9iPz9IQKS2fPJI5NTT22VV+YZHTSh/Ugl4vSZ+f4Ke84
f03T7vWUri6S5im9T5RGVEhiiTiNB0EZ5sZBxI6L3wtjL+81gNkBlD6IZqLl+cEy
IYemJADfBZKYqoDP7UmgfsVDJn94E0OI/qBqZ7Z4dzuTCAaGqfj9wnByAYWm7qIe
nX2pGvXtUOavuf7j1ok5dUHqCl8HXYwMh7GDxof9gzsVGjHVD48eEqQL1n4oBxSr
2ej9BV8Ql7a6Z7CJHrn+myLcGyes9lR/itKOq5eDQrAI48/g2dHNW/BVyQlfAsxa
+36IpwoGscawL8cxeuYKN5zjH+BsceWMiPH9ZbK0tRhU33JJh1gRSpgNb8pPjBrl
7YRTalnfiVRmWs0vOHkKaz9Y2HrzUir/b353MvmrYeAoYZRlASnmuSglpAU4lH2N
IXWVBoEfEo0zyQTdAn6sFTtNPqDvVm7oGTp1PyS4fxQBPlQJZqMfgdWuSzppML1C
SR3ghAY0cY8n5X7k7jEdNbQ2CxPhtRFEJ9JivEnY9xmCoFKAK4SncxHjznXb2043
aGzpWTizwXJIwt3Gs0Qze9rQWfIJ1w1d9v9QusUZb8upDnDkDBKfP/eM2QcwZNiz
g9R/PnmLAcK5w2Y6mzLeYMzKaK5oZRKT+xeyvffsipDQOFQ6oa9b+0Ronvztz3cN
53hY6HihPB0yrVtMqfpFti7mjrRdFCOIec4Vlz8KynZ2jzYj8JL59sI6JAu+jU/6
pc/SSQTHhGOiHf4t1O2menF2/Evq4QaaHWxYu6NhZsOEKTm4dB1pz1TvwlGtlu67
3uTmpVZqsgc+iIyBN7qOU/RwsTi4mpr5qlE0YnxTaKBTlotZKo4Y5JzQXYEXaXnQ
nsqaQqCVRxN+6e+rSK/Gjtg92Z5eNOmdbCMZ+nHMo26aBp+BiWwmCKpScbRUzDNs
Q2+1o34HwjoNGJr6+RF9FHJXvKYOzlqd25NVGKPdgRDvADb6MspcLKmhIcm5PVCn
1CuI/VTlpr72Mqvdi6C5hXuijHIOJud1vWkVdV43qcMyKw7nYBsrG+zMuH86XpW6
SPI0XzeAxwDf+nBJ0ULUj3+yDtpns5g1VAze5b2xBfZzT3k+64rCxltC3nbudbb2
GYLnBDXU7Zar5ajLv+woY1RMohhsXtM/hn2b7OakhM+lWjDqOd2WQlTPl3NqfgyP
sDdWd9DnA0i5ycGQn+pdKQaRWItKMO5XSZZHjJ/HjB/p55/Ma59oYJL4Jzr7RDm1
fHN7rznN4T3EGu85YDDTdKJSylnZOBWQYo8oR3FVGH/1PZJE9kwptsEJfInkY27o
z3G1no1jtXzKhUdTIRCJH7zUV1A4YevJzuIKCDThFzZn2eAPJYswlSzKeWaq33Z8
XX2R581AO1WIdtmnMq4X897eWMTDKqBsfIqC47pbTyHR5GZhhkBFM6H9unl/8/25
sKAI/bE4fR2z7RVjgSWR2IBvnAIpKGcc58u9U6QljUEZf+pwUzAh1kx6lH+YltSI
eRHLx2i70BvISmEe+blQM3hrxyfk2yBI/QU5Iy6v67DPCIdh0VCk/qdmoOHC+Ulb
6jw+iETOoEk6UHT4GQ0sUd3rNw9cLTEqRnPSjfzGrzIdik9Mj3lPdc0LSDJr2bIv
Wpw9AKaVuOb2bCxKp+uWh27SPbddyjfZtbYJOF+lggm87RF09ymXUkEpeYS3o3rA
VPnrEzcKkxRb/Ra8L8SU2+aP2Kb5Gl+4N3GHVXD0YWTSch3z7h8HjIUb289+x+0q
AyoHkshH1yqIN0uG+JFBpwVjsw2eqAk/oO2lfCF1r3R4JlYLEUwIrV8MPG146LPc
vK350VMMlcUd5dFqhgOrrXbBIdb4tjcW2yWjcZsSUiFoFCxK1f1v3VtJ+6bx+bMy
iXW7ydXPawO8dAOW3Pg1ssPJGmKZoNmYf8aSzupOBoF8/e/B+WgOFt25jT9LMzHR
tNhl23nViikLxvTz/ZR+pevLAPk+bgncDvCbwh6YJrM3u4BverSF7fpp6YaEJiAU
gYNRT8lpUqMd4QM5w7MfFshQveFtLi/c0pWGOCjEf2KJUaf23QuYJ6UxcegZmQbT
4fTue1dbDkGbUUqFstKRF4MPGaapZF5XvrX0409gDr3paZZW0GHEGHr1R5uHjjst
IFKPFD0b/toitBrwvuF00HJ7hzOWLtVQi0eg8tS+rCsm0DGXGe6OGl1zlnIhAnDp
ZGv2pCbTEkuADMWuU36boPh7ALU8MinqvjosiMbtF/18VK/Of3Rhg5abBKlsJGPK
G5YttpqGvxNjDgxV+NgtmHGMoCvCoEkKjvCMPSGYQ8Q3e2S+DIpqvonFsp9oVyKZ
6wZqwAg62UFc1FRyVupBN32jbpBLD1RHZAw5va9z8h4dnEP8g9Su2qdTTxmoee1v
HabPgTmwyT7dn1yG6TWnFSK2DzT2/vcGKdzKI/l1BIedRGIyJxFjC9R10WTJpSjr
XROIX1zAP4mDQEfgWtGTexG8N5LIBYzrxTBF1NSFYujTljv9/sPUd6o6qdJgFdaO
s+99fH5jYwzDJNqOcahT4gst6pdgNdHJhStMvITq2rkXYq9JRQs6NKiOTBF2yrma
KIlgukAEB1/rsFhJyZHYJCbwRlh1kzTg3zUvP3B5QSB/ftNuoc7J7NZfdkHRUPrf
bOiKizK5UScOVdzdzKFOMV6qMa/WNa96S8YXINx5bghaN66rxUrEWmx0goAXORlN
1ZooCT9l2+J1EpI0UycYqNu4q4A8YW6LoK8wzFU+JDOUOEmoTXI6mmyO0x67btcM
t1GUwuAd+weoVtSy8p2hQK3YPTxiRE7n4633RbuH6aLqe8CDhIMNQsv/42TSk22w
fPd1rrmYucVe/vkVodQxLXvOU7Jbh8nwgul8t6iTH9leAMjluzNLySmtb4FcxMLP
gEqorRA2uYIR696Jsacp44dTu+ZezzeABW9VYtJfoH1Ivv9PS32FDn9MHujwg4P+
cSf9fT+fif69y8O8jDdnssj/bXJj3XkVGwGtB0RQZqweeLlkv2McIDBXJ0e47lz2
5VXUSLtIm0d0JUTx64SSwUjMw2Yu8DGnJxWfWTMV/QBkEIBHQMqraMkYXnVVNO68
3HYxplQE1gPwp7vbmZ5jloF/ERqbSjkrJM9HEJrLV1FDzBq2HuCO9dognO5EeqHq
Whr2y8HAB8iXVlFy6da6E1xhcRqcjUAqf/vF7l4FkFriCcqVrplCEfRN3G6+OoUI
JU3mYddZ9bsK/7AEQURpohRwDju6askQPrBIycMRP+LlRo7wFV6SWJfc+tGc4puC
v5dqfOWWHp/4MTAGMUEr7Jvuf4geZnZSBn2DrdYXws5JqFB+y/mz2gtmYvywohti
z6gENenY8ymvUJVL9bWDVVMbH5xYCyLvj9fG6xtZPkm0BkP9+jSvuqSo+N/Yr6Wc
DDyGzS5G9hrTnXOKvuRqeZprT6pUx4J/EXI0vrslHrnLFXdQhsxKXKnXSvde7GwI
jNTRbrOkqXvYMoGIBgW+41QRdm0e96iYH8+/MU0aSVxKC+v6VPSZ5DB3U8VsOt3w
XcSAeQIupswm9tZrUQP+k8jpa6lq0SRgnnW/8u1LVkYfJDale3HKstnDjXxTojhu
KwMlsGOr5WACvDqwSqHdZa0Mf84tx/SkrEdbAmfr6VorhO5ASrJ0i1n/3k97RyLg
+DNCmuuHXpzL6CGa/dRNUcTchjPmMILw+ofFrqAo6mCo1mD3xnKtI9wihCk009O2
5aucmCi86jKId+6EoiHAR3mwVyAdrFPXwv5KobCAwpcO6EJEmkeshSF7I2LSuSzo
VWn2ctrDd3cOwRQbQClFRoRjn6xGdD9xfPlmTXMlc1rM77t3vBn4/9WGemHlWT8G
tvIebUPcD+Wdb9WRbZO3jGHCdlAp5n73uohLRyw8Qd3h8BVg7xxHzvYS1iIrPMj1
SEk/M42Y7LBHTObwdE13y52qsYlRaPmDtsfxQNSZxxFeLQ2Giigd7Uhs663NcZnw
MJaYw3FmkjDTFH1foORVbuHkUk/VcKfGKSwt/HRIiklPRtuHqtKjRUasemwl9tx9
PT6ahF4/GwTPkShhjvONXLdys8elw8JwIM4JhnLsevOD3iXJnklv+yJGJmF9CiNI
7e6Twbhklq/iqrwbSRkOSAiSgJTSoCeSVJEk2D35CINOpkp6gifjktxirmENix1V
k4TVvikXiE2OzoYCzm6Ixa8Pge3coIfp9T8eSWpGHFQ5mQn4JwviU3uugXudh3hh
7XF4YCI6eoX0vfd8qOb9EREJEu5uKbQUy/hNjqF4+TPW74NiA/UWZ62Uz4iwIefc
eQsq9dA9sVjQtx04gI9RwZbLrVlqwWt7Sr00QOGAGRG6E09pJOo07gnzTKvzyIWr
eeTbBAkGmsRwYernZyxYHn5iRoielwg5B2VxZd8zr1SYF79mncpbbFeCOwIN0dvS
Ue6tQ28iE6Tv5cez0qIkz/zGS8uF/HdmXJY7PLa7rqPixEQ+MspX9k5nsrPEs4tl
o/SUvMHvIg7lNByYdaEnuq3Qo3metnKST/xjQuIThhSCgN89IRlr5HJUhWJeNQ5n
mZQpyOFrU3JnF7LFWSIU8JwET39cpkvdbg9xlJcPsmVb8NBmilHRZqEwd+J1fq2v
uy21WK0G1/GKndy3dvKH7y8w7qwFf/Y0gPRurWo0p2+WqjlWWcTwk1QOqinDCUx5
bdNMlA0T4TrNLUqcWIDs/EM/4iJi9GaIBeWkto9EcUNiVWhsH2WwpgeCP1c3NJFU
a6FCfYEUR1bl2mEnOW0Lokge5IYNsx+0ScHhLUQGr5UjIikc40buTJXUKSI9ptro
sLRrujkl6kYX05MiLchOY6Nauz8xzCeRgragVq/XVim8hpNhRuya9IR9wrbpiqIH
6YNKDl4Ce4oTogXN0AbS/BqDX0vuy+gIfQ0A6AAoXbWrFbM8xNaIwsb1GI4AXVzO
ggiSpOIoFvC39oPHJuDMnZpzz33YKrmVjr+n9kHNM3yAGOm0XfykiAaBHdArvPtx
60MENaSL9Ck88JD9bPClGibb+DJFUjpFoFAxurjBEoewaUvaWt7u7KYoZMBxDOIr
fRqGpX3LnxnBwalrKZJAxDAYQ0A/VX0FoqYp9njmhp+inofDX4NDZFpIMQhru/hH
fUdUZ5caU52Y+l67TR0jWPORy+N1Zen9isGoeME4o670G0SJ0nhEVdfifEabMxl0
0zWmoFn9w5RSGIkrNq14Uk5G3YNrJ3yrkysMe/6A9vkzn4JKk86s8o14TSx5sFz4
jt/cyGi0TENoKzd9FhnznyucjGFhF+heqreLzfn/RMmGEz57sGwvqa5jHAh58qbB
/7YFa92PqhRbonOKkCKndx93AN42d8IM9kE5Naug/ATSCdPrUvK8l7YJlYLF8xVP
z4z/GnxOccnW1Hreo8ZA2EHHW8vwjyq/p+wXVL36crFbpE1Y/az6hsnt001+lCG5
98vU5FH1m6aqFInJi5KNsr4xfpHQgJrTd2BNyaSIkVZcouBa54IeZd/s9DPkeD5D
7DNsPMElYOO8ttU+I6eokRI2i7GxMY6EFHnRYz1fq0Ispwifneh+/1qtxOtWfZSS
WBWuHGeBHmYYVOHzbA/k/0bURA9VQJ9/sBpPJurQQctoENMWd5ibMGqicrTQC5/a
TT4KRprNRLE8GxbFLnO6aYXEHjxjz0je4839qJdu71eC4fz+iIPnmdX2D9W/PDnY
O8RPtqRLt46cinx+0ptlTbyytJsTRt0TtygoyIMpP4F75Eulp9LUrwz7rJOuBwwe
lju03HuyiOomm2c8Ilj8JHVkT8ozrSturM4noZ7sW/yZlAN69Q4s5yqbF5Pgu/fV
lIQE+vr/ECUFXsu18RPCtRb5klUX1lkIHfQi3BxCwXVI3+834tRhoouhdGGAx4Qz
RAD27wJM1Ow59la8SzudxQPz8cnNs9q3rX5hbDPqYosgfe2vUaBWsZyPhnsw4Wsh
Gk5qYVFtYNo1DaHatEEpekNoh173Yt1tf4PEksmrXu/bmriQH0l9MTEimjeFErG8
gzZqKJgVsKXXaPoahP4pQUDAN3Aa/CRb/3H5poSaoukfA8Gx6CZWqSJD6ISnzIVR
Ktp0k5NNnGwCnJ+r2CSLjeRTqGZspAphjvUpAogbcUdfHUz+D97ffsys/QhAyQ99
Dr6e2K2VRAs69wZ/8IptHZ3bHLrwTV9hAm6gdi3bONaKaiu4D8kOn//r0b6wjUIR
rry36vvCuvLCwylAlcbrPTfHhgktHP/lzf5meC+9WuZ0hE15j3fdgw97TOi86T2C
pyh/D0PPUPkiEhEGSq5qm2UMGAL8zykNe8lCP8gSlNJyQeK2UsNieQpsuVJdbtax
FNjIBoDAiDh3xntV46tiu9iUkNSvHapn/Lamf2TL5rq8DQbCYzZJkTmxdY8lns+h
k0ezRZpicHqNBGj9vF42+9OhYPngcONTvYVCTTYo2ckJ+LodERNFS2K1eBVcfOKh
QkWVM1k/bra9TuruhnZ8bsslJdxqXDHrVL3zOZOpAO2BNbzo5zLjs0RVVfVhKCpy
5t79Ij3E0vE7gPdUXf0AIBoPX2O3bWFd/TBI6kYvU/w3MsPQQWn5bv4gb9jazA7z
eQdZsPU1pFu9N3g0dLxvR57hpV1cW3M3pE5qs41rIpYBjc94Q+tdUx7+/tkKKUvu
NW60tHHLxyA6aPRMhjEXQsptzU2LJqXKWLDSkpCpC5+7fjebaPtZ6h+DSmzAKLUV
RULEynYo+Qsxb43gBFvMRx3THSymUlOmAKr229BoQOdds2FByO8XyLCIAbx/E73q
RXo62QraUZrhxZiOkm3FeW3/l3Op0f2BXbkFeRN5v1KEPuggPP64pOqTexMF1Pid
wvy8h+1i4/L6UX1PiJWWXpa92KKWlqMiydnj0LFQugx00zdP9BUOJL49MSwBzA56
0M+1NNGAnoQKYEAcG8AU/Ba4gvt19HJ+8ZPg0P7V7hJb6Y3XInJw7/Gqcr9m1jiK
zKRQ9fcelE+Y1WgCnJhoSR9GO+EMkXGn9SmU2axD4kQVUWa5AGjNK4QmY5o6mpxC
conAh39CSBHSPbVfGhWFSBwdCC/7jcI9Nnmk9mceUR2epfS7ATEamOhMfx7jWCL8
MSj9l/mfU8Mt8yRKeYPFIJ6mvNbfK1OLVSblNyGl+OaOh/yu388VenvTP3nmHppp
DbPGwuVfKreysAvl+LPvfCoI4FOh4z+VXrOB8xeBrfL/7NbgBUUR2kEgpMPZVQIf
7ue/MV3CdV0vnG+K41Wn9jx0pyNYJ29Mq0oc7QzKOJfICFuGw4pK7ymAHB1TSlwP
LL6euvUafQqjcR01nJ9lE0oNxH0NtbT3yHUVPj3isk8c+dzIrBDesL31O9WVST+w
5ZXdUQ29i9C/tvBvz1JFi3eHSEuqqA3FnmiJjyFrKuEeK6uhOCTCZGs8/nTpHliV
KfHWtRFw/KiCIbaT3qFqO1Cnau2lpnzyX6H425UbAwxQLMMNgy+TYBrDJs5uoGuS
7MQ23ONLXPj17CbCrainaIQ3o05wUz6eeRF9dqj5hX9VZQAKMXbPhWSI5aC79U1b
byMIxeoEEvuFqShFqghL6m3ovDP41HpmMFQKPFsD0UQPwLzTmlSiZCo62idnp/Ns
96YUmkDpom11gmEcH24iR99rKhtH2EpsYBgRYzLyx/VUI8r3Dma2bbncofaX2y+L
nVY8Qu+N3gthpsr5hXbrLePwo6mM1mEWfYhTyEmv6OloMN4CttEViY0L4IFKTovx
KugKsaSGet0+1mmIYLAtHXJGgVHkI52ffU8jR7Lu7UBdD1ulnj5XjzQtPYm4bMCc
Ft5EcLwMhp++TJyiEFiDWVgqSc/Vh1MnqteLpTGFURYyw0DQfAIwQjb8e7C22aUA
+Ts+39dYhyDKC95tCsaKeueTa0+RkXKg8/iTZDJXAyLo3aNDtYXBN1myzZE7+TCc
WaDTCHYicGUHHRh7wf7dWS0Tz76fp4ZzrbuI+SYYxZ0wuDhx84SqAAn6dsBl6Ug+
ULVKouwyKpzoXrRho3dSrB+c12W4oeBNs1AqDF9mGhFl6wXpUqfX65SlalIINx5o
P5nUOK+zB2m1ILyGWzBuEghSoIzTGvW+Ihm8xwFVbPmy33d3qWe5kAkQeLmVCv1N
jF/3qyMTdlequtg1qJ/SllMSEr3JuzdXXm6R9IGuy8mW9wG8ewXoi0BF2JTJboGa
ZMpxzPEBX3aH2+TGKt2yxol4nhES1rBkwlQ8BpT1inulvWtE4snjEW+qZEaGmRae
84Gh9M/CKtNRpx90A54612dYXZfQdbbqCinSAVvESfvhB6tHqdOtRcEfmQuAXNQl
8n9keUmboNiqFTZ/xguCWHIODLEeBxSTXsn4Nz0iofUwGcnPbTeu7B9DWpi9QmIM
R+JQjsJWzlKgV0Mkw0L76/0aQsJ5SJV5kwMb6ssQ3ZcGALJ2Cbk8dZYWjMeHrokG
1TcMnTx3iWq6Ly2+9I9fC2+BvahE+8sYz4GE4UG/xv5uaViIP623DIwfeO7/XfOA
fjwXrfAwvvbmdRdR3e+ZjIZDbba5snBSmui+/sDMCeFZKT5WFo11LyEN4gLCBu6N
I2I4LKe8EOvW1ML4B1ufor/BFRyzi07Ee3A80vvTACvlbm/oGQ7HAmPHinV31ye0
AmE6NXjNqP3aDx21ov90VKVgAa2wzLfM0afkt9PF5olAs+p0V5+HKcGloyhUAd1g
Y3ZTqIFogyFGwv+KL6COiYRpd9CUZ5i1arUQ7hReqcE3ItTP6TQGva5BLX6m9cTd
WmHYdxjnx0t/BMinhiSqpwuwdm9xuvBFVYDisleF17Q3z52c4y6Q4z7tQqm2Hg3E
IS16Y6XAGstFvMaPOUEHSd8yeLtPOZTQZNWe2bzbtxFePbYF4DMlcQXgWFOTyEHn
ziE073nm4vKlmt2jcilhnVU0KkYYbB/upTFBP35anPKdPeMpLKn6COKHmq/K/PNe
ankZDOaYRxIRF78eewYeb5BytxCUUqccbBh7n1feszCcCiAbnGqIWTPSQylLT7uC
3AHZdiM/BW7XyzZeY25+sY29HMo+pCYLzPG5Ka1seVzD2fcFRoDKpRggySFnOjPf
u2MhF84cLv6NjudvrtrjJfp9DYj8s3z9k+TuCyGZV7BbVJsCRlJnXWDTHset20uE
ZU+WD7wVsEIyLJvz0lCjhNr2hhpDrnZHZGdMdceRWhTavD/ho2cXj+2Bwi9IEqsl
Dj6vhqvDaNT2Ok326YsmdnxvhWc6xaCSkw2yUyrXnxP25g4DiZTbkp4yb7xOQ3af
zwtaRvU/w6rh6QSWKq6Edb6B9LL51DZhfOrmzBOfLf7MhO/TbRG0P0zjJr9F0k37
dd+AZMXewBHZQI30LupVY1jUnroUo4DGUCkpZ8jGcJQ5JQHC7lwbY/VlB1RHZ1Jj
K1yWm2PDyaudRYqQQz/97gLvHwRFLXtK/mPyA5YrW74tpQtmt1bD1h8vP5vpBDrD
lbFb4zlTDpF9/pkFlYTNQivvXoE09gTLsiBweooGchBe88s1d7ZuqWxsL/WsVfqZ
CDRNw1YRH+bkAyUayv8ON97iLFXoGg9lm8pOk18pEbUg9XGgqpoIwkwDXPblNNOk
iAjGwkdmERm2S6ohU2AG/VRF5YpwLwN3Y+0t7LeEns7cverS0SrGCyi7PHxMJHPv
vi7CX+j775N3l50ppOJ8jvinVLFiDxEuEgPYY7HiBKXO2nYVOgkKrnZkFVaMM6El
rqcHQT5DhwUDHKMppiPB63m+chVABhdp4amTcDdnakGOfwFOqxmR2wbdx2cTylSj
f4gKzQ78NIjomeI4FeVrczRDrE6AeTjFkvA92Q6Cdgotbte2ASGUD6G5ZKr7TaBM
0svtcUlG8PCTlVtSrBGmc6nfGoO7sWWNh2ceGGpR0hnOMHEEwsDI2mlVZTSx7Mcc
MoOHEKgrTYqo/mMDbKB+0ugzeaT3ZuO54Hv/Gca9Q5SE/Mgm1VOwsCNnbp4m6Gps
vBZc5wptPv4/bHFDCo7vEvVIwfiYyyTF5ozc4Q2zb+A3F4lvegZg5Nzn3R/hrire
YRX3YOUt9o0n3TRn6r1Y10kAvLnPfBTnNBBXtAsEv1TEwORvFWcvVrsy7Rhp73UQ
s3In3olaeFfRCar0bFOH/+eM/cTdTT6qbrnY4QiE9f6GvrAgyxCSv9W9Y+gt8y96
IOPqd5eXnJLd9nOzIhLgX+07YoDhhI5Wnbi/0Z0D/r0TcEAaICh6VZMxav8wDyii
a5VOe28RV5jkgdc03GiXkY4yyLjWbmKkiDNtLUDeH9EKfHQUq2dr6JlsrgAHN64A
uAN75eqqat7HBaPdVXls1NsB5XGAgyg59FIZ4xbBYfxUpyNrrdydHOcbq/VYOkpM
zoMsDgROcovm1waRrnI5G2F6CtmSuYaHmPhg9eIPGPQPteSHsV0eYZQNikWcP974
ARMCruTtPlTGZyTW1B3LI0TLFp8MsbXM1eGO4uPdtfZynMC5Ik5skpH8eX727wMg
A7dcSna04LR4r9V2VBcEgGa72NAuV+6xjMXk9j24US1XBMk5LYLGq41K80aFyKKb
9ZBA54M0e6HkPlxeDhZhmtKY7jwoZSurGOw/z8c9o/L+F3iGolwN8plQqwUkyPxy
v06gjuSeuu8cmtoyz0mHU1y6nnPn1EFXaBEFDfD8tO5E5JWjbKiwm6jfWIzkADe8
QyW7r1cVXGm/2Br1548L4RCL9nxCAOJX6akfnJkxOzUrP8UCUGtfQhaiLh0GHoPU
ag286/q+BSH7hMMfOTLc6JoIzol6RYnU+cJ5HQ8qkIuLnV7jyoscF7aRvUhRvNHy
SZw165jvTyyAlgtZDK4Dtkh6On2rnOOgB1Thjf0RBfrTENfNkWDVci7uDgRi2p10
uMQV454AyhzefRo8vSIOJvTL5FqBizoI483sq7Gl09G3iWbu013iNrrIimGs+ga0
MyH137WebRjWY6zSIYvhenlhPlcgljpC3YkAqm7lHthPBsZ/Lc/+qN1y0WWG3+rZ
j9fpVg0NYeCy+z3mv102bauWsdvJzI2WpN1JjoLDW3FqJKPLXLypztWMB7Y1PKN/
aMH904t30691li3t6AQp+NyJUDRTtMqJY+I0dI/HzROUCoKA2g4o3c3nh4qJnUnn
kbu7ao566DPd662OOMleZkZ/xTrYE1aocBwX/Jl3+p8XZLon6ThpNPqPxkdr/NFi
uDVf3ALqfITbyC/9h2m2xvOwoLv9ydEgEm0KzEFXfc3y+zBcNDvDsrpzIXDHdeM+
MbJ2Gqv5PMNN4yyRDERHd4kLzbliQBgF3EOu9DIsNy+YTonVF95nsU0y6pL69DAs
4/LCgyiwhJyi521Y6sb3e00+VplDUAhAirLI8lXHf0B0pLXZWQ/unwXZN3j6pObS
NifQG6l4yb5iUanukNJDhsl+yqAzoouRK8pNZkVqUZYW2BmTFC3iGy/nKtgXU250
vqMESNbA6EGYLnHyhMD/dXotkmIRtwKkSAqPmvEV8BIqT/rHEqpsptEoMcIuCSzm
Pl0fQRN9CmywgSRg6flwdDd+cjrI+NY09QGgVcHb6kG33jkGqIH5X1yUEoM1QbTT
XStOdjaqixEraGp+SFqj0P/2/0qfu33Ga+2kHBkpJ5IVqBuJLJ3EM2A0Y32FoU3F
Ym1qiUz8GhJV0R+GOBqQFquBoQQotztndFXTFO5Z8t1LoDY+nkkf/lN1WaA5nvMu
CzPC36jRlZgUcmUhAxCYHxC199Lfd1VB/LtyeDYB+kZyZMGG6HSnpDoSl7GOALNF
C427vO4+LQIszzYE4LERDIXmAzzomwpx3P19m2NWU1ZdSHePYhh6JE3LuGiRnpLz
g0229mNK8Pc39v+Kay2HTOnBVdkXQ9ITXqCC/cJbLIzGKrL+JQKm/yd/czF8qWOt
mgYynHYyUm429scOsc/1ZnMlYszEasJbxpFj7opJdaOKXgbTK3dG77vWizGHNa3Q
oYjJKdXPC390ZtL3KVlB+NAnU43V7iX610Ky1gMeLtbwawhD24JhfG0Rvd2GI6sq
BE/n9idKmlv8u+nzXHqmwMPqQzW+VnYLz90wEgmQS6mC2RMCh26l/P5ECtcUBbJa
MSsBFhAGbGlWsmFoCZSZtdGGWITZXfg7LVEDWAozIAwwO0lzL610p/2OAibsnbs8
7OuxonxT81cnLOnoPxFMQhoU9BllUsumQFeMQSruUuUGErStZ7VxS5ePGBqOL9LI
KTXJx2Aa2n1uDfbI1mBBOL/6VfoFITOCAdlDso8kkN9kZaun5wUO1rOMpPCktkzG
a4j3L5dybWQ9URAf08xPYGcWtxPpcqqNyMQMnVypgmweM4v530V5zdf1Oz4aoWrt
e4Dm8ZlgJ/bhw1CvVDrQaIIocl7kV18qbq3i+zw9bDzVss3CWvSICveAi2D4TVJl
Il9F5I0Yc+HJKfb96Xrgu5ivRc/5rhf4cQAhAYO32Ka5AZlH2phmm+ldL1vwmTI8
dW4hG/nXrnJsHEBYq7zQ8W0D+t71OPVV18LS0yKB4d5ntmpsTX+h3xjfyr9NqYs0
8KpTvCFwA5Y+hyxajoBGzg7CfA6V97vhp35sMKZNSH56Ob3H5DIFxQePho/qh7Si
EsWFvzHNgI6+dt87x4CMjTL0kA8Jcxpr8iG5rJikEGO6RKo47P1bv28cjWtj9l13
xhD/+yKR8Vqnm2tF9Qn4AMThttR1wdkIKaw7rNoqspyhz9vHHKOyJL/7VogTmwt3
nOrW+xMT8+pnwq4mz/jSYk0HdXl8cU6xulN4fG/pD8g8ie9XH4nRfq/yaiV3B+h/
BraU4S8NFmugl61weEDC+XbJz/OfYhHrGqcd6/tA/yH6fe+KUTgy/tQSlbHfQcIf
HaIXjnAD330CvwUxENkNrKD+xPZXePRqkTuJH9IiO+f25/XkQPmwxn8W0yyKnAT0
/AHsIq1zfy1kyHQcIem9dV6LgitbN2Z5NS2u851zncMzukrEnKHzCsmUMzo/eFsr
d64B+MIneh64/D953mT5d1QlExOAuSpZuNSJk8y1qyTkMWJ4OtRV5GXoAWH6iZdQ
IylkUkWVqykVFh5QvAJ/VKaytcOMhPXPK9rGp4GDIoQYecYAuu8GFCigLcdbrIJw
wsvkEcHIrdJRIi2Mjzljf6D01dQs/6YjvNe1Bo/SeWzFCdnvRVMifDFoXS5jtMWS
0HEBUyntrqwq5MISrDpM0WHXlBcjkR8A1WSiYg87ChS7DDkr+goXhvyTHQkCuCiG
rmliUmieZTyDTWE/LMBB529S9INSF/L1udhpEZInS52x7WeuwJ975V/bhrg3is+g
CItqbT18GuGYywbMGVOEJNXUF7JWFTLmYM7tk9bfezl4BRs587esVjQbTPcJfnna
WRfJxEQETu1mf6xIkXCBiYbbj3zbIm/LT0Ae1yol+kXh30AHWq5fiEyK47uSZexZ
SJOj9eG11nfM1cidQjv14i2uFlv3fcE3v2aDhDLslRP2/h3cvoJ4hHmrInunIBqm
U6zYVqyJ7vb21xmslImz3kXlSe8m27bckn3tcZJSZ5Wxg+YDeC9i9SzNeMaAoT8q
KO7TJB1x3uAL3OnB/+0GuFTg0kFMCR9/dm2atTo8ZXWHzKCb5cLSY0ozQy6BkhNg
ijjywP0G3WgFjQrTeIvfRNlpyDPaEgk9r9ExqKU4tyUUCdxU3hvhnYvtNh8K6r/a
NNoLCVVvaTx1z7bG1MeAdVFwmt8C8iGzNOuPnsUtXJnTbpwMui6h3wI0gZs6ans5
Lkexy1inKJZSFdkvirNITXCIn8KI05pfhRs9+NJaanxu1E61Y7ZHCHfRYUGpO5y6
fzVa8/BfgzduAA0m9FxgEGJ8V/y/IHJS/d9/r14tr+aXeYSz/Y6za3aLcTK+csUp
HWQBzGzrNxWpJ/N7nvvdXr2Zfn+7mZRlhZFdLXXkY3UJmjJVBtffbSZ6GTy0lev6
xrq6tImCf+7A47mPOGrfWAqQ5+iZNnK+t6Qhsfonm/l+FLebtrSOlfYU5KxvHtDn
ua3Qnpz2GSkVlNJSRGzydq2NWND3HCOtBTBWoURJY0WUvZabvPD5TItpdpiBaDHN
mcnQPLkAbL3dph3HkxZt7eYVc0nmAIRJqAxBGMXMGwBSBbDB/Q7nbqqDYia0ijfm
jT2HF4w3npyzyx0pCMlIa9UG365vinTuXqyd4d/ur5EtXmsl4zqpZwFOiOgyB5Mg
ntJg8UBhzB0IhehTysUqSSNUezojMvBOYyMTNh+cN7Gq2yicQBVnJGwD29Q74Csh
IshZx7sONJzVWGpMJPuz9K5+dvtUcKGB333ZlvvFaIswKx9MmzcutPfnfZ/szurV
8v87fu8qy1eR1GnHMW/4cSn8ygYnePrZdB5g4on5s0FO9MJijQem0qT1qOJWpPk2
Jc+FD825o71QWZDo+N+H8bWLCAWcmk1tqdjKLP7LH5hTdmDoSNedZzlVSrHHjwx2
k48r8oQIlDs6sFWE4Huk//lxo4mV2qZ2LCbE+s3mzY/XUyQw9HSNej285GQqHlf2
TpQaIeYU4QNC294vNW/6LL2o1ZvTSoGndTQpPnElDk5unnhekRUj34U1bj+nBPxZ
ELIKL96V0FdWxmcjlVABoW9iQlpVpIAr6pjh0lUovFD5TpigikNh9Apg84aom3Ma
9T6J2AoYD1kL3sCohMe5StP0FdxJpYUfsnfnuH/BV6VGiNIdasq7M9NxhvPdKKyY
P6Kj+ROLxY71kXIcWKuHrEEujSePYGrP4UhterEWp/wtWIGsZlnaNiM/Ov6lD2UU
J6U9euaAihURd8XwUCM/DiguU2vRWFH9U3Y3sZZu7d1fPvFY+jemUNqzXu1AE2FD
wItQAzxZeq7999/ELFlzv8f90nMSyyzX9BSOOFBkHu6jVq36XyLhZU3nXhg4JUo2
Tp1fPnZBVEHI4ZnZfB6iRWUid34YJ0NPbdL7ArkfveS6mjN9vBLv1MbbvoE1IYJP
u5OpCvYXRi5dfZBqHb8oeAVcvxwudNS7mXzFO8tmAUDNqhe1ox8Pr6tbqcvDXtqX
c20Hoq96Qjy65SdzkEicB3Lp+k0gtX5bnEO8FZ8uGOfuTIbjXbPjIBUxkTl+hiOK
s/kL9XL0DnklWcnAzMDRckaXC3bWusDKeRZ7x9gfYGCMtaxiFhKLqmdxdch6vg3K
chYQB6Eix4Z7+c2BRdccFXsONsk/2Hlc+LifaFZa9uDA+IT9V6FWlFMluXcmnype
6OpEaLqxdMkjOCS7wdBwv5fBlMY+4Rtz5+TtNXpyIh2SVxPthLu/pj2yh3AxqGi2
iUPvBMWZx2ldawMMc5jR9i9pzTAjxbss0TWJSJBB8uRKToPaPlvN/ALDi5dCQr8w
LKGCdFhVQeVfVYUl4gvnyremY2E7W5IQWnaXg8/7Zeha1rg5JCJQkSfbhLsekVfj
BxOf0+oSPoJ2PeiUMIFfGtphgyYbc8dfPOoh0Jgf34T5Tv+G6kM7ujOBcvlH2UVc
OFtAE5Gk20uwhxxJL2OvpNUvZv8rNFXWOtDMJ81NQiBt6bsZ3zEC83Z68m9CyzIt
ErGNATV+Je04p7IYqnDqEjwdI7Qsm6MAxTDel0U7MGkfQj1RoGaSlQG0YXI1BNRK
X/U1htc0tKcIuZYDrhKw2XncRybrs6R8maYiUpia9UnUWGyz6Qrgt23OwLjs3XxV
jH/aOWnXM4LlYkOUOXDtii6BTRKNZlDeIsxUm4BaULUnRSAy9NNZd1OYrPgSNWfg
WLgTKwGAkN9O1uClmHX/YW1K9G91E4//tgkZQ5qZwuTAqfJGoTdVXw7kHxKHaeK2
Doms6DlRNY5AqxxvrqfU3V7MCRFQemB0jaOR4DXOFWux6RJa+1YqnmdtG9D0/R8r
eRDk9D1HXWokY/EjXIuQ8/KF/cBwWWbdrjnKrShZSdYN8b9MGvrQLgIc4MtaHElE
ODlpqtESpbBh9YJ7BW3kyKxOiEAZGibz+o9lR1FZ9mZmv1GPDSu1l+CMdIWWajFn
ZGdljKQZJy8J7ImyHxoykcFvndxjJqNoQ2lpy7B8VseaUjsc34esOWjQ6JlIiBV9
YUWNxEdcQRWT/djYQ9L9ZjKJ4YWY0KkMSLLoWCBdqm5uv1MsSm8V6w4VOkOtNik+
6vB7lrixriBVuZD/ms2Q7XcsST+sYoFOTzK4GPFVE3ID66EiorCmV9BhLxwgyKX0
BGdir2n3+pLoZ1utUbqFkiDDITKBmp3Wp0fxQJhRJ6ETjfQKWsur2C2YgPyl6IGu
/9rxlfLet4eNy22AHea3JORPNjnAkUhJ3tvm4hzGCxaZ6dt0Uhb/tSie4y79V8NS
vhcU2RQPzZmsjvxobrvIIenRVAJWPJHVv6uQluixPG7K1VCEhDpZDmcIDsrghuYZ
rE9RvGhU9WfgoEGQF3WXF3LqbGI6f2Q1bo8XeiX1LCDMu5AnJg15H828WL70Mqrx
TqbyV8PhEYa5vI31KS4HhAqp7BtAo2R8bFBWk9+0mfGpOH4kwvE1/LHKQ6i+jN92
7KQxRVEAVyBWfhcOns8ggm1hWkT4RbBPm80525AcUeBJc5fCdmqq1YLlED9jWkWN
M9mQ038b1WBvb2oa4dQIcWJszSCa0IPWU3UI9jxx/DyWnmTcOqdWRt6txJM5uOw+
1wRBy3/7i9qG8jhQSZf7dstqDe3YG/xdT44AEcWDxcxNh/UqRiHF+VzPukniSg37
TOZZVn69vAa12VKJ4yMbKX27a1CnxfWKJNr/FyZkdRnYUJM3jLaB5B1wVBzcsVYD
WAEl3tO/Rpgy3gWQr2MBSCGr81JkrmgqN60DAS6Ic0+eBnUbsowC115OwQT7786Y
y7ZQoQZeSP3Qdo/2rTxUA9s9VrRe6CXAxSQKAQbOwOQUbpj9+215Mrn7ltpbyIuD
b92NDVTVBbwfC8nMSglxQNDokgEM9o9HVbRXTXjFf8eCO1mkqyknB9zE7iDmaP5G
sZ7Iw0TJLEEFiF4kU5rAo/sfxocTuxj44CgruVuxGRjAiNdMc+P+2vAMdvBHD5Fb
fXexTXfUGkpFGTCcjs0W0/NJNteh/oVxevKY3Rf3g8Z8ezjYqWarN8Lf7mULxEUu
nhIP3pAXzpwklcfqTB0efX5QjODFHpdnz+AkvrLbd1WZXJlkcI++unNU+KCDNI1k
oJi8W4567L/Dsf8GjswK+Ia6mFI6awIzd/O3uJUfMC2wzEKlBAuBhmEsMA0c5w+u
nv9WhlZgTJNUM/az1AP+X+I/3sYcJjZOi5ZyulUURnlkrddPZXDCx07idiBP0AcU
iklpDMQuscQnMTy5LMTmNy4ePWTv6cmFol76wXIVZEo5FtLVZaKzh9jFSHdN4eFc
9LGOLF2o86lpHmIFUGxCUiy0QqI8+KRqIdNQwOEDRNwgNigpDSvS2lUC3rg9uNLA
PWOKIYsa1WghehpkF/CuY2qaiFCd5waBt6NSK0c6R45YaKx8AfyH5AUIKqg/zHnN
sa8Txp0tVjFZasl/B6vGoTB5o4WFO494G46ukypP/U/HUsFoCtZSVRT/bnmvKycs
75fOkwYq/7PE+3cvDaY7c9cufHZ8qop8mCRhD1L3ZtcQ4BtMCcHCQFSccbuxZ94f
XZbBriwdaHq3W9HIo87SXRnx5qozT5R0SG9C7lbBIGF4rYyY1GIq4o17C6oJmpUN
3+BYRu6XeFFWrjQgGju6ALyzQXLNsEPnHmny937HxA8yv0PG/wH+asPbcOc+pJcM
mqHq3POUU1vBnLvWChWJLgbMiChsdSNpZEYMHnHOGEBrQfHZEnD3sh9JLvUy8TOD
pcm8/ERvAwwtPz2ResJVXbZIj5vjHlkLgboBV0cYUh3T/ggATeHGpaPGwCd1ssCs
AvTvijb81Xy9qWFyC05jcpFh72IT3BuNlwyN4kWavcokVBjdslngXk1WyyubNN5C
2Cb/LpJe4gEZPICmW/Z4tvhiT26ucYp2z2M5xMdUYMDHt9OBLJtqUCHC8f6nDyqY
b30NC7wLoZL23VMetD5l4ssFg3m2WGygRSjHxhVfzQUSSstL/w46MzCOPSk6xB4i
3f5LKpCEcjpcfo+T+Q6cxFFtNZKysUYg2HE6YphLkv6FNy0hunULswHtKPGEOa6T
5JS7M1+5FvXnfGpCeGu259SNwj2oA0yeIvw2NGH2ZcWI8+3tuIqW031cRC17aigt
xGZhj+f5XLm94piyEG5uNyt6AUGbUdcXJMhLGDhcmg7i5jmUTRSMei4un9icNNyM
ob9UW+En1BNGKQn+/SsabnLoyAjDRdUDY838t65Ioai0+/p4q9xdIfJbI/tTUlSm
vHj8vcORfP36wngWNvOL5Cb0xMt/X5UEd2TvDj+CRzKS9ESonK2Pkv1Y494DOFh+
aFMjro4wtom7ZlcGj7U8zUcPXEGD8JjrJxhDpbck3Zph+wm5WSuhxUY6irVM4KeJ
V7QIeuYXARWgMe7SXJoVRP+hejRWZTYO+C7Dnm40a51eE345iTO9fBEGpUdPW5//
Md1ex3fZgnIMKKbZQNT8u4i/XIZa7XxjxOK6xr8HYFa4pgIVjABwGcpfLKHegnDI
ATH3gg0ZqY3KYyGsPNMdgdFoZAKKJgmyfS1iAbJyJWDk3UstHoeU4y42S3S4ftvy
OlgFPJxfAg9s0cEAxcfslU2kllYDtXLap1k34q1tiq0mDJNYbVn1yRipOxd1cYNt
9R6sVEuJGR2DDHqI/Ud2APqBkzfm235vGqFzAYUGO8O9TOTwKuvr8ObCzj84MwJU
ajHs1Yw0lWsklAmbg56A8CCnyHbnjGiEfa2VeNOv78quYrYG2eZ0wBU3Mmwgau4v
Jgz2Axiz5dmbsY9rURphbfzKGsUQahUUdMNxewC3t9LP2gOYywako0bJs3wJoaUQ
2wr0DmJhPjN+LmnY0B62TzhrNm+dxQIC04OLGyBbSZ2wqdvPCG2/TgSCyvlOSxs+
bsd9MgviI+3sqAx58w0wMt3EhkyEus3a4J61VfzSBkK/votZn5cpEirBELbhFR43
VURS7oc3DFVmDjMvLk2EXCiOOoCEweZZiaVc+LU2u75yOC88ohbKzh+dkibY7tGu
BLgKUSFmuWuyKk/rejbozoHplzNwdkTglQMcfFXlvpmcoDnTRyXSda9iJpzqCwci
ZwJA4wboPHlq1HmOfz+Im3/uBH9eW0MfgR0ZyZJtd17BH0zK7iiV3Lxw9bH2bMmI
1oLlUIQW8FKmNb4VnwrowDTBzQDfwlJngv+eMYVuJ7MdRvrL231uxX/svrDCYj0J
C3KyqbPHNngoqORBNzvmiOJ93a43HcqA5VsOoy7LA2pxiov2hBm6iO9fMwNB2e+d
j7cLjsodAnQAMyQfNYoKqWBDFg5yX30PcPJTfBgVajKQt/wTk185gEWRblD1wIoK
TNDgmtfu44FswbVnJuYnoX9aVopj3QWKGs0OyDZ+xFfJftiaeZf6ErytEFrpyW6C
yUBIpQGV9Z1HnqTC3LcNg7bdZuBO59QcdwLz+NgHdTlTWFYr4uNAOmg7dCVWRl1r
pJGiz7JaAwdwRDNKL6YAUDTqgRrmw1fcDfLq0RDxylgm9NmrbK5rP2t8BUmlvA1d
fY8xMn+8UGm9oBVWJGm5lprJ07vapL9Y6jwtTc31DOHaVHM7YWT2gXfEiG6QD2K6
9Sc7qlqhBClPE/8/Xyb5C8QM9QVvVbRG5ISWWkYOXvTdVl5hmAucvWuBjCBOTlCF
9MVTQOTyACp+aEtQ1JZ0FEN9ofyGMffVfV90y0VYIVfKGzTlD5nFHYmSAZROF138
JWDqUikyvF2lWKxLZYGt1YAcL4f5n+UNB2j/9H/2F3XSGWoYpfcNkJXGkPJaxo6R
UFR+9IoGv89pRYrTl9cAbGJwZi7Lagy9VEfq3xCuuSEUwWWts+3hS0lYPpfP/3Oy
3x9/8uftX/GfW1yr9g4cN0dn/PqEnsgMOnl9zrByyrcKoO5otoLC2tXccDjHlBQN
Tbxoecuu1v4e2JWFCqmdYTDM98w5cWpooHUzDFHn7rbSzkGKJbkL97npgS34tATA
urc4L5IHMwP3H4DzP4RYB3T3HUgaArXTdsdrvv1FBryB9CnTv0TOjdJyGUEkOBmt
Wx7x4m03ha1Qs1loUwnz+T4lwU/0/xdLYFAhv4Zm0Nsrkx946/XUZtNx+9gUptrw
2FXnAdA7kTC557tXs/Qy+4ZHIlmDi2VmSvR6aGSOVK7SjouSehlGHQQL7P7kEwBn
mHvWZGLRZ90zO+2NF/fh6XTRfmWOml6+OnBQufvomwhRu6jyAGJ9CWjwOcvEfx7M
E6YTZKVqfe58/Ti2ZmYJ7xX4kNQOTjvI//WGLTwB6BMCG5lvPmKC+JmCqey5BuQO
DHiqxoEbElhhl8r4dKmMaz5KQcvKtWb1q8DzHIChTBrXLsvQGZh0GEgDxcY/GUZm
i7rwi8nS554F2QyzQB6a3fLt2+XQN+7qbJKDFav2jMxVwA5I2aCyAciqhUprsvf1
m04wgRUTq5EPNxhTl5FQiN2qceluR84ltcIt7X7kcdVCP2WqU5pBvb1eCE0/lbQ/
Gwbnx3VpJCmYN31hipQNaI8+ipnfY6IdJwi+wlkpuTdBFhQqEFioiDDt6GbhHovp
0MjGX98QBf2z136fTFSJrFLiUoWxmIpse94EFM6sQlRgB73cYH9Z0NmsOQPGTTzo
V1Htrq23MyGCxXVLWQDqz9aKJawb+kAwIl3tbw3DyIGEvmsHg+UXKenuBm8QxEZb
w7fhZmj7pDWEMZraZMCQrXfhthSiVmbMds8D69VycV5Ux2VN2GXDTzdG6tsVMVQD
wRYPVWJWHxRgT4R8eSuZk0pO3OQFEMx6sBWktwXbrAiO7HBtQ4yjVKaK4W5KGWYB
DPLrKUn2Nx9Eh5b8J74kyJgMO5xVqm7BsVZ0BW/erK7Jo+nDYmRtFcew25oEWuD+
K6ZLjcEolu/fudgpu+AJ74FVMykTm3pOsmgEHI8QIDB/QLDl+BsOqiPw84EC8+AT
o/6vrjGVF8+5qsv/gasDv8DZyptny2JhA+jHoHB9zX2GQqASjGE1eCezpr4JGEuW
JLVJNbUvo0KWfmGl8/E0J/qZZV/Jf43h3xzkAqyrpURVgC/rm45Ce43Nh3E5kmMm
NwyOyLHg5jJLZJnLqm5typYlvskzS+hUCVGxthOBxQBEuCO89Xtsz4iroKFrfrfJ
ut3l0xmqQiYCaRyS8G/l0ZTw7uol4ERLRP3Vg97TTNy2yn1X5DSBvUpIn7Mkmq1y
+65RDB8V85QXG7VRCTSAC3ViqS9hFYgbFI0u3Czb+UfyKIhyD4umvoB0pfu7i607
Pz3B/9CNKCsUJpYZKz24c++wGlDR5Z/MNhRKbY8rYquQiqsGEQsfNqbEWuvCQUjn
DO8h1UdNs/3CLdkav+lwjziwUDpgNfgc//GfDy7ZgsSdwu7bc4LUA0JPgKL1nW6i
f2agz8uDUYtYtFKeRLUg60fw+FdEBy11OFxjf7un81N3Y6lZZ7TlfnwhA4UJvuwt
kUmBmgubSkTVnA1KnXdhBsWXRZylC2sP73/2SOc12lfmKJIWpSyFhNL5lbbui37R
F3hAcjHMYbscRMPnQPj33+x4LQ/dwiVACqJsWCaKEme5rkyUVulo72psTWoORhSj
i9My9J6PS4JA3YmDOTGSk7bra1JrVlD3PKLDoTr+x/NLJWKA8PkXK7yLAvEF6CAi
wfwgOkeAaEj5IIRvXvolbrzCFbJQ6AnpDzDo3IgJlEilG4bpMMspEry8HWZuBkPQ
3/ZmX66SzCl+3v7yxwSUMwEpjRcT/lYY3PCmNKMyiP9oxI/pLoz9rQzWxjHHaBK4
vrp7qxk1qeLAr1Bl3/boIQPyZQEokXkndDdjF9+PY+Ep5cD+vpy4uh623+2/Rc9B
Z5OtdfFFXf+dTvORWBb46S8Jz1qBQcVCL5MyNd7Rq8WTEDAE0+O/nPh37pngiW1n
DxH573n/C/Fg14FuRnxi9O0K/yaOdGvGJfu7wHt+4evU9iVLvK/99u5/JoL1pGUn
ju7/ZdZjnV9O9v+11TY1cF8WEOhuU1i71b/ak2gQvi/QdYsVco230yBVhCGNQL/5
wSI0RFnVf5HiYWMnJwoOJqx80H6KI7m/zYdPxPSQ7Qq9vgYYM1b5HrtXaQzka8tH
7/IoJwlQuboG8O7QOv43H63VtsccpzI5VxYmQ4bSH/TPse4MmNrn2nM0Oxd+8pFg
TnX+s2MK25Ee8vkjGnqouRw6l7pULUSgf+AqZkqHbigFvMw0oHG7gEqjHziOIa1R
zQveX/4GL/YlmfN3FVzC+6THpI1WApsu+1/6DOSXzuh1ryMvM/wk5ZrcDp3jDRzc
VLMyAXhg7tWfXxs50+bku4FImobcQdHrOt1rP4QZcN08tsazLi3Knk1WSEOQYEMs
3ndRNmTMMzooA/OFRjnnYbCPCZwB1AxV7JVCYNDL80nnY117o7TgsKf/KHXs+0lC
HqFoolDrG1k2QmsZ/lkCvRzoOGkqddAENNSE//S9Mv9U0aWC4vLDZ2YtIHz1EONh
RDF+kEw69Nr4ofA9muaAArpfsICKmOkJsL2AwtWHwqMsCa7FLz6+SsZ4EudheTy2
msiyIMGbH5j03r3uW+xULh4ylJN/MJUJyCdSI9IMkXKhMc57UqZDMmqqkrE2uCWx
atIbASCtxtc5DD/nm0bUp4JuHrneSaWZtOL5xH6auwTW/DGaI5TC+PcmJo8YCBx+
ymDchCNhh0OtswCe+mT1RTyKPCHqXpHLOMnYaeC/+ZQHVmnQCGq/p7Zv12GafLPV
1hH98R7B9oBJvdizD3qKlKoU10dKi8M7fiRrAU5/NH0vlW90yGGIN7K5UbWIh77y
9FwVDHNEPyKpQg9qV+1wI/SGJUuPk6gSJvFErnvR+1yzGjlI5kSDMlHJ1XH+gpJD
PLHQIta5Rz70s9N2BFiSnF8gNRHfmR05dF2pT0+SXjnimpsBCjWX4CCruP8Fqbw9
Rh/np9V+Ai+BlboMruntsLTMAE8UI7jmzjH8xbl4HcUXmEpq0VlA7dOcN9Qr52ZV
XxCYVhfAcEQlWokU6mTXISXQnm8j97sGXyYxK0+Kv6XIGIlBb8LABFWklJHc86wN
Mjzwlgc1MUpNm8n082UQ4Dy4h2uRff7r9+yylXRqFcr8KKXR3mFiOzPQtRCHiffE
GzDWyclFdU8rS4m6X1mCPXbIudpKXJmRwsGWPDC4c1IT/5c5U5+KM949906mvyfu
Ron8gbzTe/gp7qbvnV9AOmuiGkCwJMFewejbf8Z7DGj9ndiwJwDghwH7NTVEPDFh
6wneT+SGZ6p/xbzpgmiUa036Mx/YcY2MhDZhxUz7BBCrzWGR/UXbrR3IdD1hyi2k
atcpJ93Fhp6sm3rbZlVtkb55OF0tDd4gcqBjRtBH2G93mnJvD64OIiq4/TKg6bkW
3HHjLVbjdvVFwJVcGYwYfmTjOBt0UQ1848r7poRuiAJCJVLsuVnoCAuvMRXWtczH
vR/wvtbkkJY3H8TaVil0LveNf9SDFO5r9TYFIdhkwMdrFcfpn+W58iPJkkJw1zR0
EOY83l1efW4ciVCNcZEm1oGYvy68LrdEMvhbdCCGQWXTDNxup3hAOzLPhgfeso5G
5U94QYTsI2/7ADtq3M6dHxu9GNnHRmk7/7YcsGMobJop3X1TBf9J2T9soPO4kPGE
qP8pyUcV+xCKcXYf9UKNnKJRE1/D4h05xVtr/cDYMEOfVdhaowW+TVniyrC+9Zjn
L2S/kZPxtL9dihobWnQbEKQxpgLmeH1MvWamS/bYKRgM94bQSam4vyQuIr3SKtj7
8YPia+OQ4houFuDPCCS3sqC4NzeQypi7s7lbX0nqMehBwAM7vz5PvNQs9CoRoHwE
IZk+ey/wEc1EoWu8bNH61AbA/z/HQCdYac0ZcButdEcydgj5nX+QxT6RjwfNUsa+
ECNik/2O5kag5vKRgKjwNUbiKdaayi4C8BaZ9M/cWwYjo8VvVduDPQJu+60pYLb5
bndhNQohwIXUUhwUtqGSXEgQNgMcKwgDe+T4c5ZcFLqArP06y4wXpMZJCpyTKZl0
L96IL/gCo7ytIURZReT8lCFuxjL9k0UubQF+utExz/iEiA/2RSG8oqR2u/ae6uvh
fL2t/lq+YHvL36VD54uyMqaxDhgMJGuEVmjpyqqZCVByMF0PK0rl9hjWtuLEQ6II
gy5VcIEEDfDU2KSVG2HLnYrRzQmNaMQAZaNqMpEj7dVi2asmnOkAIK0XFo5IDCR6
MMgdFX0JRD/ZPgONztMcluLtZgRuSd12LaTtcM1s5dBzYoHz60SUw/kAjeXpAiix
44FMa068OcgIKW/sE9gQoEU2N+5Ur6v4VE73znh7uWao5+Ae3HbnmVZMz174fq55
hPIhpjz0Nx77GMDWEPQIlsciBBvdRjNQ/qNueigcpR4gRzsOdAHYnWngvEg8grLE
05N0/u3dr+tcBzi4nRBd1mCwA+/Glm94Iw2a1qYcXWhQ5oOkzX7QA+nbUwg1j51b
irHApq/f0xFB75cCpfZcNHG+ah11YAc8ZLIyx0r7+H9LvSbotkRc4JfbALOkPV5S
x6rtL39YXIxp679AFB1wjf84YEZ2oiV/bkAw0HTC5nUKyfaKDxLW6dq85UNVFpho
DglLhR9XtCSO0HJPs+UGfNnY62+/H6IWG5Ep95iRg7JYR+jhRnq/8FXU94PWsc2F
JTlZT3OmXkSSDqjg/D6y1T/XatLo+GR7kZjFwhxLVOOrTUwrgebcqO0D6HZzWFyy
Y2vIAAx0NT18vnpvcqFTRlaYnjvXOiftx43laD8m+DNmBivn9TmiuDaO9HAonZaZ
LjFrUCE42IMrOHg8lahA4deGo+FJ2R7LmcBUOr235ZwcZ2dwKWrC9O1ZqGXxrAsi
v++oQKDkzsh+PbZxgia8uil+uMQw/Ee1J293HUuwaMPawq3FEBh4vsUhAS7TBnvJ
a7atPMueWYu5n1oV9tlhAcIPHpzUIQwD3T3Ac4zNCqyaYuYS8eKXheepkD//pEFu
FJ8djq+BpEjTf8+lK091YK7cjfWEifmGzP/X8pyRJGCjBAl6Z5wZuoeNJMATvob6
qp3FZnA5gnfRaGgWHELV9eyHe8sfs4IUFA8Bw2DhY8eanc1kft9vN+6wZkCGyFof
S0DFCzNPgXjIGtAXVOIBOM6kYrKnTtE3glUSI8Q4clfIc0wwqwI5UKrsZfxm9/pw
j9Baq35y6GcC+qm2drH5z0QXouJxVE6aZQRcyE538l9SHFLsbrc/rOwygCZF8Ykn
hbs+aWJHE5AruUKQXM9PWOYCNFbeicPC+oCFRz68FVB9mpcYOyH3XpiMIYSAgMck
nEkuDtRSZH7SXms7ritCQatxSoxnfACu9NAKGlYBG+i5/nB4ku1wLd9vLybtovsg
ahg4cXrmwmK3X5HIYqaJ4fbllY089lJy26C1+K1YlqxAkmp6IBffS8w7xIffNWVr
pL+jpucuBgGHyVmJwyfUpC/nUKnaMwKJlnnJP9QZDU8FC04hdBpKMjOgSF+a8a0E
ngJW76RfkOYJKBUoK1mZJocrmJHMOBJJhIDjArQu+5F0E2Mo6WvGBfgxHTQnhUnD
qMqCND4itUlOtLUj6816lC7qqsrghJcDSZOrurwfuiIciJxZQoH+iZiadM8PdGa0
HCK8gV3iPzbiGK29I4EMMVErhs2WGB52Hyfec/6pcHGPM+njNBFYj9vFqIafIKj9
f97kM7f9IfyrmoZ2lS6KcTKy2NUQsF1ApiXH1FEEnCd1FK1OepeBj7Sz4egpPTVI
/nIJd4+GUsa3CIhZGfWAdhwLVMxR4G/tmowVjoLdxnv/MpAGcGdIW83uodXpfuba
diiRTCpUFlo5flFMBdt+FfdHDZ28i8GwESuP23+kq6ga3QdE+nozbUrp4uKmQoPB
oK8avAJaYBS5m5El5zfRGS085vnWOp0U+BjxVBiIPrgznMNq9DUa3/e1qMxlIqQY
OFKyfPUQk8tPyhazbLZHxth42BXtWeFFvfz4IYr5cY58tQho8twyr7R0Y2Ce8pGx
e9HApIfa/nOKrmZssI1Zcj89aldkQ9NPw6aqJ9m6QeRuKsiPb8LwAM5089sulzWM
XtvezPqhdIAah3qGr+ATK0mZfzQ7DdzBG7HX6s3blupOoEZseU02OikVkNu0FqF0
wLDPOU0on0Hlsf8eECiFu5BCeCTkHtgmcWGrkHPIobx7NWZ+zDENav68o3XteVUw
BXCYmyApe8AmmRyKW41ViIKwhA++N47DqEH5pDhvLiIA+oiZnJJHFGFtZzYyH8L/
J6FpICyQDntdpiT4XxzfLm1GfLu5k8HnwQcmaNTsmLpcpe0G0YJr+YUGaFVg+QOA
IVdGtoOn4b4C/k5pcSW5KnENyXvNNGO84HbJxIVxVPeMcjcqb58M4hdoF4nDFNd5
3xgCoIYbk7RNji3hhMb3awryyVSRhH6xfxdU+2MJzBb9cgJlFafZUOZu+JS3fQaB
rTxfLHoAbFDaOsVHMK1mISUi/RbXthq2hDwS/ZqRpDuIRXRng35Wxd7lbF4pCmig
b3FUg4XOxC1kbAbHArnEb+pXrve15gKebKbqceR6o6HkoEh2NOTtX7zkEh6yeeJF
Xa5ORCKU24rABbQW8bv6HoVRoC0J44txQj/1F2OoUTUwiOVKyKdAT5AEXKaDpPN6
HkcqQoJrjRg3A0HwbkhZ06lCrPFwPCXKFvDoyihyvMwD5wD5Mmsr4mKBY5gJ6cKA
3Kgkb7cAJNDNaxUmR1+KbN5VmOtKFcK4c71crf/1xlsnNuTK6rxWW4FwF+sC58rG
A1IuctflzSwcyd07jkj0YBBofHsDtNK3K8bYVp64o2DWncwAl+r2Zkb/iGqnE9Zp
dl9KZm4rrdRVgx/lQxiFKG6UffjWIEVm3n06VwSc8F4qhg8ko/xJpJkAc6FrP4CI
gWdkcOE+ByBKOXBjDQwICmUe/eFNxzAZD9UGsG40vF8xgcKTxmNWHhIfg/GyAIl0
6xkX+5tcvM1Z86+InDGLP8PQBu7w1VExMDeyvHhR+xxRofNQ4ue5XVxIRrw52oWU
m7iIm/LsG1VlA+Ar0/ixDdeKkAYBwULlqtXMAvoQuUfR2ZsKP4HwoTxU+VPBrVdF
IpPDEotrDh5HPnaNBWDrOTKWoyEOteGJGBtuhGXbCM1mDnvB66jIChH+mZ7C1bfh
OcVcMiJSFjvnFKcsEkUbMgB5v+3MSEJiEMj3D4mKYAUz0M7io9bPp/purKlQsuoY
UngnoeXXw2eogB62C6wR4jfXObCtbHkhv+9Tt5ucSXkoXONuPnNJWal0CgRDgl2M
9eOylOeOoRcjn3AH09TypczhMIyVmF+Q8EN9wFroBTWELXVQqwFwM9NtRxAQgVhp
RoJJSqekbTcN6oczgNBF8t10tyOCAHdMHezxk8rpXZTNox1xnxoivgfoMGWAWP9y
qHZkLfaTrfjZbkIbjHn/z7pNv2c8t+44qxoeUmg8tTFCcyZVlYf8iZ3bJP8H/CMO
ptwXgqeWOSXfa8HeM0iQhYzbNmkqSpkQxt6qAlw4zrtGmTbWLkcbDNgFPC6unfv9
ZG0PPM/zYsTQrgRKQWbalfHGEQmt+z63c0cPkFV12q3uOlgktiEutqS2eMpTlsWG
woDPrcJjMEFK72MMFnimx0phxwp2xvScUeT+XBJ+y0v2fnh1sfhJ6nmOOIBLqBtk
PUQg8z0XLNbkCe7IXFyEcADTLcsygC9zOvSc4pwEtJUrpjQE2X5YebYdScJNo6Gv
WNyQqkhMdZJrIXdRY+EBAItbRooMadMVxUjmTPM+g8DMdhhgSphYIIPW6n+v/7Tp
iMdyf3g1KAWj4bd7qm9YKatglQaGNXv8VfvT4aGX2hN/DpiO5tJneK8CodBf5j7x
YzCqzDisCcoi/3pf4ykw/DBfUB7mKR46qZkvpFOxl//1bswgADdLpTBMg80oS950
zi8Kc+QT2PQ/VAEkfWjAn9TUZSdt5Dt3FgKpDGB6jCrUxnKFYybCzaUkVg5o0jz+
iGP5zJ/EBGb5nDNPvibnJoARxBx7tzXZsaDJpvauW6krxmvyh/4oU2lE/d97VAhU
RTv456CTl8WQru9cJ42DZi8aEOXLw1rCDw1Ec4er3udik95DCL+7a/tCFqa+QbF/
0gLtrgOp1a490+4u8cOsRFPItrOW0O7FB2OW9orDgCjRGHtwDvu3cUQau8Hbuniu
ZwG386VKdi+QtmojYq69NBwa/4hsLpJFrnLRW1ka3M7vcVC8ix9kLGXYoPU47gYe
IhI3PfIrUccA0zIMDXIneAQQiaLRAXIy9ffGj3XwtdPqvDpD86lnx/cl/VobCpKO
rsGDNnqKkVC/wbDNIkH6A7myaFtokvWC2lXdgz/8YelVcxak+W6jE/qTPPXmK/I5
hTXkL82ldKpO4vfYNlcObBNvGSCh3FQZt2T0TrDgie7SN0CS3/Ouq3903r4aOOAp
M7EecS3JDgBj2bIzBbmHeC+icejRl1RrYgwEwyiDjCn4e2RDvmKhjtDCkDiL99pq
+e8/xQNbOrDXAJkQ1kOckpr9sdf4cVjMaVZgHQH821nByyvUPiK/Rr4qoHcIabpy
9lqQHLb1GbZGENbl6FVDudd79ouPCqBWuK1zn8VnjbHiASugWCkatcPBqa/PAC3Q
t9rILDPGVlRncPFjq7C0MCiVFmhvV5i3YnIw2nH501hxIWITRAF9/7iYRJ4V4lKe
nCt6uIXHyJfHE5h74oQqg7sJJ+0nub2LPUfl04PmJ60mc7EhswfGNqdjc7Qs0Wy7
Hy1M3PNw/KQU+QADm3K8pb7yHbSHO885L/y+8Hjb6Ubf2Y5fThKozrLw6J6AlqeR
aV75kDWi31MbX45G5vZMG2LmPC2Ah3LWS5f51+oOQ1+ZeCadfV6Ji6FRdaFmAuz9
tNNhOSrpFADhnuPA+kZIpiaur0+c+5Jf0GUGHfctzeP8mkuiR/OWkmzTl3mRLwO/
u6+tZK/kptNpRC43t++BMmmQGlFvC1iXZzZ5bI63NEHp2Iosk7Mh0JI3KYXj/c0T
wJ+0buaNpPJvSsjlL4Hv85lvH0tqzkMxT7U28gFq5cqU7SBVOhg/JxF6zWvqyfDM
5dItrUyr2F7f4yxqB+aezlbzHsdjAEDV9wspimKPfL0hN0ju4VMRUGi4AXcjq916
iHOa9ww5Ti03AeiOJdBiItjXx+y3VMcFzeCWttRJpV5p1De+L6VnGbyffe3qzPwR
SExPCE7XdrItz3LuuyemvkotstZbqN1QTqM7A/RqKLoOu6XOSgifiz01RP+Jjvoq
GQzZC+XIJMBwVEKnzKfO7EGw0MaKd2txIYRr5Dt69Sjo7/yR+82qCeT51tb1e8YX
OVq/EUGyVVRMAZm+t8a5G5Fzy+yYnMkO/AfQWx2iuiz885Pw1sEX6Xi9X7WgShUr
iuhwy2Dq+YsKWjuFlOgDBRQg1IDap2v0gKyygF+KWH9L2UIYcbG5TMhAiun9HxhG
Q6KOpoR2Dp/4VUIGCSY97GL4P+NWmK0kWSNU29JqPCBV3scm0AYas9QSS22XoFVM
XRjhfdLzIueykV1oRFxwEqWFuWoKtMIeRhATCTSr4jvuQSyRn5MC3y5jRw8hQnED
WOe1oolxqHgUjt/zSeCigG/0Qzh6w+Gde+p+T4nScijdzxKR5/SjJpGZdD1mKrI4
gLX1khyGU4aM6ZibgTTZC+yRntjvEOzJRY+1SjUkKnKY2K+ClPLvLfSAaYC2yVoL
SllZ7qfyXBQlY8S+XbZIoP7jr1Zwubu4g4/DV4gbe+pRSSzRx3hq9FZaT/lt0c91
u+m/dCm5k+lxYZHqLg0r1qVzLEY0Bz/dc/9/EkqBJ7PwlOCoRIs1n5lsStwVsonC
F5i8Oxvf4LDRdWN+r+RSaVqDp1OcdhRcTouYEASB+jkSME2W8v5hwyXzWkjJOMej
+L4luDgg7+2D3cRHToPfUAVii4M90zQpWo8idbg1a63uq7LvoTsCFor6WbuW98it
oylj7Hovfr5eRHcCb9STmPaWUAucu55TYpsCZWs/X1gsZtQN6BFK2J2N7HY8kUnX
ZHqEhfO6+j2C7j4+qTl70OStuK49pS2UPcqWR1J8ccpYIXD90EZoncwI32zVGOro
6lQDOFO4JbadjcYqBqbAy9CQ4zunkN/hulgl0bptBdvXC0gqNr/mGPwyFVFfKIfv
H3EZesN6BBX+hvAlyM/xl0ddZCi+KXwVJKs7C8Ap0xRARjGI/4chsp79mjpwHera
CjjKLf7tr0MJzGAzeQfxtTWZ1u9d/Zo88e/fAZxiXALaZpu1E1Vh0fpI8qvfgeLH
oDDt7VeIYxJfcU6lylGANSvrwhBWUnqqDZkgrNDxva8ukJpXx3FAuzUQIfII4+MM
dZgBYIK6OO0Mh9fxL6kYjHnwm2FJGcb8Xtra53/LrkRXcNCfoJujYbciDldZ+2U2
67th3mSnx2uavRXofZL3krez8Ylm9zHuOhpkjENvR7vjrbPS7NNfPUdji9Li8Y83
j/0rVczaqZt5QpxuWuPwyoPG4MLIx+ZjhCf1/GzqnKHCDZyKWIviWXnlPiH1GLJH
BPAuzFriBLHEyO78nIBm/t4kbHu++3Grd/B/aTEzt6gRDsWKs1Q7PLzl1a6evpu5
YBYaz2srX+xXEaXXvn/+exxeV2ZXfJampLrRRiABY60iaxkU3wwnbolOiAsGg+MW
Lytvr9v+dhkGhQpnSUQhpUkWOQ9119DrBuCMaF0k411oUkky70InlybhHW8THVFU
H0pnewQ1Q5kknHWP+nQBmKr6BkCWPmh49KHgUVDeTUN2lqN92fl1SB3KbUKnciG9
9xhM4NHPjqc4PpB7eFLBbNvc2RoVBZkrWpnAk8NYOQKqzW4LXN6EbOr49hXejaoQ
xAnuffeCXlfGOeQgHsN2V/xEsXY9BP2pycdzdIM9uQtm0YriYUUi1m2XPicyNqE1
TVtOjg8gXrHTSRS8PZ9y61ltOGz9sy639WQUH3jeRdt/VG78u5zm19xVQbuaqQQ4
HGGg7MfXPMFe4CbwwrweQZkXPYcAX07HcKdUVXVOerKy5lsyJd7AFMRu7Z1sfu5I
HSbTsk/531cnVoTYwTWSHfOKfLdGBiVAIK545njmPa45xDQADhjvgUdgWpGkYl+1
OHRhTOd8c8cDgNH36pL7KT+dS0RrG5Wa9MQZKdAUreyIsGzsi9g6yE/32R2tbZwH
pnoB6tXarCvmwmR5mGGKNzARhIx1/BfihWZa2lYZrvIY21lDwnP99X26Mjg3bbsk
itXSO+EjPD0yp/2/OOwBlpBi3RB6K0YwKzPmbNN00ejMJ3L4QyeTjW9IwdndP0fJ
AGF95qGGTyOXVOAbTYPxSPuVw8utoSls+6mJLWG8r+DbR5C1xAcC2HHdmAnwowlf
eU+VJTE1T4RKA8ItDclZC2eobRyZDgTtyxIjcs6fp+xaYicGMW1PGggQiKWgbZC+
yeA0zBfm44w3S8IRNyQbAy3B75+mi0QVYuPRiXWHtX547/L+xzDYwwQe/Vltv7VN
FY9yIhLdWmwCurex3e54Dc9jNYV8gSHwIjeKpsYJUMeIv2h0ZbdhB3Q366YerlZZ
tGArM3MI2Be90kaWGY1xbRyow71feFabL79G2LA+aNJEIlbQGE3UOHtSKHQ7LDz+
C1MCO3nEMtHg4JV27hR2RchuEibZK0JvukmZr1VmyZks6PK5e1Fmkq5lMO5ShL7m
Jz/HO13zR5NtmNgueJCJJT6Pl6YbLInLbqKOAInEKMNmTbr3kZjUFUiRzB3g1VaB
iFrSSegpBrCVbux2e0J6tIsHTH+3rQ6q2zOeYymhOoNTJx4iedrWkNVes0Q92uM3
4noa/GcduO+MZmGO9aiSMBfLyV8y+SpKC1HN+JVJlUw6tnECHDeyjD+Rku81X6qu
NtvT7MV78pUVKLIAB/41PP+D2HBZEsnxYztgw11Z0THEAL5KkAyDT7qfhYydrUjY
cHnYUeMGD0iwjqN/l3YcV6G1arCpt/ag8JYNXQJaQirA3dfryBL5kL26o7dnDKAg
O/SnvFVxISUv/WzDWsna3ozg3uxHs3x5QEdst8jTCfVlWFL4qnKNe75V99vXjOcg
Q8Bwf/NQbpB27CzKS6muTW195I2tYvAbkWiU9ziljSZM4shLRsSd9KDDehoSS/Gl
THLhFrwNlh7d/39KzSX8NCXdv/QmVVeh8Twgz8p9SQRmPNlq5Xf1OX5U93TUs4em
rmSSv5aWAL2n3OYtgMN3UPPg/5YYbfTO83T5UEouE6o/gSRT5+KoGnk+21GL2Kyz
3lMU5wirShh+MjpBg2IYea22H0nEDiTYnkjUPpmoJptXCvqMPMnm9PlVfUKUpGVt
JVZRbfE5GnpjUELr/qBIDirFpE8K7H/TvPmxht43OXT8MnMnaEoyy0CkvAVfM7Li
X5TY910rVWvuzPiMzybYPhwUkNcFZ93D6IWTKFFgdM+JLije5s7Ee8hCGMeUwLyN
iC462bRzP8+EVwC/KllQ7zR+5XjSsr1TMEIKje/ybZ1GuIo0N2Nz74I4/Q+aP/bc
TzYuQouuZmU+G9AzgImyvkr7GwnHS9wIzmOcL4ZzLxLPk/YQk6mo0/BZ0JVPwN+u
GQOHbFozkK2A0s9BQpqb7Lz4Fh3znpxQb1cuqzISnfSCOr+gbM5wqrf8UQm2xSkO
/U+V9Mxnh92IPWkRpi+l3EbEzH7zCf4x3K5sYchjFqgXAzFxQcB2UgQrmUtdOVUO
hN6IJBA6fL6CqNAZKe3x89HUNi1ApZjmZQ5eGVKjOTh2PMZ/G8HCB/7HY+ksq9gh
kRbs2m22ep6Ox8rDcUVvLQTjFLzFkNBDQZBCcYU2JYSHEjVTfIQTwfWuWOM1fl8p
Y+lm3BgHxMKDI6C3K7v0yR4nj9Cd+R+0JqBBjSNUcquv7ua9I1rBzCiQVT2mj8sG
1Z6FYu5N3mMRni05BLJBigJpKgiWP9ZFRQBIJ+tk4AUhPpXkhFhC6yw2ucw0XkFr
ndx/Wn+DEWCswCJ3YARqkyJwrQf2lf9gpt2gw1fpcmX50yyBLO2cAtB6Y9V66qBB
ZrtmqlJE5Jwj1gufKag2vPkeO/7bMuGA/U9Xf8GF23XdWd/O7zv+IEu257bTTLm0
EqG4Zb4S87RP7bkv3fqxeIKMmvoJt6NIVWJpXsE7sVeuK8khaqQbJ9V5eEtnZAqC
ydazzfLJarfczo74RHT6VHc4vRJLg5I3bpxF3wblxoMQEvF1fz/IQei/c5Emwp+4
e1a/3NvvMBPlYjRKI4JzpmtsXoybcur28RXI8n4wOgls4MP/55tjlPRJBEZVgyRd
zLFVwgZZaBBwNsip05tTwdaFFGuB7HPeTfD+Z7lVlZbnrCXsgLWRhRnrXeXbxZ8w
YH0Io8od200qMdKVFjBwJmuFWBU0DCt//psKBAk27KGOuQjLvmEZi7bqLu/Ni+0X
Mtf0qt1LoGU+q9NJfydrst2MbFoq+aiNqxNSSkw30ClxJzv3mLopHVaPI3ikrVdL
htEAzKdgbw2V5v3atpyy+16TXYu7aHA1lv71joZO4yh8RzeGEzeYswg9YegJiM9X
3X+3Jz6yy+h/7uNiqf7I/SJeKPoa/qjNbA4mokJh4wNQqM4gWQ23An+e24d6qS+P
ydvmIjxA6byuGKJwh19kPMgHXwrJpZpJmtWjeDgfocLACfufI5rEYSzgQPTmzuFh
kWYO8eJiLwKOTvMHzE4NVSLGsMYWZNleFEtxN+CllbeiT2R5wmq38WXDTSrtTwNj
C9KL6/Hi9CMTcihDWgEOS2sbw00Q9nd+pPJQcuzT6FAcuTzcGAq8vcDlMKBF4UHc
xKzJyk73G1K+06wgJPQHH6+5QvUqUU6t53jCv+ZjbdHTqHwv3N6tJQPYReNwHvaa
mTlzxhUrAVY3lgwFpYQKLuoXqdnu7LtJjNnyfEEXdwDpgjAmqHOw6PpcN0w5q59O
buT7I4FuDeUrl20B/ykA2mTSs9CulTNjRysD490Ua27EdxK7gHFC0KcXehNlVtnM
7WVcnfV4mf6xDwzIhffGTOUaqSeubknCOIcf6d6Xnxo0xgfqZB/6dBfNDng7nRjw
qABfTjhwSGPKmn4MaWmvP+umgA6bCCXk1W/QiHzze7Oo0wQRqUGwtV3CKXgOZAQD
7IlWPD4VHCtt9d6b6M3XLWBZBwBnB3ZBf6rkEKhDaDP0veYVmZV9NXPxdy4ttScL
56VnkS5XeBwhzWAE+HI8pi1NKEeDwJzKXj3outwpjyptHnkn2d7M2zvQ9INXF6Wm
B09VwIPGV4tyJdiFLwPINo0OMetfyHUJPt8j4tGALKpVbPiu73bCXUrjqTzJdqQf
ySvsz0cuTo1h17xdiFvGGH3h5Iu8wwRpeO6w5TYVrQf/pB4+kuTSPwEYPt5kL3du
4E7f86RPnK/hkmxKatGmFJM05i4glkAAB4fBvReq6rK6UbHEM2Tm0i19NiX+774n
YXNn5Q38xpCInw5u9Wk86LFY1Tbycp31K31MuDtio3DzGbo4r0z/Dp4CDA8UgNrf
WpKTghwpfvCu//0JFS14arAFj9ID8ZRBo5FmQFk1RKVz2pHtGS3mRc5w2dkYdPxd
wu5M4N854GzCWSxkVZfZb/qIUlqAicR6Pjv72gYAIXTni88FGDQQczjikhivVrpA
YWTy1mv1ACS3UYIRQnhI5+Wxb46rgVXCFodP59Ze3CrR4taJzFNBDfAng09jLDtH
FnD7corsFIaFyAQK1RtFcHz1H757kI96QElxNZ86ZS6z7m55FTo5dAgqxh3H15Bs
VIuM+pvRJnngaoB7xC4eLtvxrxAGLE2sAMdfInCTPMoklL/fngcgBUxOrdXfSRNH
Y8/hvZpKwmqPPGF4fVVo570gdG9zsnr4w4N50ZvJZJDn0ajIaUQrgw/31EDXf4RP
enRsqDm8oJcrhPJuLMtf9bttLtXDfuHSRUxvYeyDmG9A1f9tivwwlM4ih3AwfBnu
5G7R3p+Oa0cLGqdi/iwtbWQo39h9YnPrngoEbIUx5uK0uGetitlD/MrbIpE6RtBd
N7QMY1kjpAy4r29vZFsRsE/UmbSesT1+/ykX8UMdbDdYg+4bOtbXexhCUKBezYt1
dm2mkB3SqafPhn/6m7SVLNzE/LsAXXMmIyIeH2b17M1x0GdoRUs/rYWA+lNPq6hg
/fHaEUGgKVwPYVU3fs5z+TMt2+nE+08idgjXdIToS1SVjRyh7NWPQKMhDEsGnQRD
WK3alJDl9VNcmLPuHgeSxoFg3MEasAaU8Kcr9JXEdWXpudH1W+JxF8tAFM6T22f6
a8puJN7HPDM6n5jyNh3Az6Z79EvBymeZXvakRBz9YCtg+2GJ+Q+Q4hA/MxV19fpO
eDlpByWw5TzZ9zgJxrklp5zmsBZFrgj1nWdUjUmjKsuZoVI+KYMFzqPe1zcX3ojT
T25+JzMxMgfU6hfvT1vvySNdhnKngX+XdeLDILSuxyPgpMrqdov2qyPQtMCdxv0r
YP09Zje/Yljz7YeH4ARHJX3xZ24Kw0YrmktNqvjUv/CLDf3JRdZ6yn9frUs4/Hf3
qkEJIzwXma6YKt0WFX5c2rcrcEhm8wLc4JR4ammukwxS+4lKQ61vex+MYTXLcDeX
HB6hF8p9KjYUAlZbqTd/SqoICKrv5iM/xfUA2qin2JPZFTszTdYDIuVE0nFiJY16
hiBSMmBobQwGXJQ5JaeK0MNFtEVsv+uvOX9tuaW4K2ZnyZYDkv8CkDfoHqAWgLT1
ErPfriC2KPnCW/8mB1SkzU1knujJMQradKdEQhZ5VN813W64+NWPmepu9fMZ9dhv
vDc3IZRRnIhbpT791rCyhwqGwhgV6xgpPhDpWboMrZ/+TyxD+5JaP27ZcstUCZAF
YPL4JKKx9e4IIQdfXrUz5Qn95LqLnhEsP/SJWgRvjM+O2le72xYXQ8qNGAexiuCU
iwcvnXoZEV9RaQ67DUX7OKJ6l5LZg/17aFquWyec1XdOr1J7ocfEwGQACuWXrz6I
4TRmeRWHQWCB+Rr+OAqpAWBurpgzhJ/ud7Ym+7qrZlnOkL/wusMcLWMq0Ohmd1Re
tVafx9uAZlBZyyP4C2n/ZeyzW1j0RIqIHQa6eg6ZEDZB3/vHJRM5tsxG+BhFLXfb
ASMfW7dvzocKCunT7wUtTNSv9NT/U8NreO5ugOsW1gkX9jmjGPPkWVnhdVgDvyOc
f6rLFRFyylydXiTG26Pkf4PKO5AYU+0+EqfDke3uQ1ShRcYFp3oV1sSC/044NRlV
phA7aDMgvWoZuT8eY8uSkCtUj/SiDBP5zzL79l2k4ICN8sfI+AjiRI2dDptC1DnS
F5Srecxg+JKGyadeiBKMgfhMOyUwLoFnsG6P3FqFFyufTPDBUaGYbeXA1tmyctIw
h6UTclCVN3WD5lSefU9GpJIqLcPu/3+/aIF0UXk3cpJJSCJk7hmcHNYDJkT9AVaD
ThOxBsnqIgtJvqZI81VflutL284nk6NN0JGuFEeXjmhhgfpJMuNMKC42ASmFVkML
3RHCl3XJ5LZpFV/wNLu8KToMddCicbbR+CsFhmdwfsH3N0PQmzOJqoB5aymkfUCb
DiVB1k+amGZcOXDMwo40Wd16p/Xv3IoXdorbTPzqwfUPweI7Y1wGbYoKvFKMtXHr
UT75fP7GPUiiWMvZCPxWA6PgAORGMyeS5TeRRL+JiBgZweX49jIeeHMskCD2ERUX
DGQtda+glA3JmPJh8ok84mvGIvGVtvFq86ctU2AXg/2FrCPXy2v/t1IO8U+X8PN8
xi14iE1yMbFR6a23jFmTY1cA9wIK8UtKGmB1Ci5GfuRLIaruU0qrJway6Ez5j4sy
zNsxq9dvr65H/xk7UK9Nov8rYGyFm1LwJ5jJIC3EzHGNIOOiw01NMDpHmFoVgxvB
Z62OuE2NnBo0PKQRmZVhHxm4t6TAicfVryj90Hq9GCgJm/BYIPPRdr5fp/m6RVH9
9uNXpyCKx/hqxpPOMDKODN5ynOlnPZxmH57wXrn6Z3/y3wzTxx+yt4D3UQ50BmOJ
IMu3NuzHr5gocnI3moP1BwKT1r8XFXxl0mhF761PgSQzOMIcj8G5+GjKu9vMvSsa
79oquXec/PKdkaGSK3db6gdf/DqfNRXegbBBqQ4t1VrMThlU2NHsK+cKY/7BYLGF
hHyECGJ0GeUjnKMJNrmb36CTlM+dp/BggIitBj27DSFtY7PSOOS+XSBWfqy5K7KT
B5YMa+xZb/mW2U5OwSDpkAX93AiPGGilUkLUBWhkv6LJhGeNYHhCSwVIYU9PnZwQ
a+I2UeScEdKs4ca66tahnbhrc0sLGrA4+w+AlZn6tKM/Nww0kbkoZMz6zP3pqYRg
gL2Rccjx5lCJsFFGuPnFfci+SL/brgV0XGTNIGkyEqtbmym6SixBMsFssKAj+/H7
EgZ8B9IfWechNt0bMdfcVm2bisFqbXzE+OPPTSz1DmBj02CXHyg22rBxwuiWKWzn
dzq18yBN221n0KvysMfv6Xyd4pEEEoEJYph+Rl8bPFgzFTH0BYCz5SbOm9UBZDdD
Fi3e1EaWpuL/oKHknt06nIPoy/qao2VLqOVc/PiwgfvKw+FoPdoQQe2/cEdL7t7Y
SjPOvYJPa48KWNbrjRiV/VTKDitMYML5TTk71wcThEE0QA/bUm03IxlfP9KcCOcl
QD9iQwgZ7edqgFtjr84/1aRSgkWcCkawYuqKXweAy14xjvkj57HQovNkiNbYEM5n
x504ztnclgM10tGb24K82AyEAEI8a3eHM5sAnSwIsAlNOlCtFpX44vj8MiJrtlOP
E1dskKoCXzZXUnmyxpQvo8+0TQxiS0kwoF9A22si9G2kn2LQuM0vi1wI/SKb93OH
iOwS+ludPu8ex40helPR5mPDGN2mNOk5YIraVhxZJjdR8AJaiGl4IDQzNqzUGQ6h
+L7e/0l8F9L4ff4Klt+XbUo+DeV0vBaKNWvzUUurgotoWicbR6qmvY2URMnT5NyK
MaQCq1QBd/0KK+T5zIpa8PyTHo3iB+3WkSGbILJ7mBSbc3p2TfOHDb5+dqKvW8m0
J35QZeZ9EU+IqgK839xAID3SoHzwPLibnQhPfD0v0ZkEoRWzGAUHQaoIGlAULYb7
512onc/l0T2+XErKpUMBVpxvbuJpU+RWKohWQHhNXaDeU1MAJVD+pBd4bNkNKXt5
smqWv+VvRu76+SmDeYIdSJhSmgNLNln9Rx0glYePtNMxUQNDqmvMDneSPZ8gNLZO
0Ow4e+Gh6zEuSUkAMWjOOrVfxCdT7ESQVZfdLtVLl5nMCmKzLvitbuTBjJ2j20PI
6P/Be3wZbmBRdbolU6bRIOD6/HEuCG7p4SNNs5/u0S9GmE9tVDBbUzTSZiri1nhY
t9eHyfMfl82sAbg//QegBREIIJoHrNSy5zj0qaycRpwWwsWQZZdMqSJ+kSOhzig5
2d08eBjHSDLF+CB8nCDjZGFMg+Td3GTWSV+h8inTfdINArWuoIWhZgBSge+vhBIY
8z8sXyiJ/ob4pDLtTF6xJrvGUSilGiPdPu48bojaO2xBkcnpc/lLZ/NmZlY5JrTX
eqW8BEoITw3vMPmq7XH0rsWptpzjYNh2dnF7mHMRXZiPvjUlpAJMq5f6OOO5lbuV
KzvsEY1P5jO//jmCduNZRCPmF67OgqDyts7IQOABHactQa/+UM5LN37z2AGI7wWU
WcKeOkAxq0d8+qgtZ9YhRdg1V2K2XSA8gS1atOqlglTrjh/3j6yeJ2tzegYCwuR0
D+2UApU5dOl2VGzkndF6JfKhUk43CHg7ad2dBQBxtPmDqPncvvGV9XBc9JrD9fGn
KOlmJI3/6sPO6h0zmf1wDmnFa+n6Sor88IJNnYpY9LbPam/A/Az3OCrC5BS5/LPm
SIbxoZekb/WdL0Xfoi6GAhPvZByES6BxbKYs5g6KCINX1oTDOrMAGB4cAO63Up0G
9WSec/QmXhraRHBdKIZDtZv3225rbmi8+OjZD5jTUTp/25sOKvaHlR3WmJmc660/
zVV0vQMDAlTh5uvpWpFnNuc0GsrHJVxXoBtIj1yjm8xp8PjO1+Vqy7UmXKbEuBE7
QewPHc8Nb26LjHfu7+c+sQGXBvfUmyRZSiEB3YBlSBDLA3aQBDDvcblM7iB78euC
sbOurDXKQoV4oFtGuJNaPOV2LSU5TE/+Y6204HYB3kceGu/9Tv1awvZUWj5aeWYV
nca46TAPS6XE5JwgxtsPVmnYWP8DlapRZkXXOLjAcI3v5DiJ4Hq9CPnXeZvt7Ayh
gZ4uR3n+ETzju9gIne5QOdXc8G6nSF3KEfbNQnK6Oh8joPkUvfzwjxO/Z/rWb/ZZ
gVtpyDdgOERrd+4/TrkqOJ3AyfQzJUmrnUyt6l3IneNPZCM/EsOg6V+R00cRgqnF
rRS9JzE67eJkIcB/Dbf3AjaDDppMNaVNP6YCXfUdUjsA9idNwQHPBr98RK0vXydj
6LmBxImpg4Cho1QjPU8GkCQFbGuybf0rRLirrhuXs6xUsErBdyPPIua2td7Ynhaw
YW8ZYrB6xl1JrAUPrauU+CCMnyHE1XK4UEpsfuf3ZLRO3zjtnVT6aj5GcCXp8FEn
UMratCwXTiysDv4ME3TWKZRii1nN+t/2fPszYQxNl0vY1CbVfl+FC1VEhU7oOpWL
T1wha7lbMGIInJUw620T5CqVfuH6ouoZORa+vsCE3jsQEQDrTPv4+/gEtfRFekIJ
LxYCGLl9wA/OFQI7sMcjPn9S1oiDIm7lS8jTdtjol+snxWMWORV07yTVxqMfRoX6
gWj3Znty8ad+e7uB9vAsUrHFyPrgUamyR51Zp1ORruzPrr78RJ38z26JAoqYnkgh
njI5mJ0YRKRTkMzEQwNcgp+NotTpT5oh4a1JVKZxBumLc0LxgNtSVcgpDE6iFvIy
v7R8Tr7RxyP97VOta0lI1ifC3L4URnbSeI04hiN6CJTNSZtbTtcpKJ4VMAGoJORW
Z/StqxEy6OLnNetmwVqws/MZE5yC5ZbfOzcfsL2iFPuwzu+7zMRVAr2mNzx6cfd/
JbYr4UeaMeUz3kBMioscqaclD7/EGisFtksh7AtmdcOPcb/OKGPtxMS2EjqK7Jzx
zQgaYv/RNVAUZ968LmXnLoGMrlhrK0/4QQq3HTwYBEO1RcRJ+bo7GDr8AVuYnhjL
h40Qm4WVLTgKtRyHUxpd2jLO0am+8PsM1E1Kl/xq5X/rsPFI1LAN6LjyhzJWTvM+
7Fs/PoZDbgrxd3iI25hDciixEGLJkhBrGsTPcllY1AyOik9ajUqBaSDpLp29UoKN
WoUBFtIcUOAqJVAo9jyKDayEwN8RVWWkNk6iHNWb2tXhYYDhB0s+/+YQxqIjs/xY
W19KXCOeBTTqWqJUng1OAbWdc3RjdV2G7fAa8Scc1iiA/I7ZOwh7aphv+vyG/PdY
X34JFWFbE3CXYbezmTb5+NICn7qhnpiyb7Xx9H1Fqg/kQVz83hZx91Igi23QiUWv
wBYJqOlaCoz5zBPhzPiru4lvsSa6a7Hbub8JLF32rzCYOita6VquaKwASiKioRi6
tQkfejHLgYY8BhdJhyHaTxB7aNK/3OjLiB7wjRj7I1486chZrLoe1sN1R6R0jt1k
BLAJnaHPcPBth2WtRLJy6PcwsgrU2XBPmXmkln6TL3CbFyhDVV9GSCRY7PPvnrz/
0nlc9WEl1XruON4if+fQdebikG1efDZlGLuuGOeNE2OQUSlUpE5DQa6zIgvTXlN2
P8xR+7Du28ZU0q2H87vQUyd9Iu5oxhEzfWSY1GofV+PBeoBgN6zmUJGCnIOWG3kv
eI4eGMG43bW9xxr1wSHrjBS6BXANtEgbKvxD3ckmCOeVkD1tsDM6Sjc4Y7lcvmLX
HlUW0FvbW5O1CjHvI5kGvCQmRe5ja3ZWtP1mC1F4xhb/L3mi+r3wn9Mw1dtngdH0
UJzghxqJbJPnYYbbj1CeiAXp5w1E5ObpkbqRVx7NwDMA4FwoPdiKGhUYs5EJLU4a
gKfIj+/QGLL3VvuX4FGIkVoygBaYIVgzcaDBIKU6I7n9mw3r1h127r6DYMxHVTIT
GvRtUNLzH0JVIKu2PpLhG3c82RQ8X6mJacvXJezvp93yRUy6N9QDJLswCKOcaUc4
iMnr/lWM6VlPYUyq8fPQNYG586LZe3YEeiHkDg/bNhTLDobmfTbu93f5Wvr/F+cH
WOk61GRgD+4feEh+NIr2lz2b2DrFLL9JjyxjbdaB+bqHYgoi03TlZu472Oumen3m
exUy0mVAWOrZCJ42EQ2UjuFtcjZqKn1mrRMyDdX7bWYBx9Kr4DlNbF1Ed8U9ywIX
U/HH0r8yrX761xrNwJ7jAulCikMpGRZ1nKMqMQldxEvALePmVjD3o7X9F7Ex6zlf
YwCkPR8GFPuSCPXisKWp7Pi4knd+oHXX2aPepQWd3F36DWdYQxK2tYhs1hZqv9zX
9sGu4I/BfFf3Kx0sieIxYnQZyDOoBtUrWOzguRS7hccQjsZX3eKmacUvr3u+alwh
YewU88SNv5VCY7jXk/AB7M+qf4nLXzrJJqGV64kHBrufzn/3/hXEiHKZtcJn3f6T
p2FAANMJgNh6FkDk/QySFx2Lu4O/wLkjgdtWKle8nu+ILJAf6s3x2S8Qd17E/ipc
SD04co0biFIN67tWco4JHj/S/UHDTmBUib43yBzIUSPztZL6AyYS/05yNgwMStZh
5VbqGOLV8iIp0fKM8N3yhjERn1jiPnGd7vPHylk6RvN9vwFjfXKANdU5LcuxEUg5
w43arhz4lS1/G8zInSl2reEEMGCSbXYmJfMCb+0K+m7zKHbONrWjsxmrbGJ8gPgu
Fdj1EXWe1+E8e1Eckq/phlmNO3+I26cktwgm3tb4f98SoQ9EK66peJfuAExC8awA
RckJ2v5FwnpNj6S5eyPryaKvuL6wGdZIigpKV0wSHfEA6QsM5pAa6gg6OQ8bl2KA
FStWxRTg4gxu+yW0/D8NcW5GGXnOJ4qRIGMO67oxu+p0Oz1zhvLoH2Oi1P4w7VWk
fN1PEVFei+eP/JN1mB+qJ6J94gV/xxdFpjDokaSicqV39bjz6mCqU0YZdl9vH2eq
1PsVf1C5uwrZYxCr1KAqqzuUq/TO/GTygosksykTzF2Cz6QJNYkCjnzSWbGFZPem
usmoylDO122L7aMGF1AnBmpzSmcTWiiqWbFuUZQN70Ja/5dpaI4GbxkQS2Qq44Jd
mDYJ0lWcMegZ1BRF74dpcRCllA1Ltj/ZqRHPGiKbYaJRuW9OAz/XUQR8SWJqJNTe
mmNnau7X4sDQV42Hycxl9frJ75hoO6EuWOQFfaZ1lnPdjAccDDhol460aomuv1GH
BGYXi4w98otbgsLGb4aD36sfaGPOx/Q9cZmhm5uez/U771fK0poTGnli05hzHdjC
qUcVc/5Y+fGxait+4/rddKxSxds0zMDpKymUMMra1NGPa24dSxU2hV35j8otBUrr
vH0V5rQSLIAyj8JGBhl5hwNzIniD4f/bI/zVH+eWzVT+Tfyo/cFMv9seo9KMf03i
d0UbTxESg0FRpFMHt1SAT56LEweZO+L5GRiRxOZr1bf+nr6RYfjrea0TTKNWZl8X
Z+hCpu7utqO0i3AmvJMHjsgoBHWqwXPcm74cxcmo53NQulvQ+E8V04Z6fJLVG6rE
GqJViLHph5u1a416nVHfgUXYaIA2Aobv5NqI1WQsYNzz2/xzmi0BPvI/ebm65ijM
uu8DRC+1t4jo72BNBxcf5YNaP6A3i9nvR3QtRdkdgOqlemS/HmWDJAoQ35wKadUn
nao4szDBAFfK9zesYOz4EHgf5cmXPpcxUQuduyUENeQ7/J1qhk49cgAK2PrAsI4Q
BAC3eHMNupNOBM3/CDXL5rBijEd5POKmmbGguva3GMKX6oxDeMpetRcOtZPo+w28
5KEu4QpJW+1OGj6sexBuiELO5yiD4+zZCmBKXIY5P3xX5U63s46bTfJ9beqxqKv7
nTdqaO/+s8mmYEm7O3Q/owW+kSWqiv2ZqZxbcauDlihByvHVI5P9mc9DE6Ph+RNJ
iPJarCvAgZUucquaiRlvx+qKztT2GTu/+TKzEdsNeTTxmJ/tGub3eBKLvM/II5Tc
MsCt4kYpTVuKlxvKUEUPMHhs8torMWxw2bdJbDsj8OPL63jVzwGpLAyU0mXh5YTB
gKlfTibGzjPfU0bWbRjOeWegx+105sR3D3BiHvY0D7DJ2AAbbXQrlmXo7nRKfAVc
dbVeFh5llfWNON5HnpdBWXOVIfAONZqPjA6/RWQXpnOMvG1iFlb5MTMxi/MvbFNy
FQHoYplXCfP2vVnIbavQ7HMars8PqR8I+PiksTCkP3jIXnGGHlrxmAwcWsV6PH7B
bgoYpSulY7kzYgeUFBpGCczNxFwGVclx69VfLaB/BsaUbWXkXnvhZoCBBuVuop4b
/PwZH6IoMNrR5++h54uPn9GGDzF/SahSGsO6cnmMsyDSecPKGoLIal+hZEhZj9yD
MEj+CEz73HGbwP6YmT5PAyLARR86XEZjihx0Kvka3KC+pcHD95Oz7t/O3bmBnDL6
MBWnSK3bVKK80bBnu98juMxATj/ilyfNmsMKXXlK4wEujy32WVyVkIhRaaV3bv+o
veJAzSghLZoelGbkxgHQoz05WoST7b4hQK9+jInMXSFAFDQH07EBPZmCk3owe/N7
5fuCZEtGtVuwna8cZRPc4YGM0KkBAuE6eDpD7nR7vyJZ0bSzqte1Hyi5UtPlJiP7
TkV1e0kl0AhTFGRPn/nM5xKfKD9Ohgr8icfGGGm5H2WCKi2//ghMPFoEgLqqdBxt
TCD9WcExhHf1foA6FmYWkC7MiBHX+uZhkaJbKF0JBRBZMScnozkdGnqCHzrtadUb
xypDGVFLTGI3y07fCfxsp/eGoYDpoVVBrM5z+898ZEax1o+JTM+RjK5j5O5dKlM2
YOVln0KmXnRArpeRJNdWhq+IcrpI7arGX2wbCsMJcGnWQiOE4qulZYfjopQeFW/F
RUCsd9hrnDNTf0KlWqkCe4PRIsaBGESS3dC63yCMaHbRq+ErK4XZG5GYl6chm+7v
xrOrpJQvwoQXWgyBwQ//BKoMF4x6AA9MmZPImQbMXGx4sKbgo503gSTgwnj6TAXR
HDAJ5hJFERj3+kh2E5GqQUB24o8xGC0Zx+VkC+DrFqxpEQv6bXRDCOscvC4xD+Xg
/6o2D8cIRPVOq3S9J2yRRxe2unz3xF5GBCXWnmc93kRXM2CJ0DCKRwEq/ez85phy
deSjVfm2bb0GAthBKbBHzWZwMaN4Qd1gHDlV6wiGwstWNkN2q48fBwhDbu9lRy+M
8GDr4apCDtsFe4UEE2j+wxToLwNd3L6qntgOLS8LfnKHti3nnzv7+yUMnXA6lEb7
k5E9tnREoHlyQkZC7ebH8ttG1ZzX0iOlmytbROHlh8yLSQAr61LX3/ymnzqmoGlb
uaRLAnxzS/ZOXELIfS5x6ZxALq2j2sQuxEBcPJvPyII+IJIPP4ciF7mO/tRqoqea
Pdb+5/TOQVo/9VRxvu6gm8uzo++RvDoxXHQuChmPvvIFu4vxBSoUxCcjZM+WyAFl
q0A8NVcqRf/oSNBOlfFbvIa3t8rpdXiaMT//gqfrvC1U84BiVwY0nRvfE31f/BY0
9dMBXvuXtj5qDdcZBGM2viizYLR8sX+RkQSARkyHFhREYXKPILDkDJpSNHva05NC
tohqp33KUpWkE8Emj5EsfIyaWXkxIv1x/0OHzsxOUz1fb7nHCbJmDhacdtPtjXaO
C7+EFThZAo50PWjZILtmSMOKP/m/7qa1Spabor/CFVfZACs08gXdDCsv6Np0uhyb
/oCL0nflUkwFb1ql3SPaiAdOpyrvO3gGx3Np/+qpeQxweL+L8EOZZkhX+RnkxKrJ
btU9KpyS6X+47wvC13oLtIbxybGrxbWFQ1Juou19j18Z6BX6Y8yjk54OLJ7l9AKr
v/WU+pyJJupm5NCOC3RRWdui7YtCK87BCAwAebYBuK5q7dsgYi59TPrmnCFxNH5I
9N5flDKJ6rmPIU2UoszKltIRHNzWOyy04Wbpx+55cvJPksBmVY1osznMPbtRrKhl
tjAZRu+rRVXoBmCzCiTO6uuCE6jYIcnvPvrQOmihW3zZ0fLS2fYGyNrHM2kvKVNx
Yw1nGd1nFKRzdzeBk6CpZ8FrdUvTV0ulyV0+wL1aqURLXf2eu/JcLLjktvlEZdB8
NE+Yz03B9y3jRlXupbTTc3s94zuTd5QXoHoLjJEKDqvHM+mmXFrLi6zGYaElQeur
aGsOCHpVJch3kPWobUzOHP1TuxworDXl8L8GN4mhrJjXmrOeuly+YkfFrsYPM+eV
AlbFxhXdAJkjGjs12qLnCHnSRoXZCwLlRdQQXFU2y3WbEvGVXTiu8MvodGs2ELin
QIcLLETLAIFJ0FMYFAP/dyRVhsqQIDP7afogdZm2in88qmTxbBsGwNxW+mUHLL3U
NdP/1kSEUMKDcCxbuZExoZqX3kfc88RLYfSG9qzg7fGmsxV9ZfY0jqiPdsYd+Ow9
491Hg2O3uN8n05sGRXSuA/7M1He2GConjWyU5+HOfdAp4Q0dDEwAuRV6OoNcLEQ+
JkzvqNJAQL18UQJP9W3KvACvpyyTnr3m40sDtgBhK/J1pmQSICGgjDbm/MPujt11
iOM1HTJce09ehVamVrhGWFWJFpvvkcY7Z7NsmUS98j+NuBX9XqiXrlZUenqh2kPH
pzokOe9yL57DmWHZ4uI2YHPy+UpORQuVYkPQrTQNBT5H7yK6ICVSoUVZ78zAS398
/UvJD1vFrbhjrzI6RXw4m6OLd84S4Vx7kTK9phvPCMEpadZ4um5Kt4hehmNk4ncf
yh1vG0j6a/EPeHT0XSDFzyDoDJ7f2E25IQRZWeWwoXYd8NVU3UiR4qCj89ScX3+C
4k8AyaQ1tW7NYQPcRjsPsNpQQgw7vFYCuXR5Gl6XqsQXtV49wUsLWF5WZVRo8BxJ
uV3u6QiwEKTjaUyvaZh1qsl5CiBRLlpACQKkcCYryln2XnEvUgMtKH9ysvOSBjJI
IAt0Mn6za0M17HV0T8xEP7jKjhz70TRKNbC+y6rICyzDPu6QMVLekRUOHx1CVG1I
Wv9NTfInUgJ11E0NUf/ZarbtRldQWYmsTa9knDXSTgVYiHyl8U74Np5k/o5Jiq5w
E7lfoImpVAkpbt8GcMiWJnLqtL1w/ta41hCYWhsLYCt6d7l10zFEIVi6grI9Pzyz
TfNELbxDzX/fGOqFJ29y/aBznwRaJiu7GQ1Hdd/3RspusotWef28qDUeqI2dRlwV
5tD9ZWfAlK0W0rcu4Cd9idKPrh6FrMfjvzhBZswwANr4KK+4VOITItTJwNzMTRHw
IphhpediSHXPMV1SKrB1Qp35cgYYJGqs9PmzMR4JhNSitJ3T8VrWXqhSL5TBy8fs
zyJZJcEfihotPbOgFDYc8BU02AoMjiiE4BOgZddPrGyjJ8sAHalWMScEG+4dH9kE
w6vENLo0X/ShA9Bb6Rxpqs2Zl7AOgguS0Pu1nz6THb93sScEtIqu69O85fK2feIT
rM0wnL5ctaWlaQgFtrFVDT1SGOjEjD/Nrn/rChFvjUJrPLE0IMLhwTsKi4O8bJoo
65HD4ZxFsjisPBg5fRr8akHFBJyKHrwwAcetRz2UeIPHl5Xi3vXlDdbwxrEs1NM/
0lt91fXggC5m6lZP8KwwCCUDq1+8C6PkyH5W8bF4jheou4S4+RxCEXEio+OUIzq8
uRTGYTDnTl7eCAVK0XcRN4aFqXnCwoYSwlXpcNoKkp+7uOiC0C5CKW2a9kSNVJb9
Oqj/Po22UPyUa1GRtnqWcRUm2ESXo2SPWRBD87BjRi+7Sswb9lXD41q79O5BNZSW
Uz00hfKFhpAgRZKTZEw98tZCxLwJaCv+S71kMXYn2m0tDqs6GwSt2eXCy03DtC75
qwY2YOcJ3bnccfAVjnBB0w5kCZ9M7ieXFuKhq5IMR/jV0IWYtmcWQ1hlayvP5PXi
icKfgruhBwcgCfkxeYJVCvMOMUUwAfnkqzl+pSuXUHBvMSviZHlp/GAs3wlQfCff
bWTK0ozjr38M7lXUBFhH0nxBAsgA6PwBeaafLcaPgzasu2kKx7D+GoWRwKB4lL2r
NedEdgu4ODRuU9LAO0lPmNQpJfacjZT2gdPIVKUb3yBAM7RYAqMD38QluHXA15uq
xBMm5wZ6ZMJSCxc2XpNomukjR8jsAFoW0Yn7f2ea1XILZSzEzMRy02isihD8A21C
nGtFQPUdSexEEQ4vmEIjZS8NpqVZhnbko9OrIRZcHvm0ug8oBRKH6Zllvi3lBXKo
F42NyO0av2wIbGjYFGo7dJpaoh3anc5jc6g2a9J7zfriwUjHEjxdBK9pMAgWb7Ti
sKMCmFyiZuFc1SeHrQkkgU/OHP4DRjtqYsBv9B9deMpcYxqIeC7BjDO6bTRGlaXx
DjTzlT55TgWGV8wrPzYL786wEfBLHE3dAopV2YTqbuSlMOb0s9GsgfNRfaSqoZts
6hM4+Gz04ZNHyo21zSWZ9VblLnC/dnjmiVMjDsSwkwgY3ZC8OzCAtfr/M7tCyK4t
iYSA5pfptqbf9LvZdp2ZfAWYYPCgibcNMzEPjy5tHJIMwyhWOo/2r3+YpN6dfudz
wNtwvIwVYbTRP7R8OzcKKiWg3pNNADRqX1CF2W98uThkZ+GcQ9vDl70KuFKm4go9
nq+D0fe/GVSqgTo/lwwaZEoSGp1SKIm1BZ6p8nhwKCnsgNQegTjghiP/C5YPbggk
etej8x5ryLOUUCosigELn0tbzVfwrVrLPQVzjW9x85MmMxkRZ3D9mSUCc/pVHOH/
ju1KwPsCr9oFkd2tAkwMHsXNEJRS/43VwENQq2TfDXswaSRWcTZWl4B0t/iSpozk
b0FCFCQwZ0elZteQhJsvs++/5WWTMGb3qv2jCy2w2/C2bspJMkH9chcUpo61eOA1
5gWM6juF/VmFD1GJ350oblSo5DubTo8CMIulZ0KIIGF/UM6QhEBIyRd6lbOeD4Sm
tL5pA8UUirePqzPbDvWegLSLQ7nG9yeE9J338g06ZDIZAircgM/bpXwCnHwQBf00
a37Fr2yPAiN+0XcqK9Pz7GeDSVElkldFuTW2NJfcGFo0M9G/jaMyuwG5rlLmRfyz
MTl1773lbKMDDn2aKZH6cfZ17S1xu6qhY1joR7bHXBSquKrASEgHzbEE4YefbKGX
zHsfLpWCxxeuM3O7BgZlvkMXW9Cu8zH7nwZYmaNFZDoTtndvIymHiUnkKfGyFOd3
VHtHABv2uALWsZpVVYs0NrVrbohERoWsNDtDvzZfzlfUrajCSUTFpWRwMf5QPdtl
cw6fk0L1jg+PGx6vAEc+CL6UC32KgruEN0UdZB/IiPJf707wzn688DCeRkNU9TXx
hw+8PeLHNae7NfK5BgZ8NZ0cXckARFYL6fdTCXCemqstO5QHfvQ+7AUHEGgvOvUz
wLscRh5ZYaZZnRkBuhcstS5Uxrs9BxY6A99GHWMYk2tOEWbvhdJOV+i13ilN/Vb5
yEALn+Y4SMV6pzycec5K3qxPbtV4WwGovCBnMeUDysNGd8mZTpQxJscFtRl4trxY
BQcy2gosndLcwL8cXl/+eJNxNgjuafkles+uf1/6yfHXzRbjrTk8jOqLqsEfH9Xb
n8qjT9XyxQ+beSMVWozRXD9bU0otX7zZ+5Uu+lpOZC/SoDXfrhi2dRlZTBSwdzOx
K8NTFgalMd/P4GqM5T2StnI2G7lgZqbY/AjMY2t7vYWdcijGq+/2XU2T3r416l8d
A/sbq6zr+PebwoW29zSfygUuu8BUEca/Uy0Tt50Vh409dRDY3Lk89IYk8cSa1ha6
+41obVqW7wGnNQ7gZo7rkVcxB7EuJUzLPkgjwXLzs7BSfLLQDc0oZ/7mR83jgsgG
jY/Pb2p1gY4D+xf0LJu+bBfmOCYDaazVWeNb7eHVgpku1QOvmoECPRQaducCt38P
zg3KBx5AMs91sWYmNW+aNV5M4FVm0Db3XvYqCIPzGuC8qCBYG/hKzETmnQq1NppP
M6YrNdnViCfP9HIcJgu7e6mTUnQyiTbzQEsWqrjJr7ebC5dlkgx2mKsA2kgHrLYn
wkR08KeI/gRKbnxt3v52Oi6kJCZcPUUqgb8aFFpsReUS8kFBvzO3gdF/p1fKB4md
A1jfrVozQxNTRHddcxT6ImbsvjOQoUzRW6gaNhFDhlJH4yDLP/fpGRF2Rv4x0BHf
W1ZgIplAEIAKi1jm63rmIwjWF1U1MeNFjcofkvePGjMtqh7SSjHeIPbvYFgf7AsE
zypOR5XGenAWIpyPSXuWtXsMepcypF/nHGim9iHfw4Sd4P+VlO+5hIQM6UvAvl4q
YFiET45qyfGdby21k1CII6BkyokuzUmV8zvtgxwGB0IlMwY3ET1p6zHgvMVMe6sl
ChpJfftz9d5ZdHGOjvlS+RdlTuMF6ralBhzPHAJn+vNzyZ2CpmIF5aGv/7JgOh1Y
59PuEIgAM3ynCytJQCD++O4eObHLl2M85kTWFR4pJ/pRgobDAa+jDTEsa+jq4M85
zHVcipeTjiIO1KxeBYSa0X9EOR+TVIN7izxfDyWNHsJ6A32W8BVVuPgtYQvDKqZk
DrhDmmGzFQMiXrm6m7ifZ6bnNZP2EL8NXw/FzHMMhcnZ3mFBtAqBLJo4mMOVgqKY
YONdLRFb0Zu+++AEbswh9OZVzBMTE7R8Xe+YGFWhJszdxaNagM57lqgjq6KljhnZ
tLcfwX8iWOPac9fc7PqDJJbKTKOAugwaUUXJ2Tk3lrb4uSKYwQzrBcVvLtnePcqg
b+SrHyM+g8MvMPny/MmjSPLuEPQoUSrpocf03EgsrbrT4vAqIKVorhAMEw1hYyFK
4urXonFuKfEh31aEX49zmAJ8ra8+UCZDQtzxHuNUSE+atOsYIZtXdQUt5hacwlmN
ZNzV13PCpTgTTZP1d+AcCNOGzscJ9XXjaVAWNOpAmTRn65P3arjU3wmsmtQWoJJa
DbDU2DFif7jrd/DFrPlCnE9gNzJ/LczrNdIS+rUvByxKhdfuou/IbW8UM8qYWIb7
ouIVtjqehSx1XM9q3Lp5id0WO08l1frbGTL+CSK8Zr3U7GhZ2oL9n9J8BNlNOEKA
yiq5adNKy13r+Iq/Kbw+Ei3CGZxS3BFdUAoA2742RfZWW+seBLDjLFungnLFNVzm
wQeTGfg6su0Kh8li/0jmVV6UNrXqFGQUwxoydr8E3z4JkpWmmcntHCYez80lS6hP
eVGY3YMFBRG4SMQ6E8xMFiYjJrDMtsNiF56UoAtO1H2iqhNLSZBm80+GvlLEXIPi
bZRoUjwyICD39xCjtE9FX0+Kv0+Dv55zFGoM7Dyd8I4y6w0Bdq5YFQFvaNNHoqs6
Pkqaz3klHpq8PaAUHsPtQBpmXcGSJdM1DCu57ROl9FAyB2Vj0DJsK6xDstFYdoFp
yd9cfUSkaf413eVT3nzgprOSWpSPP6r2I4DHpA2vIldfG8hobIbSXzMD/dLUube6
ZxYlqHHIGTIa4eVxZw2gMwinzSCwagsyWez8QAMvzF8yjChkzfKfP5ZDPSKCEuXB
hl0C/n8/501mMFPqRzLMTYd8TMvDkeI+uitYTERrthhSkEd5ED43o3TWXAwtq4Jh
h1pWecIFAeXIChUox+QZlFvW4JyY1wvVPaU6vz3EZskONptYRjENhqXUjtEa8/fn
yN+4pVdE+3v2pIsX2qEQqMf7meeVdmb4y0qyyBH63tVWRP2VIgsV7DijxL40F5eq
1UBznMhsbjkvFAVPUXCa/vV1ONETVsAESRrMnvZhm6n3Me7jHZi2aTuNJKGPc3ld
9Dh/mI2SzLRUw77MLrCI93XYpF1Lsdqbe+OfoWisCfkfNj3hoIdiQbPYB0INzx+8
xvpWqN2Di0DsE72ZiZEtLBXUpD7AhoajWUOQuKAXsul0mdlTbpQuzkgQsS/y+Cqx
Xwc8cOtr2v2o5C/QWqlDlvdLY0AfRTqaGMWshMk1+iFxNgxMe0npoElgxzZVJY7P
ND1uzs0nAtFVUchJjl2zjcZ79GH9Q2dEBXJjx6rmjlnKTXnzMuMWmuEI+pvWJTmA
AzT5SPlYvcL8tlqisOVHdyy9Py7nJXxE6i0JkoPUWG4QW0BJtqRjmuRfR1AU4Nbr
8k7W6Cg2ApiwnxIvMcmvGViMe2pjvc7figFpY1LC0BwE6i646xUzFK248GXh9Vig
RqpG2hOXYBAMwzPARsVf0Agq612NNQSJHsNH1JwBaFYaSvgqtd/e6U0R3KqjnG8r
z2VGZLkG5X1yOp9ysLSGyRkg4N84apb0WZEAeJCKurJqdE4P5katNRIQ4dM4HbJB
X3QJvHWeQ5ugKjJENiznz7a6Ulb8aeYM5iKFTM/KwwhjYQQcbspQ2D6GzdF1u/wz
YGsQ+WFrft7On+lclqKGLxS2tq/fe13n4dOwuUv/+diuQp+8Wl5j4oFqjjk+M7jB
X8Gpw/1UWPMIFvH8mYwgmP8mW5NTmOpTBspSy2nEyiXQ7DTs2CLIlGOtPcfo9Z5j
+YoXMOyfskkKrhCzig5J8mQpIUecLxrRPhfWySRyV2KoZOD2zmm5GyqNAv0WERBv
gYebFJH/VGb4cyt43Q+ZeIaLaRJNcTM4Ei4leJiMEktIXdew1vp0gn8SMYvPQ+CM
liS5SlglHwCPINXwDV8SEQ2dnTXr65Ny0rxruOboZtp6ZquuV5e68gb4fWtKRjYp
bGH3HIUh2BECrpHXMWZIIrU6RIsV5bOrxG7Hj0KkKjap6IzkBKTeWtqKyc2AeDrc
9kW6yedbJh71UI2yyTARLynjAG7Nz0gWaf248a2L/JnCnUxF3ELcArpxbZFlv4VX
hLjWHsaHwGjnLibYGctDVnIfitoy1ZQGAy1zJTFiMZH+QM9zlKgAiMoEB8QxNTtz
hjKn0LgwV+WnwzuIIrnQ12MObnWZxOlC1zHAdfNue9jxWsxhYTpuqlsCp95CTqb1
DJN5nBsj8YE7Zn4cNo09V0Ad4Qnepw9nXdYxGodYxuTtzojoMlhm35eUjnnR2thu
t6JYqwFg1CxTO6JzOa+wGcjOpeGtzOrDdKTd4IEDdBm0AsEhKEQx049XsAnpb93/
f+caTYhXZLWpBmUGEOYkIxVHIhP84COxy3skorzMeyTz1jYuA0GsoWujw94/YN46
EFTnbCQWkpf3KDSThgY1QGHJ50ARvTxFuVsaKfBNaN32lol4Clq8amC2UjIimtbc
pPxXUsEgV70M+17Sbokw4RH8J+RCQbxrdzAv97FL73iVPsYUhd/NxrEob1zKQPbB
3aVs0lyZlR7I2zKVxNxM4LRYro90C+z0VMvsGaCfYEgPeiApcAI1QpcxwCJH+1A5
JGGQ7Fq9qcOkUqVAxcWx3X1Cr9L+eZTIS03iK+SuIs+IRic3piRayXUPAQMM/Cbh
W2MPC17/PiYJimt11eGoreyguvrmEcNxp0Juo7P9a9yibT1+fJU4muq0WkJjS9RS
Le+68F5m6LljYLDKlN1d/MGar7I/WCgkrL9LVKeh3Fx6VfGoNa997kO0cG8oUetg
aMrL0Ng62a2qgz3G0gKGE4ABcpT/icaSAXOoUVhju4f2BYoKDIDy8EN5PwUFXf8Z
tWp9vNzCO0pPQc20rp/XrAAcW1bOTAsrHLEDr96qIJuxE1yzpB/kQRAN7Q0cQJ2Y
UHpLgBhMWArqAuiIBefzayniTFgElIP2ZA1NlmztR2u4Ya05UXxCwd47Gl4KrShz
7qc2lQA0fEuXaoRYXdpkO3AqVRPdcLXpR1NgGNWsYElkOp7m/Dh0RKCdA6Uox6Bp
GEK1Mlu6n9YCDRDFpWsOHfsV//RqHErgb/88DCaL9bAuJlTDSndHZfEeZxzSzIXC
4qnWw6w4/4s+eU4qzO/YfbtHpYZDC2w0nw6aEw5/V0SpOsixcjmy2AWIsGcxplWl
L5B9xDTQ8KstD30h6/yjdtbhStkeiEnlHA6uaq4GIywOsiYI/7xru9c7dgV9G5k0
EcSrDaGZvx4OdTgPw6n1pWjNWAJLYWfMxfe2ADkkWQwl8wdKXLWJSya9cWzXu6rP
7ppmeMQGyijjoEyUbpkryHVRuY84Pubkiz5BWA9t6R8/1SMvGNEWE1bB7rr0nqb7
mkGL2/DV/qGR0kx6ad67cYsEPvulXv/PnigC6ZBvqM6zjIHpV0ipDNo4I9UJYJSE
ZwtnV74v+331M4dR+5/1RI/m5S0sC6sakOVOjZSfCh8yUcz00ptqZcyZk9LWKrns
U1EhWcjoUGAF0movaUK+zYnmClpRnx7R1eaYuEpqA51VYqJGrOTqIA1gLA7l0IjE
LfL8rFBSMKMZeREq0TVigjsEokFiVU4SQ65Lh6qkv5gWk6y1XZIrPXSN73lleBEp
RprqxBIbZV8AoDTNlcgc3aKpsC/iFKESYaCZf3KpiLLQjZj89EVUQO/drkLJqWh/
Vb3hFjAyps6lAaHX/eTpYHO0/x9tO2YVj9Io7JmhLridVVuHKeltPQl7Oc46kcfk
2Qp3eqFolKGMWPlaLm0mAAfjsRYz+m/iL0EGa6m1SYZiJntNYOcanQTq+oEEn7jj
WdZrb361yO1YPacC+pTV4NmN4NjwEDGPkHr3MUa3ZQJCc6yAk2z1k+nPbhxvFAgv
QmGedZ7R0SWg4dSi1f6zZSZVZvP/yNW8z1rh9+H4N2RDs5VH3wZ9aOcp5EnW3nNo
Yl+nK75ur+FASu8FZc4HhzgVBmqDXch5wfkBSSuCBGSoiVgd+CfwhypGtsaB3aOx
FvA8tkoa0mejYK/Z5lJX5OSSrkVF7xQ31zXGUFj7nsFKipQbs8Br2anjW38mStYr
oiWlvZYJCfcGl2x4j3xklJHu71sApbuUlLyb/wdiPnW6j9vLXuUD/1vDYxDTYuCz
RZ3wVDW/WhANq3RJ4rqByZhBbfW15/1cjoW5siuA1RBvDO172dso4LxDeCTizexW
XctXvtThCE+RFiDf+mcsgCyDr8aOI4Lu1duPXyb385webcO6OtzQRkuv7HYQH7uv
rnReK3sb6YhD1klB/IH5Tq8mFOpCtRgYlmH8FHMNMdkMWM4c+UMW5+mp6mva570O
WB5Kki2P9nQ9t+r7X91dw+xSCPesNq8hizl4stVP10Da+D3pzAwFYaEE5A9h5BKU
5589nVtBHKTTYjFZswHa6NGYfko1M/ed6npcq5IS9A/fueHXn55IGPReYnMq7PC2
0HLE/GnKcvQKE4+eQnDszTdqF0HohRcLvWoEnwGVDwsOW4ITfHo0ql3PLPhE19HG
XuLK4+E9S6iBSLYrvpcruHoeDkmiuRrJovpXc5BmbD7F0NTszPmknagBZ3g1BtuZ
BtjsytWYXUwUhc5kuA9sBHMdZ7jB2Tp5Vc+liqvbUOeLmeKXxnEFcXUShE/Ivy8B
72+Kvx7yoTEjCBFMx5TM7dqbx+kCOOepKJr3/tSVwJc1oQfmmZ0OoiCLpzVNWBql
t0PEqdlq5r83pbp5cKRq6LWfmlNpwz87cRNIRA4krFd+1gY7ov7KBy1GrEZ/cwNQ
TWJwoPN2hXkqqZsMKqlmVxHnGv+Gjg0Mo3TshEZcNEheaoFFvNBvI1pn4ld1bNty
FhOgAUYHp2KH1MR22lMmdxW8uFiqsoedRVb3SB9qSv2tDHHeWon9J1dTy8oJbqfm
5SVc1jQgphsCM9Mck9q6uYah0Y9GjDw1PoBpRvccfeBAm9M58E+ZQn03vjC0E2iZ
kSwcriUPNxjkogXLlVw5hTVkfuWw6XTMU0mrFErIKlUp82guxqODcihw/z5I7yTl
g01LUVsa9NNpZpiXJLqCD/tz5PARtddNksKfcG0hWOqw82kKOkgr9Nd0nlnEw52K
zqbVKB5oGNahe0CIixEfWTk0+ndsZvI1aDLDYmiIy+OlY4U/46QKaz1QViZDhvbf
fa+j8p8/9awlZn92MbGJ0qCdo4rI36PFNPIjVz1Zr8qlwTYJqQdhIs9ZGTA0NBzP
TH0xTlZ6JurlnwRxtA4qPgJIcpp59lrFoOgVVmm20363BQKu12MDHCqds7OnZ4Di
WOma+zluQkjsskdXh1WHgHeSM67v5LwmZObjM7e8yZk3sqZnJledmEc5TWeoAAiW
V1pEDg0XV41dxxG46tXZrZ+YLt8dPA53DFmus8mfzKrHPwW0w0X3qOmiKnQfFBkm
xVHcUrIyjoKA09Eb+MzO3qtCpLGwYnDRZpJRqcPcSOzAwavq0jS75EJrp1IpVnoF
A/IuJwWVavlwbXXhKXm0E06rGxrAsMfb/N2tj0QZVnYwDk43e9J6ijFIwwuq1Qdb
h76bQ2badih355EJTGvdgHIdyzAWF0mmxnLephBLQFZlZMl2MtC6+pW47ebR7A7c
ZX7aHNoKEbVvy296IvtiokVA6289Q0K4607mSckozOSb8XVkPj3/q9gFpP+Nx2IK
oGZF96MKmH+cLc9gHblQU5O7iSHpsm4zk2ijTH5jaywPnbvs9+FqIjcgJ9Dgd/iL
8qLqLAJVEBmDR66ws/CtcnMCmPU7uWtFJfF020tFZdcQFdDb/5br0ja/CM45Q8ir
TGurRqoSLttwjd7/ifZo2pBt8IM+I91FqVLDVxRW3tqPX0t/szMYfZDMQ5wyq/JY
fkIvy1V9WPXXVmSWT0M30eorbWZSORU/g7v86oIEWWwv4XCq6l0bT1EvJT/8VaJL
Mu8W/DOvMjRrQO048R9BL+ImK/69QKiaVs2/rvhNmLrEsyirZVh05CJ0gJPh34vz
JN/zYScTBYDM9V1yMexhTLzeanpBEvaBaF1j9P8gSj9IblwP6VL6c6PKWyxdo0P+
ow0T2Kc90Z4fg3aKriPhmkdNWcXcByO5JdZicEPIEBI8bduEhqcO4jZRRkOk1v1S
OQGufXzsrOU7qtI5V8+k60wsie8u9SCoMpetyOh7ePDK2ikDQsI3nKoBYe6NL05f
sRzY+vHHg3PlHmX7T9t94X0kMBE7WPz9wIHKCU4b5WLnNTXlc3FGsq2d1iTutMEQ
BEFDJbmRQo2Ea973Lkj/9yQm0vV7PnLMusH2qEPfdwdrEPTGYZ9eJuKp7ljTiRqt
ttrp8iQNM3dNC5kXezaxe3m69ZhINO5CkpSXsSkQrb4zOAwp72SNuuZo0YtaC7Vd
APwFSuvH9JQRHtnjTrek8Smma0s5lv/OPCMd4s0T8DxsZqEVy7djPYkceDNfFuYA
Y/ysXr0zGu5LKJq0FqklKf6k437uJQ36zbouMdQUsFrdRDY0JBI+jacEm6dHesIv
SL1AXo3Yr0x7YA6I9ruHdslCWeITHwdf/6QC1Cs1Hx0oNyJBGB1XtkWLqEt1oUFP
0zDYhgFABi+uwQ2jQnLNnlgfCFwAGytZ/ulHA3dXm7N++ICSUzpek17RpQmM53O+
s3Sw5GeL+6VSok4OPp4Ve7wuU0ANSQXtXfuttTRNn5tOCWjePxwxVR4vD8nVwBe1
FwRdZCULk7k4iEhSS5t1R5PdEIbtOoTPxlNf9OSnay4WFK8RhTG18rd8ut3i41gy
+kAjGlYuh88nxut6zs1vohU2yvrrZwGvV3cz3OASUWbitZx0XIK6pasDQsk6H1DZ
2wuABYa7y8F2xKXtyJBRlIjP4tt9nNI743wwfZK8Lobose+ndIdCTGLdCNoJKkJd
vfD2EQXOf7VzVIWmafVeP9h3uo1xmQ0yoZSBMEBqCREGeBj/wf13fiwdpAh6/6l+
5lWP1FAd16ukl4pq7I5aqzmJmSlmmrtg4EW65nrXssKLHt0iKRtlkD+G5Vjlvg2f
jZteMMYNgAKyVV51l1zpJFF/a65oG9EBYswvs0qJ9Qvl+PW8+gaw7Ucm2pF5DCVZ
b88wnVkFdCHTNGrSYr8TGbqU6ehrNFxnoGa7YRW1YbAJAsCY1fomBL0l7daaRcYb
Xvbjk/TgWTjZoAjxKAqLv836cAHDYmGcc1srVWt6DmfO4suaGZCoH9N8412DlyjE
h59MSrtIQ+xXRRH81WKJFMC2olkVmMqum9Hdr7zQMsGsXsiLnu13CMcUCvm49Kb1
UX8VNDy9cUmBdOH2gU9jBuAJYNkkrd4jmZmJyDjtFyoj6PLuSI9kEUA1P5x7Quql
kf62+zdz0brBgmwxYuWJVBpSV/iue9mxTMluLP8KAZ0VTTMdBqAkO8O/tN7CKIg1
mrj0UWGN86nazOTHJptqGAkIPdb14ZPZXH/fahbOEw3pu78KwpSmZ8WHXENsch3C
7BSLnALdqXRYHfc3058KqnbolGSTr/MRBGGj43OHxBWcM0Zw8uU7xkgLIouDwHMK
1F4hqnMkaR4NJC26DfhZUj/A0FZj5HPQObSGJFQjzE6PFeP4T5dazBt3RjuD/A4D
DUfRnHJjvpVtpg+oFwr2JMwf7kxpx1+v5GAPpwMkc0CXq3/pN0Jsr3gtAvBu9303
dmbRwSPvRncQRgDRA/z15GVTKbgKM+kdLkg1qYNkBctWOo7UnjlvPDKX7JWv6uw4
3oaXmVm0FvD33nOodozXBJgmpiGYiRZWDMnL7KV7ByudTmgQKwuIrjIP9N+olXrt
oRutXBfI37C8W5rMC00VmjVSfNUYsht6qHvLe+8ThldJRvIRITh4XxoJe0e8XRFs
xxbNttaEbnxREGiANv7k4GKxkkM6oGqqTPaERQlluBiNBUGbDm1wIwYNXyRcHqql
fcIi3vVpICQOoJWggEIJvWGAmgWLg2HAyP3hggM/C9t/RhQbjPoxukNYO+fns9iw
RBm4VR/AZi30OtvLOL6n9OzKZrpkznCmJd4289cRqsxG6pl778NdB6OSRt8LLW7u
uylYv/hHgL6b8MzchRKF5XRWasnWgekfWO3ivKsAUR3CGCjBc6a+saU/UgrnUmGd
3QzltMK1MrxYzTUcZUymC/EfCk7+RAmgxRgPzB7DYVTBT05toQ3K23WySVugt+xS
CRPNB/ThGKN1WFonRjtYzV8UEiV+hEhmh1q1MVYh5Czx48EM6+CbuTHl3aqlm1HD
JMpvb5QOhw63+kqTKXNlcm0e0YTgKSbyWpWBw8Km3wIod1TJPDZNgYeDM25ng+NT
5MrMlwlqGhVoZQaQE4+rB0xStZzjaMGINPPhu0HrwL8KU+Y2OrHz1vdHFNHpcXKu
MKN8IJY+ZLjUih5MoYbcu9VAOMU2lbKs12bZsskU/CyMmCJShNRFvUa8gtD9354u
Lfz2sksfhwaiKn/7FEUoXfIWJARY9YJGhCHa91/Aa4JQPvNKHUWHWup31UEoHs4j
dRAzxuyzHCyQ5eAQ0+A9EaE9JLCWn0oupwzy1r8bcyjSwFQFKPMC59fmA5ReFMjr
ScdtgxJoG4Bd2mvnMcwibJGmGc0HBWvMQLWjw3LpqhcF2YJZV46yaCJ2Ki9zdUhM
JNJVDkbEcRbFQgJYAJnnYICkMhdsF2pec2LDpisTvCKAr5pYM1muocDlu+sPgpAE
AzZVBR8qkj4I3WB3BWiqaxchcOs0dVtRl5WUDgXkxu2vlT9a01WhY2MfY5s3Vlgq
4uw/d02VD6sc4y3u1dHO7PvBimKhKqay/m3aPAGyoGcA7d0Bgywh543h16DsrTlJ
qWKLgdVaprbHGDp6ftPpYBeZtYUkTcs/mnW83ok8KtsPwRCfKNmWaNnIArFFjmuO
KXz9hODcnoGUEgDCM/h1riVpKp3cvp9VhQ9Stpxv30/t0pcQwPl3nppynY6M7uS7
2cBrEknrJr6YzSua5qTwZ9krgDsLjf1VTPtoFsMlDDmjb10tzERU2l98QJ01vvHK
xrqBVBnMxkAmvR+WgCWnK6hGyWIlL4h2DODXUGP6hPH5bucSvtMrukb6tecnHi0t
flxLG0dYI/fqf55ngHPyKZ88r6apMyWf69G2+gknNw2nyTyKL0JqhtC89zbqsD8P
Q3KIdQ0wpFe3XM8kPlu3h8NBVM/hDCbRN5SaYfpiKXMdFw83InTLoGckhNOXyXnT
fsPXsEVaA/t1z1f/woTLaywNRXGlURL6ZMfAH8IRkEkgxt4tauATrSr2Du8pQCuN
U99g1jax3gsT30WXP/bP9/2nDN57XkfhnNEbrPRSncdpnEwoinZ4F4YSPRE6lnJf
Tyvhe/8GANcS5IrRIhPXv2JzbBc6LxpJFmc6VdW05gtbyvRCZ2kgUx/jn1SrQKTD
i3G8yHE6BTlHblHbFOWWMNSWegyqFRsesebm6d7l3DEQf7rGFZwdUYqrEIbLTfjz
HLXGe7FBY7MCm+il+PR07V8N0qlsfP1BpNrCdnqd8Lgfp4OOi8ukIagyS+hC1e5E
XRk0AewjHTUDMDtostR8dEVThIj4NtyQH3RlLqTjcqjiM+jYFBHorzq4wwCYCZsR
z9rmI9V2X6CrCoac1z7lLsS4Xry9RViFa5RGqgQY6vbncGX0lX0wCA20q13dvnOf
mbvnrePqTpNXiQobN8hZkYjLqgcIu54ltEKSvyRhnF4MWx0U1aisiBlViCY6Us30
GmEwcvBBDbFSAHMj0eeKNFnvTg6CxOxk4auMFRRZ+ak36sN32MCtd8F96RbOoN9Z
FysJWCuiaJ8R6Ff1Pg31K4UdMc3cCDpzHWQt7/88omiN6aqrEf+Qm8IM24vfOQAz
uJCMgs66U5PaCv088mCU+RleuMOS/Bcy3YA3jp3LcLQn3TbdR/YDupH9PZJQtssO
gYg5Zu/4gmADitVHmY5s7lf1vy0UL5QnjW4EsJURNYdQo07Z1KB9SyJhCBoeV4W6
z72MRRDAL7JRr44M+xhKDVFmeZZglmAzi/urhyKdjPARV6pLqcwW9Obc9kir6a1m
Qe56wvOSQnfnT3rbVoYI7Gm1bKMk6NKWqX8H3YkTr1nSyguS7gMf6K7kfytt10c3
8YYT1txfL7Mjmsj1qEQV6HEClA6nFETxgI2poWWa8dtvOCiCq2dm0JNYcAWbAAOt
uVh97piLu2dxZJkf5DeyIdeF8yq8H9cEYwYXHtxhHeHtXLvxCwlgj4n2DvuG+wQd
THCAsPSXPZsW5f4vs4fjko5Xbp65v9EpBpIPD2sKICvHqVEkTjbDSAcfWxXzMwI1
+A9sigICkLB0+eptsYcGh6WZFI7+KYG44vapdmsBtjVP3W1gLfuiAjb7WaQnZF95
Nxibj31PPZZxDmgG95Pb9uOf1BHcBfAgF7jgjqgJwv5bVPYm6guPxLQZ1r/fxfpp
Un0J9+A2v5vTW/hz4kSDOLFp1zP6+8no5PFbK1CmAjyRDlDFHcvJKsaLB+F91SIU
EKLx47qF6dVCEHZjsyaAfiLtQdS+dAqlKWx7wF5Di2psDgcZcPIEngkGuFjPrzAp
ehgBn/OMBMARM+2M0bm8hkWjVwPz8EYGTRv4187lVxLboZ5qbffz3NLwsJtRBbhG
x7GEVsvms5S8pHloXV3Qt+Ur1eX0rM9GxhOacRtXbagvLvhsr/qWYVZfzSkSZJIO
FvW3uc5c6zk3TiJlsZlFmqXDrrsAYS7kcvFvTQAr9uiz3Y0B1IZOnbvfwRmXtnIZ
d8x5Yfre9d7tlH0N8reld3BV/aCNTXajCBIqtu/uxMSl5lmx1lHZpISNfV/Qw9Xg
UGMj3Le+dyFPXLHSj51huA+omKpZIikx0M4NgCaNtKIwIJFIcoZ5jwphtof2opa9
1VWuD2yB4WAo2gy4o4nTGG+WgZyJD6bPWfjD6ei2DC4D1iio0GBTcdKy4lbiEgZ6
VemBlncD5KXgUJ0+ZDTkCgtXWZI8cS2h/xzUjp9OacI877zqiqpI54dk4ZvIaISt
lhGHkOUiFHWOJgn/PxhWuMTvQwIiNksR460L72j/1saBnvI1cHoEznZ0RzPLpKRu
cr5p/se1+p1yroeOyhxZOPjMCm6G1WZm4ir6xpU5ylzNGf0aJhdgbiZ+5B99CTZB
NPIa96UZzShVq7Wu0LfzfvXofyCZFRsGSBSt504QlhVJNZ5jqC96HlflP7VvXwc3
QBMHVDo9S2s95UAFteXybD353hz3ay31J0jWN6NR+V7Dl5I24kugjNJtwbhG/mOW
bIqv1H/27wf2OVo+FsG02lXO26Plxw1SMJ+oJi2E+5I8Cje8vJNMb8U0tDAwNcBA
W7ciDOj4PihfPRJX8Sl7CSIiOZq9sjaiwldPcKCKHChUfJd23PxzjMPn6nkr/6lX
gxJs7SAyR6lFBKumzKKGSSUs3f8MppEnXDR4uUIB9lpFF9SBJZ+s/+A/ffLeQVxO
6CSMQWFIap0iAb6OaHUdPvoYqHo9MIfsKJAjohLd84L7YFtNqQAnPddrVU0Bna3+
9WPY84aMj0FMXhgM8vThf8EcO7QzeO+G7e7yBgqAI/Bh7psXOlEYGNoD8mMZA1or
UFNvreq6MK8IDdoz3x8tf6pV8zfW9/V/K4XY812JzKjlErzYXcvsw6HA0AM9mTAI
kfJg6LY9azI3ZtDRLKY1vm+252LvkjBKYM5u6WlhU6+9qB0bIUYOoL8mcAc6FmfB
3bfcUjbcXfPWW36NaRhhSp8wNZz1OjY+Uh6UdVvfmmNJ0EHdj5EjbRsfnAKGcuHR
uHuNWYWtrpLmZ5/zo4LcOTw19HEMwHYhn5eGG0y9eyk=
`protect end_protected