`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 12176 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/59UwEX+aE7FohaWu0/8IpTj7mav863zUNIsgIH2BWb
Abd9opeuBjbGF/waQMI2vMJTwD1ie1YueHc3nSNpEh4OXp8P5ybZFY89uyGz3ztU
W1EsuUnchJoQgbHZ/sLbgtGRgsrAFn+ZoIeGN1d6RAF2wAESJmYP8zw+p00RvjZ5
heIpmLmrzD5nzvK4jElYdCUVOwZta+uD/pnzZmXEnthUwtWUCgki/griyvUnPVTs
QjxjbGbIOZPBxHbXB7pcS7DYYOn8SHV+DLS63TcFfPhaK8ylGVtoGINOaJVIgGbL
ZU2uiYsknlHT8qCuMOHz01omWPdxM4PqtTD6DyPgmgq/U+QwkJmy27IJyCby4YB3
Oh7+/ah1zzvbCZDgnlzrNMYBt/lygGBXRFoRiiNVHSRzre1u9DqYFisj28osmUal
Cj6LF7qD7hKSrAgTgrpjp4sX5T6UK9CElJdwU5iIt5tBTMaZjgyvvA1mu/ylI7Ev
XFtXRiJjnkU1GSP0tX0naDTQNpA/yJYbnySK4lvyBQodhwoJmAJhme4IWAZVRtwJ
REyGJiRahoLk3wJloU59YOQIwZg8VdFPmQfC+SvF8XdQ/gmjX+1OdC6TsPYefhBf
qLYo26RotfWv6pQI87/h7lE23SdXZoidu7Mxwvym6mC3DublxzgiDfG3kLhtGwF7
k6N6go0L7zn8LSrgGANVDKIwEonGe8EKA8NyP5PFG8F7dfcBreVkYzcVyvjwnHEz
Klvu1ohdq/frCzFs/rbA/qOTJHV3E0A74+06dowualgC1sxN6BbOUB6rG5L4OLsl
ri85Kt6zAlozANuqyiMVOQj1hfbAOO3JMbSzhGjHWhozqP8fVmzYQY9rxyptwFmj
l3KbL4zQcOenhtL4LUBoJkSSOYnSASOJF5p2T/o6z/jt+Lb8fkP+427jH+DFYEag
J/oHSQGnKzj7Xd0/EwirfY3jrauxyLNnMZAFcJivtUI9x9ZbuKKt/kGIMk3F/YvI
9DBo3o4KKE28iB5VRd1Gq1LM4ie41U39xP6IeXEIk2NVzRu6tV+7FcZVKF989+aW
p6EurqRNsLUq1l9puZKbVgVwMrLrEPNuEsYTYATBKJPts6RxaMgaS7pfXBev5V/Z
wzmASvGpLn2T19IXciOkyR+zzR3Z8W1kmjta4glOtr3edbrHze6P6YTsJ9XXthiU
PVUKCf1/0I4fFlvSJ6bg8ABwNzKo40+ualtCHmTEtMEtnBwta838vcj6lQYeAKep
XE2yODfmqeEME4u1/LEoB6+thoPbU15qmkj7Lnvu+2G25gmuytb0UXLUUfFf+zmd
0ZUbFZln+9L1tylkdGKHN7NQOtlj+S5m1gWq9yUnY+yFWZZETN0kA6f/ebUaW16O
krZVDlqFGNKpOYIO5T2v5fxuNWEOA1Xac29lvezcyQcYK7RTIUnd3mD7KFknMxnk
IjgKeBdyKKysuvT7puEmLbXAWB9z1IA8ORKjm6Rvr5eilIRXXQvpVvmRu0s6R3hI
lzfQ17FB8NXSNdcGFbDS5mTIj4IoxGCjesINh6GLsfUkrYwseUAr/8EuynPWhlzk
+NR9uE/eSdisD0w7LfDwwOzPF4s4H5CGvMhXVFVlJuNQEUuzpLtkYkzfEuz3gPwM
ruapFc/pCrLksUS0Gpp8HM6eBr2wJca7DfGDXxJN5Ow6pgCKJ+uvyu7UbbyCwc5F
3C1CQ5x5ysOTAQFeNdZCCct8tlTS9XzW1ZL7acohJIjRooLhWd9RkUqldYKyAo6G
WbK5DZ4wp5dxBqqVe25uXv/Pcz+dQ5QIhyrWQxyY5Qb76PwTgdF7HAI19FesdIdt
2C4OCzFAaFj8ET66h2Ezv/4BGepZG95copPZJLJn0VPeI1iYHRonDBpwEzvyEPlX
5zy/Fktm0Ib7exhQN1itsIML4Ot4JPNjN9Jlqlsacg3pybxvJCxvm2K8HxcdUCb5
zB1wwWcJjlr3fsypxnD6B939VgVfSVx4kYcMLGG+YY/cwlEpbd/VGW5U1W3mykqu
9HPJ06rO4LokKozM7fK7Y/b3qoLxpPzQcZFgSYVoqq3tnzCJUsXtwyUqQ4ox/S97
WrGHAW2pgx/GKvReqaW4KgT5q6Rq63Ptjc0rHOw3GRu1YwJQgH1+A1XWIZw7UQqG
nfD7KucBSqv0beZGkQOerpDFuP3ayW6FuXzRaWF6uC0oxEiu2M2HYhRCj6dJpzmP
/oERdN24+fFKRQ9lTCP8MP26EkDOC9cM8AcXfEmi2ziPQFx644jo4DKI5rd9c26b
aL3/27Bxq7WjGiOxDcYEcBCQuXLzTY+9pmVpo4d6QwhmTlMfBI6vbmQnjZwDrxC3
Qwxek7WMCNsgqG17pjjugD7I986msKd/C7xuUc/NsUHvjEYzySmu80lJBGWMJxzT
+qyjiLeCdF5QVnpR6YolDpzLonhhNvrMyS2b02fXT3ZUpfwMEmDWx76maV9Pkt9h
ndL5jFi1vRUq0fgW9Qz3R3/cTYq1Tb2JVcuHmBqnNIzrAKhJEz+dMR+P43ur4cfl
H/CXB8gDpYXJisJRznA2rXI8JYOkaceMPW7gnGlqtHO/9tzJ9O+rIuJgp4yDAVkI
N9FQaFifryCwIewGcjAeFPcJn3pcfbzE7/TVof7nsCYiDvGWfjVOKgqEC/85bahx
2R4ZNSCF3sfCaSeKRwBe0gFE9fPXd9dpvpSGOaJ+TEOjSbxkH2b2SDr6oA/AlEcu
KrkMmmeB6H5wx9f1647bk6lTxgkeqoFdV+uwmZJwqYOAeX8YrrZJTXFozbn0twYf
CvcvLNb/q8c8+c5L2Wcfl+dQOuwrXj4JiFaRRssn6Zn28hWr6Zp2TnEEAz9pfcm7
itV1+pBo3Xb0rS0GxF5oEwt12fiUeNQDfWU2S3Hly+sCsyMpz+7mfXuON495dS9d
HX+3zzD7bOWCAHY9wP/LCZ093SEQaUJDYlt1cXUUWX4+CSIx6XNr390iLvz1mURx
OXvwpSDekFRde00jO5/v+OyVmkI/4ZQQS8fJJBxgQn0y4v1jCr5KphcsvbqL2wCS
/4MfCAIe7PYgmzGidp7Ar0xnT5VtsQQqy2mgdCHlnryQfZYhfGKHxBnnbAo6H9EH
MFzCAK6p6qv/xAMeZVSbXCkJOroS7xGif5gBqMC9dWru0GV6V+kPOJQg0awjU5f5
bk4tl2E9canUkJRdOW6gVmb2iCSF6va2LeQ8I6alSYze7ZfbEdR2QawRulQd6Vn0
gSB18g7Q2NtHH7o0LYPKjFwCXVWSJ0n0Xe8jjY2nMSiWLqwl5XchlRf094NBCGgH
eQPpgyDs3E9lE0cQaX8BdjLom6/YeFe8Uz2A8/MVPCoxIRlh6Mvz8HWTo6g5CDlY
WkkKDeLlzHpQnx2K1BCxwfOgFykj/OOLC/CB5LxteAjBb2CIu2A0w0NQ/eO8V5jS
EREJo7heoYxEqXzZ+w/6N+LeacrhRgtm+jbcSojnjAAWxHIyYu77vufXGBeeX23L
IoRMOVwWrEBfGKCPYN9rqsknNFaXjzCl8nx7SFxNAzigoWs/qT54iSsMMcEHgm87
2YnJaZ4Ewv9C0sXk61rQQqpPlcDPu2JetfGYFRpNn42b2nSZOaYml7oCrWkYPDPV
vVW7lxDjw8wcE2MOCuMh4ecx1G1Hn8clI5YMHXStNOYfWe3RKeaqboz09LQJJ6CX
2QcJcZlHLZN0cVvuy9lW0cDMPVA7GJ/DdYbSrXfMkNwBmrtv0VpR7jKFTXK+VUdk
+dqUSCGfFQyq7+9yQU5qtrBoZCuahtI5fAyvYz2r4g8CQp1ioUnhlQtL02QpmTEV
DANMGKw+VR9f72BF4SfWkJ7eXpPRKNHt8N+yVVclIgPFXhq9zAegUYEnxaWwUJqx
UEPljvRNBv4AkxIWgABF3G0lP37wye704XinRC3qf++oI/4l1tZqq0XcZZ72PQw1
uDTT0KEkbijFUBJ7VZ5wDMTC2T4O0hhOvXbfxXN71eZHqfjb/2rYA2hM5Z1qA4lR
a4GVH6VIATTK44fx1iR+q/R7MbBpCo1czEAWQkR+qAJ8iX8UIaXawt7BmFanpiEu
HWTFzNzgtafWUjDih+FnaWiafODxvMY5lapDb51l3lpJGkNdJRt8xGXXHWeK6V1Q
5G+QWIP/waEYdkHdgkoQYN7SYjCgcx2kHj/FBVoru9/FmA0S3jvPrs8wGu2dXQxu
WvYrJ33K0hMeDrpo9pMMLr2baVp7hjL2TfX75At1nBIADL0nBMYCNI9E8NaFIGr2
OVlqlqC6GqY292oPMz2eksWl4vNd8Yf2qmq1TW6EJnRwnNePULFCaNFD+M05kdaw
l4JpfM2eipE77gRznvjtNub2yblsoKrT07Gk0FAoeQRk+e09BOqO1p378teuRRRq
61ixej3SV3LzunOIuUSPSqoYtztO/817Xsmg9uWH3hqamuhcOeQ3DAEg69PyhqD2
0OFYNHa7/GUW3hN3VoZH9ag5jqzldmWTb1SmOYwYffMCcubTch17/GiiIu+YITSh
vjHok6C1+0Hl421WHGvGkYZ9qnmkuU1ofDhMvHGiTjte7DBMdjNmMsYZ9jjFDM/Q
DAMGud06Ilq/KYOuKOjSMfgVGJhOUZixlCpNmUODB0SpLqAGyx/oqhdUCnGenGjj
u7huNcNulQ7MfDJOP1AguW0qLhyhKvlEWwNfNPYlYYvmkykxJyAKKD0j8uHByvCz
Fsik5VJBnCxQGSjdeGh8pd1PnSvbt4T4RKzFl9MGEUY30xE6/BoC0GrcBb+BvbkM
vlrDOFXUt1rRkCAxhAu22/hpbRVyfMM06oD5ue1ebERRZb9MrrKzUipo4xlQTaK3
KrfhiZOHLdXap522Uw3iDkMR6lvi3JCjK+B1ShlXoNju3hQW+jmv+l+7WfQbP8eq
G1ka9RO8cc5GeSbmv0v8ZNCZx4bAzzNnKgeKayT2HdCoOW4hvY6hNzFBVMtGOGPG
7cyCczNrR/8UvF8qzKf/1PYqovoeQ/6sKYfT7ScZZFtGD+XBp4TgJ/vtra3Fa+oE
0EWApNcd6hz11Rh1E75akQ2lG0cRS6eNoiDzUwQlnegjs+xGS4ucFpdmpoDygWob
k3hh4Vck8DpI8LqYNn4br/lQIGtyxdNAH7QSue032vjrAdQpybjRRWAhEjHPla5J
0HNxTbZbryzG5WPaG6Xz3hlUNNxU1DiYIypT6+QZjbUowxjQ/HVTMUlV19eXX+Xg
UBuAAq1j1429Cix0Z574uWgh7an5WGVxjAFA18rAP3F7asq4pvKm1svZT3Ij0RiC
Ry9ixsFqFhlWUGPXDCvVHChMsfTVyS2yO5OFX+JwnnQGqxBVcbkTuW5dlmpgqDem
hR2BgOGjISxJM7K/k5Rglzv7RZJXwnWSZz/AAGityY/xUKrTScnMTMkMNoT+EMq3
JIN18T/P/kAXYV+c37WIT9op8S7meErIfNIaplQFv846vNs8MxPy15C803TSlJIt
UXsOSkOlVA2CmzCcHfKJ+s2Ha8mqI+rfTw0rBJPmI76doJK/XaQy+TvLcQtyVru+
wffIriwjQL/vGPetHkN0M0iLXEpQyg308WaSJj5eB/FtDSmKQdKfkcEee93bIs6m
2UOlSjpb10m8T40btzaezttXO5w0OqGgJsUiDbLmv35T5Z0elHzTjB36Hlp1LlEG
6ByZa/3Hs/Bud+RvNispjFpl9tA8Vxa0nHUVpfaiUK5QQpaRsuGRYx5Iwwlj2NlF
P423ySDnqFQLR0dA8ec1BTk4xVUIEJdZ68uBgMEySGiCm9oZ1qAn92leP/cJUA3n
2jHOPbf4ctD1+/8vNZ8uoA+90xoxkdotKY1Or9RQB8gHyp26iNxNi/ZsEbejHg8j
hH8zGeGq3oWeW9oHQn8rJ6scWCTE9UFldDYdcET7J71U6zm47hBckjYffLQOpDsP
OWo8xayQPjNLbLQU8NjmG8w8V5SeXJ+QeoOmwrK59KMFd4/NFii61//1YbQ9dLsV
q25yA7q9u5uXMjh2drqxTDrHDJbWdQiI5PYzHLSymQl6so9b0P63yOAWe7ufy4UZ
fCbJQ9WfVpvEuSkyJm0mAdESg47YPNrYbZS5DReYyuw7tWtPj4V0jU78WTLph66g
AiEb/LQ+pKLu+EyIG/jA39KR7CY2tKACbr2tTv5HS5bBodTUA5V/4tjYl91HezRo
xaGgFpnNB+dy7GlEQjm3QbNK9l9PVZeCKoHVt5QxAUZVQldQlphiPxRJKYZwHPgK
zq0Rvj1Dn60OzsG3QTzS+HTY/Al4p/kk3k9/Jam6vREGnU0o+hts/YshTw+q+Luf
2ZZcPntiW8dGk39nb2a4+y3AaPuYmhpzfPrHoasjly+dfuhijaaX/3SpMf4K93/w
c8L84NaAMdiUx5cfpRtaFKG2jMOFlEMmWxAxGGejZkrc7kD11IkmcDGFYTvLTNtr
1Q536CbC5XMgZoHVrhCkNVOo+b/YoTkS61aaYQKpli5o8zogtpWpZXWqo+bfvgTN
HbafQCw5vxQvvy8GUEIpyNSdyojQMuEwNMer1fM1Z8rT0+3mwaYl85LpYCfLL+ci
5JaQoog9D7/Hp8upnUCRNPjBb5dRAC+y5dxUUzsUeFKCOOXBkgoxupPIfDE2WTgP
ym8iADqoH5G1vB7yAWng6DvsNP2a4HtfF6KIg/mmbylpToIqNZbwhW2cuuVst9lW
u1Ji4O3q8vUV3yWInxYTAzBCg8fPm5T79FV++19dEDxWoY3PjYMFjIsPLAjqKHUY
fYy82IQvSujuupdVhtlkswuTRtc6PWNA/X39NI0/TjPCzLQJzx0IPN8n5PZYL900
FInZMpujOiou2wnZMODPqLnz5EG/U0ZOcbjJRodWRESrAfNiw3fJKgqZGb5VezxA
CgqYxNXzb36JQGDnyG2VnuOEyk2FSis65yoBWqPouZLtirKrLrMfMgEAAJ98UAuO
Jb3B34gyN+wU6hyEYfqS5n6e7O5iu03u9hRlmIEkfvYsPeMXufYqoSBDYjX3Ve7H
NInchH7vcNGfLlGaO1HbyogF4nRbgPbDxmWNyugFsPWrbZjpY73krBrHnYbnLo2l
c0r08HfZfV5czLJQB4/vB7gKZYtmmk6RE5D3oD9y2hPvdur9STELa7MeXr9vr17Z
Ub+/UYs4rkEoMKpbfxKQzrWOg3lQiXmvX0WFBhnuh+Omx/EzIEeT05228BJyyWqs
tblkeOV6iruWgMvYmh9vShUazLqKC+gjb64CPGlM/qv/3gth6/qAlO1JdKeOcg7l
Qq4yp6va3TaMhf9smkquFhr9KGDeTT8CmOcpcjevBBGdP8pi8+auCQZrHP4B9s+C
hEEZUAs3ZTkxKDIl9AL28V+82O3xnsX7c3WwGu91ncdvH4TNKlMRXBF+7sKI+/Kc
hLj1m7LMg9jrnWRUzRaaUC5kwKgy5QT7/ijJ4kTbLgsHjHLmYwej9jBjbVXtSipj
zb9m6Ya8M4cv0QO5ZpQdaeeoYnM1s5SfFrc2REWRolQgDottdzsL6R3+3TKK3954
FZs0zZhkg6NbKa0zxQ6Ikyk+rggTMjq2vJmBH08Kvmt5usZtqa6ZVwqPYfyMuHmu
s9UDyhUUnMPB5D+euShExWXxFZcdoavBLYIa4QPW1pG9q7ktz05SPS4Qx7bCI6ZT
+S0hpe+oKknV/bNVEOJfBCL5pe5Ba2gTiIkvBVMNUFwJwmLcY45+cqqoEbELIX3U
F1B8m2dnjncpG56dsHc39/bI7/9LR+8BEj/micLOLjV+hGUjhnSWb3xelA5NCE/o
FEuinSksYi+GnNdMMgGdJyC5JerVkp/SGsQItAzRcM1C3UFL8kQCmmiftilEtRjF
TTk8uVb0PZVeAfWQheWJCZM5X8Dv47T96eSidewQoe/afDWf4fijCRP7WZ1ficeQ
QFymtfvMU2cPWTY29fMCKj4WR7v1ThLyRMJ85KQt4CYWkiB2iT3rA0wgRdpfdLxj
iNALyoWeGxEyAR58ClEbVNkIj4D+MPHKzhY817DAS6NwE4arjb8qIzLmU+yHBhjr
7gsu7L3yhLncucwaB/EuZseI8RuuVdUEZNTNQc41H6HCS2ZQfnVfSjvQ+8xvJ3DP
Uf2UtFWgypkIBOp6908lzYSE731UXYLoqZiCRNtceh0ve34ek4SoTOn0HZAIYnT4
PmQO2imZgRTW/XWyQiVxamLj0RfueQhjjz2RQzcsGXL0W8lkcO9a7zT/QKypd2A2
s2/eOpLWTWHIBolQLgLv9bLGU0ELhORjGszZjPRi63mWOT237C+pAEn59w93l33K
kG/11sPm0ILY/0zF2GzZ+ZaJH0VXwyPfNfRB5PU3VTGfcGLOgl1Or3KrjJVdzD+4
z0TgUxuL7qKD6cZCjCHrvP4KV7uTqJgwDYSecI4LoFcJs6D5mKXgr1XmzTsui2Ay
RUqEKL+BNsMlfcHpWob2yZb6ZM7CSJgKAEdxtwl/pXK4cBLTpr9I9Wsu5vNrpFrz
sohnQUszDMuk3yllbU5+fUAbQKPIxZVcQMMrEDVmTYiGRlptEN1KXezTd/A+3gzT
D7evJv4WZyRcujCwLtpcTYkaxrVICi55fhfjN/G4HDUWXL1aq4P4ZiICBrMb/Xc9
1FpxMjOGcdtbimjrBN1aGAZRdy+podhlWy7muADYZaBK9psr36n5geuOHMozLP4h
L8bLtQz5hvHjg1Pvhj5tUStKRAJF4XT9HsZhYMbKOidV01KU/sN6iih42j8r6ulS
twQEdQWfGwP4qfGMJm9n+9IbaQ7uHKlNmiiZ92ucr9YC9T+cmDZocTb6IoVKWThv
akF3r3Kj2E2dxCO36n1JsQEly0/bfe5wF1tE4VoY76j/rA3LDsN3zapqvzX4Juwi
lDZEw3UawrZljQtzKM5l7SbKpEaCg5uxWv7Llyh0ayf6tCYsM/kuKegybRDKMb+v
K4kWvqZD2sLSw6wgLxuaZqNj0RQl5yLHGMNT87Ty0Ht5rrPkdR7O6EhTOP+ucw3e
ap8TMdj93t6IVnZ7NS/HdvnjbkgUoJZ3WWtYDQs0DBsFyA2yuIV4XVtZl+sD++Sc
mHzchI1iI5Ps0fEF0aEQCGw0mzHpa5g05Lp+MC47dM+lyq0AN7KlnBFCZCv31i0N
+Ivd9WdE7j2EyhHNmAPrXN6N53XXYfK9FYLCT2c1QISWQe+6HH42WoCUA17vmgms
M1vzuycEEMlJZjjFJfhXoRxg0MfDQGE7BjZ+qXn24fiaXTZcYzI00NOr/JjqZhAn
xQIOvIM4mHvFAO2Fq6Jf7CtGubpZeCFsXIwt5FyT6R6Ca/hpb7Uz+CcSU2h8thJ1
FfiOH8/2IujzpNTZCS92l/izVIkJAfyk2YId0FT6MatZ++PNbYs/4NWtQPL0ZxOg
0iVHf1F/EhUg/Vw2NrTcEfNQeXBXbozhTJDHIFYcVUzyMbOBgwVpH/2c3wbzAzNc
benRta6lcePdu/8xpMq06oCrZG0ge0OxYNBDqBaZk4Yw/bxNSV5BDH2NpqQNHrQb
Q0G6tVynsi4c72X4e/C8Gro8KJk+Ssjp8ElQu3JWN5cjXIEleTiue1CdeyNqboXO
qMMZ2Kko1KTQdtOuY90f669o0lzdd3nim86T/WVjxvQ7IzjBHz80Ac6AQ/kXnzvW
oCCduRGf/is3u9fTvzechzSiAKIyeKeGKRRcFOXzgrsMWHMibgHTRuamHVILPx1r
SxEK9MJ2YZ/UunI1zixsPNq7Azzm2/97bj40f7I3CgQTtJ4nzLpFizEYWowtvHo5
4sYIYwb2hWNqH6zMRtBy+Gd+TDGF929fh+aBKLDFeMMr1ZwJFFWo6SxvLxWi3RN4
xWYljnPe2xGstoEX5Cm4EYfo4RfP/xzGVPMJ2fHLaW4bg6qoBH/V+Hc6cDY+D2KJ
9NeElJ1iZLZrRt3N3oqDz+oALMQh9g4TVSQt4/Sr1b1mtFjHsJ4PpTjwBND6lwuq
E8HinXcyTo8vNo4QYmW7x3CTS91i5I6GNze1ymqETCfuR01DZ4W8iIrq8nYe606t
dNOLxgPuX7uEW7CZmeVoUvZYkAnU0NmREIJrXICIMgtIjT/X8bxHSac9kYS24byb
A95uHdYU1GZlvpAe8TZF17GeeZQwxlMHRX9XD+JG8egTjGPA1GYtMKTkVmJ8wJrX
uEdeIQrXKRw+Bwet3uKp9lnqC2d7rNy2seJykqb/7fpCZ7fD6eSPt8c1mjj8+h9z
qc8fhEt0YGuNqPHTSlUM+XmBdQhjG/Ua5yCUggLne0EYyhD74GkGrFwlOT48R+Zx
tjwgw4qmqE4N0/lefxySN9EWHolNkRyDPFzM8r87CyNlKM1RsBu1R4tCTItlwzVm
o/WP+8j6GakZLj01FqAFsat/4u4lxJN83t4Ht0BV+aM3+m8XA7rINCK9+wDY6x8V
8LEsbuD7R/aSvw7XnhjJD1/jWdkhQzVmcFX31Z+2u7BjNYYgVHX3VMjJhLzU/P00
SaEwiXNLnYHpD/73dqh5woZdB9tAbrN8pzbGZ5MaCWU2iUM2SdMJ0l7bnOJlH900
U9cP9yr8isQniM6o/3Pkt9nFYQQVcA3Tlric+7voh2t5/o0OwuZfPJordsRsbRaX
Q2DhwtA0nPQ/FwzHVmDk9usw5U7Rre6OJJHXA1en2Py+OShAGIEnq1c452LRWCtf
www8oqNV4KDLfEDGTpdM85jjGR4+0wLvL9GIP0nvUPnUtG1xAZjysTu18476a+r3
6endCtECNn8OyYCLLwzAeKfqgmwvO8QE/Y2n+2VGKoL3l5PUF3BPLgoRYfbXpBsL
Qa7JMWY70nXKVuUwVsRoS/UywHaf7uezrsPsVdfTgTDsh1iQXs7+WmO8WG8/wDdb
aoTB2USJ/X+dVf2+V+PygzBR5JdEGUllmwntPqThaZCyeC2cW+j1LyOksz7631Si
g73wgIrnC0Ck8XhjXyyKM9lNud7hUc4k5mpIyiJiYBuKME5u9chndKD2xgxi37ui
EX63SmMy1duS2Ysa8oRcPWTz8uQUChuRrLPktcaa0NZ4nD8nN1Pa0O6XBXIHDCD/
UdKekr8m1zhZveOxEbcJo4sSayXP8vAoNqOH5kVfy1xKPVtx7wxOxkQFGeO583OE
08+eWEkDAJ4+2x1so0shP19My8PW2DJ4RR89cUsOOLdrHGA8RaViIO/46lYE183E
cEz7ULh1OZxA42pUqnW6sxecM9gpQAJXOxeuVKFFmUPyoW7Gk+QvrENmJuolxb01
4Hi+qTMrD8zPl6vKQYRfjJ72aKfn+46aag7X5xiezIaRHyju27Goip0VcGt/j00o
6AHo5q+Vi7GxFBZpKu3FP1XmC7UbXuIujx3V/peuaxcs/Vulo+qyWdW0TTrrSfjb
Ma29/x0W/BvXhSUp0xG2Q1ER2Fr6EsnUr7pxx9O0dYsiOk7vB/Q1728IIY9dzatU
DF+QEz80zQ2mRuYESETwOd0FuTuG5RKHt9GInaaGrCPr9c47TaCPZSCiK2mHR51g
kfXREEINc1fi+Nf1cOPFQdlF8QW3hhlO4WPIyNwM4laBS6TzYkRyt1mkU3DQDbwQ
tnLqlsqYfGNvw90f16/gMA7cNZGPaMuB8Ng7Ap35KgjRP+vILA+1T5DnZmDCoQLu
3uUFdE/J9L/m0Yz0oWOMxRKUkwij2gYpb6TYMrpcqSo9EyIS7lyJKVlmO61sXiwm
MgCcnUsJUBr0/bUpV/LIhEZb/AQipindTHAk3YoXmewSHdfptoI1TPHgUgrVG67L
2WC8YHdpYRbJGmI/Q3Xt+E14L8KFZlMzJw+FnA1eHcseL8NpeCfUb8HzxIhWmxsA
usl2l++SfOCGF+PSnxCWKM9Y+j4RI4aYw3p9KbCeABRaCGdUlGtkQ389/Llqksc5
SeCcZZhrlmzOVUUXyMKj2cDJB0ITDUDK+bj1QS8AVU3Efp9JAO3x+rMLci98N7wc
YIq2ZEN76cw+XU2Qu4CSua0WiV+hwTS3kN0wsh3cr6yfRrFWMSAUrlGJTlHCTZzR
pyU17AkRTedugnclF33uC66wTZuWuYvD76+JXogV1W+Hms6LjyHA6loDYhvQz4Km
TJtzO0165XkKKh3NmARYyjTp+Mfro/1Ufpf/AWb6iDuSpMJV+7xVJLbphtSneHcu
6Z6bdR4/Wera6Mf1FKBcPPPhhidCTXjXfj0tEqKl8eoJ6z+LEOQssJlOFsN13EZC
FGMGJPq+Ke+rGTZewRpU1j6mV+MYCF4Dtd7HyfCuH1jPNEwOD3h93GQu/90/digB
iruZDGykYnhZA/VZ6b41Baq8dQtey2XqD8DW9LTtH8HPgP8hkcP5lCkEpgWjJIZH
mVG25n4pa8EGZ0Vsv4dIEEt4nDTO4oxepRevWuUKvg02RhLrYT+s1d7Ivq5u3jvf
4YdTUOLrbcRt8NhvJYScI8EuYGYqOqV5Tew86SbEXvB6FRmmKnEeh8vkGBVWfrfl
E1NB7E5pHZrR2Pa5WtriPW+koCIXEruyn0o8F29wve1rsxKnmCzTznKhyjjkiCgu
hYHE6bVSiEVI1HcvRz5TeCHQhdlXU24WYQRI9BXgfn/CrAmiCRfWY3bF7D28+5FQ
VCJwC2ruiNWN6/7Ph6ZnGrn7wTEfBF3Qrha2j8jsvTAYqUcn4CfWbw2F/ULSrcU+
U1YH5zz9/IzXxn5L/n5bndpe+VOPdMeSL4tDFCJiDQI2LQajTsEv0gG7u608qJ7f
cgpnQJKmo0h4JF3e4FW4l1PI6ba13YjELogZZcwkZpxs6kPctv1vL2pDjKr0mV6N
GO9dsmb7yb2ejFeEAH54/1IW7KaALUcJjsIpff8z8q6YUpKykrslVCCxexpvY34F
hB0Wx4A9l3Ed2oYMF4PI916XfXOfGbDYxqR6gLx5aIFoQnbkkKARnMwyVglyeu0F
uNs902pSnhobtDI1YtGBPFwOlnfFsiLXkdj3akbcGQInUR1lFksxjlEI4vuSOAZ2
K1v4jCxW/vIbgyUMchNvL6bLEth316gRSOA3KpZAhhGYfCcXFvwUtIvnAT6imvjI
IwKWBUJlRWq7qEGxz23hPylDn9G9/oc7awvuJm7rhCd2KVYIkmoLazmcc2Y35IOG
MBsoA0joUFCIAQet70/LgWM7+reh/45QM5csmKze+CQSBIjTQCXguziYItYSUe+b
9DTJ8xo/fhjd8IBqkakvmkA/yT0b52tbx7TLREUe3CkEl9wrEGixErDa13cfSlsQ
6kp/ko7RhKGEal1d+aoPFRo6exLs4U5uT4YIXYeXWZgXItNFDgoS+4Pw8zaAgNCG
V36Zj5FvBV8kpIoGOp8+abksAbS/0DV59S2q77i/c3yYohjtUqmvMzluD4tZIxab
jxDTOP10VauKec4rtrAAemvSU1QGilCpNLQLxWdScA/n/nGRDZdqkKB9YoWNkEaU
gz3ow2uhmNVrBpMVzK+Z8lOymQihs9uqno7ua3noU3bW47xlSYGNpQL1K9RdyOcr
vZgyR8nD5DrKDVBZkMuMIM0VFwz/p2DBWxm5VI6mfADBQQJ4PWZVI1g1DRFCfBsK
6Za28Wl5bL//FfTJEWmLe6znfU41mGoYTcqWmREcAiRyDwLabUfE/75seUuXIm8d
RRNPzMeFM1bNFV55HfuQYpZmXtqJnXwM5GGn2sgMtBabjfj3yAYZB1vYWimNCz5H
4oQ4l0polE/Eu4PgZPmgDRyNbOpmm5f+M3SFPxcyoLlyewipbnmBTIBIwSTMP03O
TEVuIvzJpIhIS4z/5z95Xz1o1j0VPOkabT2KYpxeFiU20ztFR6DtrSrVobJ7dk3d
fyL5kqVLa79/GH+/t/cZgZlrrhtEbwYaix3ZAhy1O7pDjB6uMJQCA+5g+Q5W/8VJ
Ig4+ilQl4yuUb+XUVKqna40/r+lzq3HsmG4Ma8ePPyQ8CdmK3pRJ70Xbp3xn2iEI
bmniKCroA1iG/JQJt5cQMZgyMq8lovo3fJ9aHRnRrjH1igge4HNAaLcu+xkD7Y29
7IVzZxck/14r3SKyBHO8Utr4K5E6YwKuT51e5VNzNWIY0yXZJR+QfZfFuxg9phuc
ai6EpWZ9BhgJ2vid8hhEOWGmr0KruSNUsHoo7m0WfJRJSYdD1xrILBTrmfCLxJtc
yVIG/o8ZBUpyK64hSmhtT8LZpuQmN22A2Rzy1JxLd2q9DcuHIba3omZ+vKC9vaVY
9hvhpjbC+nFO7QZifCAhHPydQBQUpIuvVtCLb+x0thKdeLA1MDd+SaABCLsPM0eQ
IKlufeyMfA9HmBSuFc5W+VzpXZtH2QuzmKqe2y6Q+TX2gxcHWblmpVLWVH1xElRH
JPN0NdFva+zBdRO37HmWDh56ojCA0ZByEZGZm2OfS89FhbdehqccpTiw9QwxOwtA
qTCyjbVtgoi/UL2MLN4lNl+sl9R9tmomj2oMsSkvcaq0so7HBhLA1vD6IsZJsSRP
OY0/IlYwrRjHIZ8w/v5l+MqOjJe0ljN51uXAyQSfZssI8AVWmvv8Uva4s0npS+nK
PXbKPQ1+Teradq173TcDt7KLZu0foJLc085v51w5GRKQiizVk9TjGRpF+PxX+aE2
GC+94dRuiOJ14WTxF6o0iMqc+87k6fb+/MUW7J3iAA50GiwugUELCUoweAX1w+5r
MFWVJ6pjRdx9pvwAMk4K3W3mDnaOYELYfPuNFDL9TvzQkU8IVvlusjXXmaFgzOMh
Nu14mA/Y4TcBL/FAsmrl5k0gc5teOVvFuwEFuDyj59RzER+HlZhhC5pZXrGc/Cqe
Ddm2n23zaofu7xgAiWYNjkzS/adcg1j6UG/2LLySgle+drUSfu7XVJFUnQ9TDY5g
+58MS5SEyxzyz7lGt1ChATJA4GSav6mHlhIY09CyL6VrHeGPoyJZOH7BOtEd0lvV
SEkfzqgLs3sVc9Wm+4tu9rbny3eba9DOPuYLiumPntOSBR0AS28lyg+TmGM+lnbS
U/WLfrurxwwSEfSYv5Wt0OJBLWhq+WBIx8qZERNhSWXEGHvy+S2e2kSPSVzqbdV3
GfdYg/8zawe6WzQD5JXdrAoG2kA87CI/LVjatT3dU2hCSGHZpKPAikyEu//cD58d
G3dj3JjbTTHBCZqffkpyTGlL3/H3WCB8Df/zBQX5iwlk0N+XK3W4q3gf/mEsVca5
AJGZ2kZS9oVEYuonp7YBNoHCq8hUlmQ8YOG6PgFGjWFCYCNsyabx1nHRk51O/bgM
iWBgSTjMo1WGO7O+h5ODUM7iVQIx5dzhS+FUtgumOA1UIHr03FyEUKmYrMKUuHjo
uC7aC90GG93HRLC25BVUHBa3v6G7LOxG16NAXJNUdP1i9TRnOGuhZvzJ9LZaS++e
lri4HpxuHpW+sKWbR/yybJIUwTSNiJg4UELiEV1tDyiDy4iPSVXO5LMFEmyeq3QW
n2uM8Dm55Ql7vEj5UAPtghyDUsDT+jhHQbSs0D081xMrEd3vFYODRDw2pFvxgJat
r3wKaumvESbiwF1gVq0SGiSWseft+Z85jWjYJVCZtqMSG4D81Z0Dzr88/CQcGoD9
/aojzo96/OpFM2NYG9pfvFKVfgZOufOYqd8mr3r+iyJgTRHw3yWPluutWUzOd8Gp
wmVjmkpcDTNcmW2wjQ3ocyVzInEyplhgUxhakQhl36XqlxZdSUnEl6aOIWDAhFvl
Vv2bzAsPklhHa1VU/rxl+V7sy7ghdfOzASD0WTnsyZOSLEd/olFHyDluG1vkibMa
YJJ7KETi10DQPyve29LjtFOOYl5R8M0wzD8T45/HY/1TOcZHy9ExhzZcwWkVhoBt
cut96yYQmXHviq+gmG1CWoUAPrxkwc8dwBeAXZtsTToTHXw2S8o8ZkKmhgErCrMd
58pDVRQ0eB3Ly7ppbajNhtadprF8fH8hhE/6wymHEkjAutTjqcplpqLlO2/ez98b
aelT8/Rnl+JYB/SE+CIQChSKa0QR7FeKuX81BmSpFipZ7jqFxFIjP994SQUlqhv9
fO4O8AfJ+7oQAHiPrrOeuoK79H/rDW/NLJa64xhzyx1ausVO6BPLkMQ6z4Td018A
C3uvlaM7d4kf2EK6MRoO3c1iaLD6CQc78l+dCHSZFe3Pik2bjZ8P+XklniVqUMQs
K8LLLq+qqhzxvlys04GH7Y9UQmT/CuNHeYYXo4H0XxTV9WTb9qzUHILQM9BC0a2n
AGjY3dYbIfI9RAME1UQOJwBLyeYX5ZOm69Dezb/XNRU=
`protect end_protected