`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 12752 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/9huKRhRMtvnNqb3Z+UU7TahEoHV+T8U3P3ufru7l1O
3DlgtZzb9QxCbOjthp9+wDkjygH0eUfDrEl1ovhZG63HvizNTnrLsyTy3LzmP4w0
qgqLcNd3d/R6m4hKBKTOswRNOdfGo14Sd/wxm9gRR3dccrHKPlLwv6nONXxZwBpW
EbVQGQWQzJXUF0mxt7mnaifnWkibHVzQKA2WbI7PNnkz5bJhLvKFX/kTYXOnqjml
bA37RaU1ezkyofMIuJFLNTLJvaWsinNAt9dybO1eJl/XkpO/+EBzt9aQan8rbkr/
PxBuJC9Ajp8OGLpuv8j2mBsKXzTxakCP9XsuWsMSqZRAUfdrwjg1EAG1w2cNPbU0
riROYHYvx4Yh3jEkTY5BddsjJkubhyXNbwULxg4IxR4lUqzWjhf8XswQ9uECka1Q
7wlMagMIy7jXULilIPQCs7NJh1WL8vngU6zsN4BE1rezSkx4WljDuJ/5LUsF++/E
YEoKWmhJpEVra0SAaZEu3bbevWoVPxtcBZOPsT2jXgQMSDEWUFWQmYAyLJ+z8npk
6uP/RuAYa0y+Xqf0T4wgEHBrs+a/g6EqdvF7mzWnmW8sejJKn8vhOqfEIVJlV7rT
QsJ6BctyNPWDzEO51SbjzXAjP4yLb3o7u9zluyY7dWht6WkvkL+3olHAYZrC7uSL
qnwOXiY7RWghJmqG8nODIBEUaNdads4G9RqA52Z6cvirtd2DCvn5g1b1Rs0XXEaZ
cnpV/gWJ66XkU/p4Jxg2FrwBBEhgw40GpjC1wa5zPK7h7odkBPqRe/HjQxtgKSNI
sREReyTC2P7/6icpDmPcJI037OFYMjVX1QEAan1yI3rYJPJgS4fxCYmVKr/qEmU0
K+GY/68ZLgrsS3rFRI9IXHHzyi9VMT4EKHp3F5wrwqOBhE6oiKvutvUZxBWYuYlU
0IqCMqA9Q8G/ME/xVSMPpc2uTlei0oZhi3BYaJsXwWeCqVPv/B/oU0YPMnDUZPaF
PLl0g28y17AZ3d/yRO2hFn4ptaTnJNIYB/ePp9RNkfK8F3hAitPDDzyjZoOlnkGn
schE3khPwqGqWQUSYYA8syYKjcyjqgxuEiU0rsaVvvZ8I+HDskEQCorM2P06tXEh
kBL48Y1gnYMBw86tqnDIaH18M8X6Cdx/VFiqL71mHByU4uW90mzAZBhkqNb6qhhC
W8lv7dpTNmmACfPTtodQZzTOYAMyaAx7C918yi8Ox0TBXA6icPM1Vte4Z7JNDQtu
pRiNCQTnjq/moI1TU3H7s4tjsYA7sScmz+7FiXK4dgcutRszeJpedq7khoo+rtoc
smMkVKDd8+7wlMIyy9lKVv7fjzlhTGSPB9Z0z/e5G+kDEK9DLgsFk6M9Pd6F51Qn
+773K51pNW5lVMF+23QLPITjNhJfABfFtkZ3JIRbTYClv43SW9NO+Ug7SqgqZk3p
xZwDGyrIETdXUt7jKVCtf+I9Hshq5Ui0f/OH6mpHJHyphRUbtECHJPh26W+Ug8bB
D+dtYQxsu3SIWoKbpcSO3lArwW+qGZlFVhJkK1JpjYqrLMKGZM0xLrLYj2sHs4Y2
30CK0gQA1Oj/6XLBBfRIlqkGRUPgP7riLNOachhe2szogxp2Y8eXINEbMJNVmVpt
UPIvfAJkQws7tfn88NuCaDOOuyzqgZPSupWWHunF1167VGgTzM57WEkoBP1RaAJh
4zT9W47MCyEo1rOAZGiS6VktV+Uv8A25hYmdXamzpNpvtTEV87uZm6v+vJDaO2gZ
rXZiPmAi2xj1bDRzJYnWfw61cJciriwKE4v0QwooiqA/qmpHU83w2/8qgJBLUHm/
cWS+e2t/RJ4gsz2G3CDjwwtod87iw+QRyG8ZboTioBMpesycbdZDuB3OT5fzfz47
csoskpjnGD/aQVU/DwAAC0UAU37vBayXgQ2ud5dond4WuBydkp+W9TdH34tMklIr
yN9CvG+Og5+biTLU5xn0xvi5rEitD6mu8jVM+E8c1WFExLc7FiqGb0EM1WqxH5k5
DjwmwO9yuLOx3HK0WGf9Ud+b5hgEfuj/nH/BP29WwvJ7thOjBY3bC+uX6boUk/ns
9PKDVnQXu4f6o9aORJ5JSRSlqKyRfc7Ze+Wz8MmYblLRT5F8STakNpULUF2a/uA1
I7fGLgIotiRuesil/agCgixzgsx9efVZ3nbEWlizpU/Hw3R/itR2bw+Hc/Y8G+Py
3FJmIFtt/QtdOSDXgLUZ5w7REZEUvbOGGjrQrXtPltODEBSpPHxwTsa91CY+7YOr
OBn+OhtuqjTm37EGM/ngDwanw0HLALpcP0GYmX/gVBgvAhxDhqv2/A+EhXJ9z05U
pQ4eQcL9nodVZTdmi8kg3q7DreIi9ikvmWRxNb4dbK4Kb2Fk01D8f7NFcc89P3lh
GrvnIcJ1gRUkKMbE+3GKJRcoI3JbQcek80lt8MY291aoKbPcqljkH8ds9L1+ShZ4
0jE58qugJ0jmqL9brKGN3DhOFkSsExSrKu4ohYx7UD35C3M/mqU32Z/2+AEk0zi0
xRLOa6wJefbOgpTMps6JASPoHbaHGG6pTtpKblb9h4TV9VTdApSvcWxZu6nMMb0Y
Vl3wiL/I9j7wUSMSdnbDN223B84cXjpPrS5EgTcUf20TUk7KioLC6CXuhdJMyAez
j7iO17FE5EbeUjYK2lCrhCfd7v/owMeRQuqkzVI5OYDY7aZHFI8J6GGpOGowbR7u
3Jc8uiBmkODR0ycn+OqleSC3sH69+7zClTCOwXoaj8ynQZ12knEOChP/1CAeYpSa
lCZBuqPLp4j5ebM7lpsgE/jk640GAz/T5jjiqDib+4s1q5vVzS5wRmcgRt73UskR
j/gclMPzUGfbCqEYPoeVbEaSPTBO5NsfdjlfGnhm28wxYy3jLNkTId4ivJCr1UnL
+6iMHOBD9p+P1uXrvHgAPvxUYENY13qpArVHf/D7Ln4HR79kEGYpJHqZxGVu6vh0
28CytGgeL5sTLxUIuV9sd4bLAWNf5XTKsdpLDaYxfsgbXgDq1cLgoZdDmp5sCVUD
lm5pGl04R1zFZTVbEepRzaQzIX0f4Hbq/Yz2kIIm0LfbZE/cuYrTGvYue09zrIeS
mzsK/YTwGscWdZbuOKR4mJIh+8iOEQBnynCYE/zEuTQORwmELFPaGhUqT44Q/ef/
vEOfykJ8kLRvfkx1suRSUgUToNkz9bAoVc5LF21OYsBj2UwP8funA+uNQtZpAxrd
yMqXLyHdI16V6/+v/zvulnFtYixLP9W/Rz1GkZlontewUTJkVTAe9us2Qot8ek9r
o3E5+TsrfQNoTaWmXkLlCHY03n+3k2QYBWj5ETn7BRLNokq7UgBvvXanDKfk2H2u
kwjDZ1FIIxbN68eISZo2ukkslbfVh2ywg6i1C4OK3GCZGDKgibF6IpamOSntSECe
8CPBAXCjqYCFAG8zB2CzeHOs/KLhlVjDyP4khM7y2Nb79kS6iAIMYEKMD0EpAXjx
eosozNLoS0PosIIcjcCXoVzrENj0djz3oCJjNdPP7ybtTfr0kMDNAbUvWBlx+Wof
40YBz7kL8JfBWHuyFyGJ++w4F0Hu2VhGvtEK3ORerO2Lc+6WM3LAi0hrUgBag3iw
PRrLAnYxOM9E/8ph/f/DKjKPf/0WSVqrR/6SiSzqeagF59kQgr0+HgFAzoLj8jVU
T7+ML9RDJNmukX9jYX1SIxqL8rS/FoU8GnTNI3YGjg89X6dBQ1vPQukLDu4zJ6lM
0fYaYQ2SrCvT+LgDwJyhje8ml1csTNR9r+VB91ugFgE7Us8IOH+HRx8b52jzM7bv
e+AnkKa4r1cea3691jk0FLFNtsdmdoAkgrEiJopAXj0SeDl3TC2onDDRaqZEyhTD
fXW5KEn7VNFt2aE7M4B6U61rO7FfNfic3FyO49guQ6qBcTwPM7ZHFgdEIUZonQYo
GTTp8gJN3kmVI8+bBdEvPSv/tKqueF9jOgLHfvCnz+czWPvy5fPbRT7BCf6v88Hy
FRFuj7xVtcWBdlFw1FlGpEDyt8yj3bGMu9mh67E4H9P07P6Vv8pbIOuR4aLRAgAv
Q5DqVOYptRU/kLWY2j0vy7PHp1JuxvKzk6vdGnwA/zFiBVNTAtNuVYoGSeJ0VrO0
WG7wjK9LjIaoPPsIgI33Vxsae6/ixDXnKrY1Gn7DSyYoTUVrhajw9R2u6KfBm5Ku
iazDZv1OWA70pMNMFRzvX7LVfA/xH41qxJuld3Zc3cZFRTwZsPlnOWFiwVhsGSaK
rrdx8+cswERi7Vt3vLv3enP200Ljh2mCRZDNdwuVcBXClNH2vxFxmVhfdN5Rj7gW
OBZoTOftaFH+gTtXLof0lbatkOBD1P0CEf8Ks2L1h3x9WJ55iA0xY7b5OEceztsX
g5BvYEMcEQX9XkyrR6h9dBE3y2uakGTNJg7zr9hsUX5G5ifZVHa4R1rd34dCbWn0
R0ucW9/liVbjoPAtcH9EONf+KOPTgMGsQxC5BckPSa2aUFJwL9VuTB8qs4PWm+p5
RIe8uv505xNmuJo2C5ZhbasmtlgHmNqrhTaEshiSGqTLeSO6LVRbfFUqsVzAUd/p
Y2mAckeIHjd0XA37D8NEsn8THdGKFHsB/he543yY82rs2R9qZ6LGyubwdsJzKDQk
D/vlZpjcwK0uTAnQK8pINNb4JecOH9PYWV71t8Z3bPgPSpGI5YFKbAtgFF6s3vn3
xqXCTHMW5MIiiiXDyFrXTuH13a4pwi/qQbwoUXbEECvgguAWJhaDjq9Fg6jVvIh+
38gBx7y53Nqe4+G5CT7M8r7m2emILQlJseltJiyQSWpP0Fh+/wfnowlxlNQu7QPg
ZRvuWGeEblkTnLVfPXjFl++tjFlIhYmxEKe55Drhnn6iLewxXIyfznX4k0JxaYAx
OgrjUS5u8g1pEf6ti9DeXTxpkEVQTjzLuYWW875l1hoj7hh5qRVn+8PtXkppRV/7
CDFzt5eU9x5d5t7/64lkCIsSXX2Cnmq2ap3QmWZE57wAmboHx7LC6dhC6yVsLpyk
Z9iLOkYyAh/1GgvvW3qXah8j73sCvHk6hHOGNh7WxUOQZxgXuEY2as306w8PEohn
e9Lry+VBBqJ2AoSEoyRNNV0YvolZNboTFlkTxeoWwyYnW51jxWJI/Po4dR438bsX
VMUOfnGustsAot2du6M4ERl00MMH8hgnCKNy13rZ0ucnq879WOl6ofRMOuR0eZCx
v79VP9Xyq90AwwAPnYeJNqMuntUIvOQY1gF9BkUGaZwrHlFhM2q87fX4hDlrJC3Z
USEzf2z0lqhOGvAtAl/tFNC9Pqn2iUC2Sme15hbiDlDq9gg3A7gz9CZvlGJwqKt0
KuMVPXg2Gyo+qvRvkOiGMQgDKmUyeDnqa1Tr7sVAZZd96glwn9QquLjhVBEjQ3Ch
duV3iJzI0UCs126ubO6qkE+dp8zWeDx9agecyY/2TsejEnT+TFhiiW3OPjpEwS5G
Q4Xl67svreUl066V6SOSZ9KvYU5XhI4X9FqsHGMQ6VuMR5D+mUDu0oPByW59wAoI
xyoAG+v3fcAJr9kshAntmP5oNDu9hQ4UyyG1FB8WatE0xd/ksZWiYiyti1A5Rdps
b1Yt9lh6V6/5sohiWOmc9Uq36Eirq/BVzzKQxHGfyqT652KpeklF3wpDYi2DvNJ4
C0tkMNTtpkkmqBK8vlQMFofW16E/Z9wFsyYntrd9R5KnVsGUpWlwx6K/0Nfk/Mmi
CaLA6not/BN3UEbAO9MI8GhOGxTYYfMexfZXdbixwqFSgNC8Kt9PqEwQrDCLkZR3
fmNIwfx757GDjN1B8xdDf/1VD7cgGapldMMxv67GGauaIzDcfxIB5YCOdDN8KmS2
LRTZLOP/1srQVrm1+jkS7Y/DNQrfoo1DLZjXvQ49zH3sRqw042CauEpaX0HNQ8Qs
aZilgKz3tM+QqYJyEKp3OcUhSf5QD7NkQJ5ncXDMgUU296uyWgNbz9rHJb1R+Vkw
LjS88dapi/NhyOtjq+jjUvxsAHRHXQJBVKTWHl7q93Vx/q3WNVu4sx6/uUZMTBDh
zswKpAHnq/SrhRJPXl2ZsL1/tb7qk+LgI/BTF1DbhW26Dz3t5c3yDSNSZGCI619k
lpZaLnG7Z3aGgQFfiXHiO66cGStTYnZW7uiBaAbopGZVQmpOpePM5//vg6cGfFK0
ZKs4Gtgu2npi3HJvBCkjxfGbR9Y+EJDs3g/PR9JMLPA8Sy3I7Q9ujPxwLYhWfFAH
Qx9snZKl2aSrUKe3e2yhDONh61SHPgTYR2tWWCUiXnofzyx6xfF6lGEHh4DuLQzz
Ntae0maQ4yriYI+av7QjWlD7+KHgszVKK7XLBg2hRjTStdwRLn9b2m2Wa0oUwf2+
7yPJVD7jd5hvyp3yxj9BMVA6sa9KQU4ElodxDBSXmD5D2mGJwwk+9TvhrfZp5N/8
qz/A91Ysn4oc22ZplYCMwMDunYcYgyM4hr12HWFptDoTohmjd53psRwxxSJsa4IL
BAfOaAGapaXh6zIUB9dbw7akgzmp5X0UxdPiTLOowIY/zRK6BYssZPoqmbrYr164
RuqBQ9CoVP6S/rBLWnoxcYCuJTw8ZOe+/S2x797qN3fEdqI91PIi/+rtYikb9Xnh
jLXQ1hDzEw38LhK6xVAZQRU59JiK6bNcKRj0XzhbcXenxSCb76JhAzeuj8pwrGlQ
cDOTZNibnUVk9AR5Qks/JPzCfoxoisIq2dPyfL0Nxd1Oha23wpue9giTW5Smtjxp
m6PO6CuYDYFnOBamT8bZDXUoX9/OiCPNRZtoDllhBb3MZERfAtbNKbkg3XHiZTS4
bMLQOP2Bth9S4GhQaCdpq6mY/umbxsVCE6pZvDmzWDqHwYVlVWQ+MR1OwEBoQIgz
wG5o7iPPV6LvmtLIqnMjdgqX3OSgTu7ina3/rXW7m92BDOgoL8j9UpcE26Mj4cLj
7AiFf3f2zQBSIWyHzG6+3V5tNbKoEYuqLboL7y3on9hw7N3qpJYCcXavSfCx+dZG
sf0S5i18VoYyA/CQteIlPfqNx1hyuzb9eYSqEFp1R4jGjk/NtWr1gI+JQbXsY963
6c2yM9omkgAeT7vvpDOBFpVUCnNyLTOnz7DsWHjgioVQaTQFEALNEhRe1D4ixwVm
47Rpiniwn7//gOz8zSkdFh6a24zr+hdka5OUa4DRfPB216EyERaIK6RwCe3Z6r2k
5YYm9aUFwkFbm0R+aR/+hEAdMbdrCKN+VQfDk8BqErqvm+5XihE6J/NR2Emcr+tw
jeuEzPEv9e0oCMdZe4Vx4siVf0vV286dtJh/vh6RTUp0k2oKQ7AIMQ6+Z5dBP6U+
+6dX3VjSexBRfNX6OglZEsD5LmTeqqigivosNZNTc36gyYzoUjHyt2XqwiXqYnG7
dw8EffvxW5MtcpqEr1iXdoLAk9nLDHEE51AfvAs1AZ5JmHqQgsDtSwEkrsqj84Td
EQ81mdOl5cBGDFP1njziVmWWSPu4JREDBI07n16mdiA7uirCDtxOqDotIxV+M/EG
VZmdG0dMuba/BTRykOX24OYcPrgPZ/ss8ND2o70KMjMuZdA2w/OaaRT7oNsxw9u/
h6dzokNIMtk9laVZH/W5TC1fWqmBNere6GsrS+DFFEy38FB+kBGeq/lCIe7dEZ0w
iHl4QpSdOqFWNmzLXp6CYgoTthwLELfvbOMuYkALs7Dh806X//nJjxinRCVoCBld
AbsGA7JjzWmHQp9z9ETxzC5AMKuJl4Z015jKu/WthCXffCBdGYbZSa0uet49fq/C
RtNdtsnOZBhtNov/IOLs2pve7Pp17rGuzGRic8cYea3MAEQ/U+blplze9dTwbgxC
dMSRcpSmgx+P64L2jCxEdttdTJ36t8GCxWQrchUpjmZCMVN1NRq4CXc/KIghZK+C
9WGudgJ1LxXL0oki2wZ/C0yEjAWftsHTwXy2cpObIiGkpz4EXfh6dKH5nzlwu7Xt
n+NvX6cEtXmNLu0DsUjNj6oL5dYkmEEIhOw+WDzsQLa+I10st1HdiMRPpOo746en
XU0hFhNXi7oCg+AYX/WGqQPMf9/nZPHtqyNWFyeDq/UvyZK32LLi19WanCFQC2N1
DJ2AnxU7aw5ke7Q+H9WMhW7jnoQ1fumw/VMtyrZgu6PYypu9LJXLcYepQa98ZjXb
xMQ+GIGAycTACYQr15ujgZ1yzJ4zT0twrtbvbG/ZMN8rUkd9PFazIU41AvojrZHN
ZWKUG7DFn8gcWrxvXgi4CJDfkvtLefkxY+OOSffwaukcKX7x3PSpLLWnhG19B0R0
zG78VguJiDnSZ0e4tcrkvnSVFcotEUK6iwcT6HmNs6uKt3D3VIJXmDTk1BuFckFq
sM4YrWcvmUpu0Y87LAkGfZ+B0BUbDOP8RN5oJxKEyyKT8RWyYf7oy6ipcBuPvpsQ
yBLlDhxEeIHVWHH3ApbKheJ0B71/uQRzedgMoYOfEriXU+uzl0Iquygkmh7/NzFN
2j3fzHoj8x4ECwDVADMb7LnvBDmuAljOeLEOvQZAeyZkAKQXpi+Lpr58b7r0flnD
Pc5ArSYjJFTENBmyVOFHMz4eMnytmvLvAyEjmrtsnT0M/GyICfdobqiiv6dxyxz3
m8dyMEzaSYLW0Yi68UXkbNZqjmkwo609fkwTJHpfpJQKl1g06IS6tzyEPSTSiVfJ
uluPKfuEp/eftpSTW4rOVUPNTkRJdL1lWgBh8durH9+NuXcEgWZtGW+A/1zHH7yD
3mYtYM5afWvlJd9MtiJfMQevujPWIPIj/MTMGWoGT4QlK7GLasOO0+wG6HWWvDOF
oUhG1abHa9gNK9TnlrciQXWGVP+cLy4vWk5AncEs+8C3IXHnfEx8XQoIOxpWObol
QrMoIy+HA7zOf+nU7mj2j7FinWiwMenWt7oZwaIy1YayMs8LLCfTpV75tkr2BHpr
d6ol9RqRz4qTKV6Ynldt2z0h8TyCKMNughyC2bbxk/fagOGdxgEF/S+hxZu22tzH
gmAMsWN690BiaV9476RgxsPytxnI9c5D+xzD6sqvJAsRpzLimjT3797ffgbwTEil
9nNsUqRmgaU5MqUAg0taSYu+SR1h2ejCq0IYzrz2ao5IiCJqHiGKn3GfqgrfVTLV
AmtBXyT0By2dxYG+70jMlmF6aJ7X+QbQSygeGUFmnQNEB2YyvTBdpu47DaF2DPh9
Eada039qwvQbauppI3GqVJvlwc0L61OW7vb0e6v69djGutze7eRllw8Gfua0QWFl
aZYOdyHi4syS3A+09ZsOU8cJMTOUEcHNgpxpcMZkn5OMZhWVQrAWmfkMq7k+eDpM
zZPubsjgkKlHcmLmRvL85SgEfhdbIlpVdB6qkvNX9/QPhSnJocUv5PtFhhgt7PRg
es8j09vLbEBr3Fpv6lKXMBeCpz5Z9G6oWSeJOmNx/ba6JZ/Dba0Rkr/VAzMPLqHI
gNLK0FYWldsCoLt79MFOEJb2ebOkZHoHnmfmxxj32iqT3BzvwqqDpG7PgJOm8f8j
A8CR4L+tJTlzOLQs5S3A7Vp6uI2wzddVxxofV0GYRli/xgPiSyt8+iYfxFb3xLFG
sk81TrrE9Bomi9Q19SmYmYbjkh2feXhaQrw+k9BwZJyffNbeONfhKkeyPmwBv3KH
qjwCaUQcbaSgxW76bTHjDdFKpuWknNBx4IPjQRN8iSgb2eFMRy2KwcfnU/n6i2Jm
y8AGh/6XqQw07/yEmLjqcdAxUtkOv0MsDEoKKlYhXgCxdaP4j4hsv966myKCWPAH
aFu8GSx5Ypuw7NkWyaW5CMBm8NP2yHLZJNYGLXxSAsfoR4gO7R8H4kOjHZ42Rdwy
HpHBNDsQF0VbEq/cV9LTNIujPxSwfYOrC4g1NCwdDUHtmZYdsqLHDD7YxJLA4zrb
WFIgXmgwPetrzVwWPbo/LyCyfigQIo1LQym6wGmOnXZhYoFEqnNVGlSj+UGW5Nfi
Ft7EW8Or5vtmWE5KLCWaKHF9AFNDZn23ZOyfEF03MBalhq7h9sRKCXLggkD7wX94
EHxgja6WthH3Bsy0z6FquYxBXyr8AMPIWS8LzOZYpzdM/CZ3Xw2M/h7j2hEov9k/
BxLIJS+WJksui/Qia2y04jLhE3RAzJ8R6Y9v9u2B6stJZxwY6IHtrjoEpAGTSk39
NSEipo2BCHDZalg+V41x5bDUlA2TVbxIsAGYvDP6nUMqt0K7HPfISjAAKuXGr6Is
prmYHfEVtIWVxXbjTeGQcgeTOCuvrk4J9tZqOEw1hBGou52hoOmiepAZ02VZSx64
J58sF6F3RTStdAbpkdcemknY5ANNaXM7fEwDrrN+k+2GQ5dLG1yceveMINWMrEJc
l1PqYfG/m/bCfz0/SXnOddUDK/sRqwed1904rKfeY1mvVqnDa50DFHElmZXhP6H0
aq4Ab1TSt83W+N8+Feq40iDRup0pIgYIKniUUZzsmrPFToqq5rcmb2Z+paouBVtn
ZRU9rD0gkECVFVff0Y4wDEXHxvwG8JkwCQhz40M1Of6yEG30i7kirRrmjaYm5Svn
fM+hsaKka0GaJJm4jV/mRkJR0RsG2s6EjE1jp1JnUrjsQtAbcgNZ2fZqzujcBbeO
1x6v42aF0YcRxx4NU3ITWDf2b6YBoBnb8lrjgH7yYKUC6MzPlso/xbZ03Jyr9Isp
5uPVsuhG6HLeAGINfLpeYCZuUmWTQOKFCuep5s/v7B4iCS54u3CKflryrnWnRvZJ
y7uVmEMBRpB7k8WqXHaIktQ5MIdXvYXTW2pasbC8yTa1lVpqUUUjXtE6crN6zan1
rSFmx/NV7TjlZkUoiNrReiEnPRcZGVgymrKifqRmbjgdNAlBvU9teJblvLnn6Wrb
VtUbgq2vkaFTDSZFdTVfKW28eOxQscEMemqV8017gwfUvmNBB/Fok010RLsun+0A
soA3TRmPN4zn5mCdXuHSekINWM9aBJardVTs20QuDngP6LRmN6ls0RYErdgsrPrS
IjdeVbNx5DH8F2c+dw09xJ8n3ALaACDEsnesD8lXo6UAlrV5WT3fbghtEAd2H380
n9mDiYyLT4xG5yMpupI0tUtZB0QCtHYzKlptlvtrTl2HU5vw0EYF9cqnOVE30jkk
WuyIpvI+Qs0Cfq4VKofLLhiXpkaJj7gN63aq84/pJQif67wmf/PrprWIwNr2LEyL
2kGsMoJxjSJyLtu8xUF/WmEuFsVweWlEI4m8ZQmqWWZOTQlUi28oCw9wFV9bLcif
9iaEMy2uJTzG0AA/MTfHgZbgOTSH9t9d6SkxBsMKP3/c1Q4TxTa86iIZa99OTpBB
ndVOrFN/D/rS18WHN8Iqb9fS9Vhh0QWGszJRNqKsK4oWuuVGooHXMKcrAdbHAvjH
ijwY+hsjSFaiaCPFRUTls5LbHoz2KVEBN/Ck5HoBEeLu1zjcpB8WwI8szCoRLAIy
lPBYveiGHITZ53kutC8A3j3dZ+nqp9C10DfvO7qSHnXkClXosMiY9w+ovdj1FN0W
WjBqLlTzB/XwaZ7ghvF8nQhnk2VbkIy5XM0wakzFcNb0F1JhM1dgoU9zgDlAqp0c
nRXXr0N1OerkMpRztbEVZgxDlVjlCr4M6x19ib+cFjMJ3abuDP1PXti711GIcd33
mwXpz7hCUizbvHIcMGpZw5WRfx+0odKREEycyp9Q7ItrUPBHGzXQCP102L2oQMtq
8pHRdv9irRmKRZ6XilOoYC8YkKU4Flsx8iEHIwu30FTGln+JS+nCYMEEcFhzKOcZ
zjpLKDPtgjxmwkzYiusY/DYSWGVEnDmucSatDmlazfXk0qkpf7FTM490//sduxI9
gHNHchtWXtIGpNqjzSAZy5U1zWjPLqlbOCa2Qe6Bf5roDn+pzPqCDXowLSrQaa/G
F6Xekjt3DjaNcg8m7Ew5eFnjPcvhOWTtrnIUFF59HuhFyo//Y2Nx3BU3NMdI6kU2
800PLvtB4MZX6AAv6XFHovlKOFMStTbdruon2tldRqr+z8jwybPX6cHyM96BPk1n
opwYsTLtUN+u9yrMobUyXgLXiZ3eh9ZNAFs9aqNyouPwysNCtijsO2WvEcmov1Mf
8UnC7FhN+frccI6Vk34au+DvZCkwq+RVAIajFszcctuHxgMHrhydP84l4W6ZO3if
2Vww4Ly8P7t+AMR8rQvsW4Gc+JNre5fvinJgbc7Xr9G3Pw9/gr2pZ7FjoykiK2/y
UHX75F4FUmXL8WlyIgEBFpM44l4WJfFXTKpBxfr/aR+b9MmHjrsq6ITCQrF+Hoe7
bmFvSFBs+4xE6BYeH9GZEpQf9wWMdiYE48PPqUdlyrV9vW/o2/2qM3d6H+75n24g
P1H+dcLuTvLj3ALEA39rQ9bEDE3si+JA6zcPDwixIODI4urpmRBXmnJzO5rLIn/8
/JnLH57uvWa0F5hTYos4WQr3ftLTmt8S148MASbTcYlI/6QyVHvUFw18CNWL3C5g
IqZCtq/yGynxMBPvFhu1WjFp46l89Pwbv8999QKXO/L4AePxvoZMutJ5RvxWPSwi
I537YoQXAnaa14+E5bzS4a2AY6k6OpsWmpk6rGdxRYG3UHwgoMNCVrNreD5Tz63n
MCkgD9v+XQIziESCHay4nmKxcR3Hs19qGt3cKGE0EoytMIkIOhnV815WLPtrcwIH
sIMxtsXin7MvLrFnNsYDkMfbWJtfMmxZVAsSvx6yNDZFwPt2aomIjTPcr7yUUbxq
JVUTe9h+RpUIxyUIJsL/5z+pECYhOYllE/i25cytyk1JXSMxB6am2Bt1rxT1sUKe
zO7JBqtunTx3A8n4LMQVV9Yk32rjKY23WZ3vd3SK9z0qUJEdZKm4U5a/gyhXWl87
8PDZolrzMNFD/iKkkOUUAAcwfT3DR3IkQSloftayn2loj/mjEeN3k7NiDD00A5kr
9Z3LeBwBCNJEeT9fJi5hWjmeCZ9Cv21xVzAIlD3flZR7OkCb5NNEMCfprpcVmsmc
RhkPltzT1ChBBJ1yjWazZ4ONrEv4iQgEWnJZtcErtRijx0WQUAgwm5ZLTsgj33Qp
wzzXJed209tcZQ8Qvz1kWVp1vt6Svc+BDAOZRTsPbBD1iLeDGaSI4fALFzV2zH9O
1dIFn7eayC7UUgFgTotBbSRyTXIo/VREJ0al7QLPe0UXa9S7mntl4shTnXrM/sp7
+xFjDwQhCOHxglNUHL7tSlVYeG+535FIOTJouCiDcH9kQYoPjg1X35UVVAIPAGMs
gpzHyQCmAQakBT8sfczctcwd1syWD11yiJtMHTS6PN1kOAvmh3qL3KgomYptTByZ
/oV9t3erF+bjHzhOZ9noUH9pBXEy+rjCBDEZATxGXU7Q+iTqXO3oQ3RO3XHF1NKg
9f3JOt21mGH2Y51BmCw4lJ1jg9jRoPdvBVrjMC/84tcfpGDU6AOlEah3QIcWUVAG
RMWzM68ayAbeiAeApuLPwb3u6pve6l777Df8j2D8NPOY8FUR01F+MmiPnUnuE5uH
KcVswPjXn6y9/jOwq20yFE8Wz/fhCIiqU2dLkXVO0rZVUVasG4+fdyWSsqi1XYzh
qKJQcliECvVxMahroI61JAQrLCS7uUMSqBTRkOX71ny1xdnSIg9bOuQXUlDbpvwc
8xFg5z187hG39IPFgPgwdd+Oi2icd9hN8O4i9Op4vNKv5KQl3X66BpLl7Ro565pv
Q+i6dYjYElQNbtqVzii/TVJZBh54Y/wQlFG1ERlDnqrLTP+zO45rVkKkeNeB7yXp
vR/oRhWe1c0DcyBTFvRsSXZzx40kwkhyGZ4XtP8m0kMKRTOBULYyLmim35tWAWOY
FxVdJdMImWxQDQV7iVbyjRHO/B5N7wuvHaqwgWYOFvbEc571sU+fp9VOU5ql4C4E
IQNPjPrbxd8Bb9E1NvJv6a7kXdq9M+mYvmKVLhdMMVU14p2P4MS7vsZ54SNtHbth
3z9wcEMjSbWCk9V6vW9MSXsVjV2zzftlGzayfuZh+F8xGG3dF8t0fXEOUabwhT7R
EeBXImzJ9PTmodr9O0eMFBmh2FNORKEiRPd3FSB80pswVYZscUDHIE4HxVDtcMph
k5YWiic/f6TBVcQ9kjzDzGdbafuQhcL/aYed4bjvIqoGRxnbVs7ae3b8pj+cqIG3
zk0md2SAZrVXRPS+ZRY+VRP7bSUSFJkCJTT9MNWnRn/OoBsrZ1PANMsXmZhTZH5c
njSbjmzcXxLJ9Zn/JVg+OAmDJXtYnqwIrGpjuoVUzXb+IdEFwifQbsGWlO3aoMv7
nqc6Zchfv/20B4mb7G774tfJdcNSOTtjpXt+x6FZI95EI7h+AYViYVtPRpvSfr7Z
cKXTwW+Xh1+arL5DV5AAHZis1kOQgpbbe1sOmTirehQ0EmCRftB+WH3zZyOiKmHl
8wypkeqzPmdWBBWklnmaR971VVPdAHok6P72aLctOUP46nAazraGNVsBWZSRsGbn
JtcP9+Nw8eXfHh8UH2F3i+NSyJ4xW7Zoi+E1Ntdt6qohrxccaPhSvpnTmc5qhSZw
0pK8hT5+ha4d2SoGCRExdcEiyQnL31ZRbBRv/hPM0dABlsWyzJaUAvU2y7O1gh+J
D3t84o+W0eCovxen74kakmCAihtax1nwPGVSFQJ4Z4pWxFZ1XuSTb0T1hyFHa+mz
KZKnPDgULGHgNt183DYPmMYLZOG9hol/T9cHJv/k8iDX0P4OEezRtUtPZ6vw0HAm
1LWuK/2DwbQARJEooxkASOMtAr14w2gpqBB9LndJefZolIhR0gg+fwaDLv+BlBbR
6CqK7FXpxaSEkMKmCJ4xbQOW3oSdicjG+Ly27tqsmFsSfiPjkzF1eSvQ8e30Mh55
q1kiqH0rZ9WGHUaL23LBEvB6AtVMDo/dsp4snoa6QhrOadhgMEpDmSeYCmjsjomp
1AGUH0O1Ieb7LVio45rdDpBNXsCfPb6CjwzcQRqmwnNfEdaMjEjcOS6a7GIXNzYM
vYc+N4rRB0saGGz/IedNCCgbLgUNL4pQ4IuAmZ2U6xPUS3jkAfNFYjKLK/VUwmaf
azTzbX8EHYT29ndvsxTb+i9GVh2aSUFhzbFIQf+Wvty3kGRmfBRD8wevV/XDDS9o
ZiCc49lBwNshdOFOVdavD9xhYtcMsri4Ewfb6Hk0TV1/VjgJdW8oaKYTmTW7Ywy2
sQfLUKyrw9qsfkX3JkQxDzd6tw8bdRP0pjjaJZ3tZ1Nq900IDniCsn3+0jEIHtOz
HI5StTDlGcI1tGQCTqE77FFvdcvLur0giMk8Nc6cRSrbj9/dntZZtTAEpEL80Do0
eCL2fggecUk5W1e0KYB1DccWS8opVCn/dc5AR9qw/GlbmDD+v0pKiby0nOzsMRYj
sAA6G624mZ2e/qbcY4kE8Miw8mW5KMSAQWgbD0//kNXevQi+jsxVGAwkEqdUqKfg
ABImbJb0snRMbpI3rrV0cu4FkeQNaaExcccAfhBAtUZp3wG5hjZSG45BEvJpQcV0
2Ntp7qcmUdAorpts85xQsHBw19SxuS/h39H0CZ0KFeX3hmhts0RgWnmTPdgim6Lh
HfjHxQIYBybYNR1siOJLMxcD2sN/lRLa3PJm9JlHMNeylcsa5vf7FdzFlyGx1HgG
KNN4h8NH99vekNm54z/bLn+goSC32dSDqBwri4S98I+bXr5kev6gjU60duMSPMh0
yPYL8Y7QzD8/B1k4sMA9U3ZmCgYX9XOODDNaOEspr+ye73Rqp/4dsyz/tlJ7L4jM
3RXXuWLLI0LaVH1Kmu9vko3Uk8aL6qpC8h0wJaNWmCFvHNBaddD8NLpEuUkSPuwV
AESsPJ5kgRvZUHrjtq29r/8fhUoY2EhUVAELwWnYP94ckP/bLmn0R0gHTvllvqN8
MKBGDaFr9zN7epY3Omz60dZsIO5njuXu2mkNO4zBlKb+/fhrCORNZCtvrYW4sw9G
7y7mUBMtHidIhdglBaFJFAyMhHNIeavNRw4ulsMIXMjguSkpDUobmAoqgPq7ZZNh
nJ8VU0FMhG9VYD7s2X3ZT0aP8kfo/EX+fZt76orp8RCy7tlWL9OTuAJwjhVguuzf
SApKizsmXsLRePVWavkvwUTSGwpBdUphPhwDTe3AyGmWlQpASNHT+JxAgSAtdveu
6dJI/9bVnJ4m75SDmB1JRlGUa7KmOoQm862eNDc7EaxmjQGMC3Jf4YoJ/CcODNu3
G+mEU2Wz2ltyjwYpR0l+7YRVzrXsPEkZhlqm3e8JxI0y6eNGhCoRP3VMWuHMoUas
ZWdwdXpfGbzJHM0LbVbneAaTGPy0d2Q6GNcXqNeLEKPfU6V/qdj+uVqpTy4j/Edm
YWN9G95JLWnU/95jnW3CcL8b8UIm4PzP6vTq+IhCDy2j6w9yGfN4OHGSVD5BkrFY
aYTvV0akxSxcDEw2kvXYZzrPbGZ3fYEOL7RzWXbiE8M7SYys2ltRl4Sks2Y3YqIc
uDVC48mF8VU01LjS2R4dtZao6bBKy3tChrT8QMn1bdybtO6zgqyv0Eum+DHE0186
YW6fdI9IqzsLc7DivYlWDfGnthZNlEUPAa9xKBxYxdWOOUW+lDQwksbTboyLB7ZG
lu4S2OAcElsUWDcg4jugQTGyi3ESLNV6j5fhlOY+7fCnuSJjSzgLfqNuvfl2ZS0T
QregbxM4Tl/vhyd7lECyQW8e4rtWfA+FNz+l2nLPC+HGHJII1heBdSAuYWlLcYnG
ybPxnOajTYEZSVPmxdRTpPNz0FXcOohDNSKSop4/xirV2OW9zJWM3QAf4aJ1wdeV
wwS1E7UrOsezrRhM5dRMllCfeghnXdOCxRaK5gbvXgiuqb4kmLYksEzmf4FhlaDK
2oBbpr155/1tUrec8w0hO46p3ZIsnr2Ol1FdMG8vzKZj6DcmTvpWSZVPiAcsDyIY
nGl+S3t6Rgjl3dvkdw8d09OGm84ED7SvGU5Ql8FWwzTyqHr86XwogleovZCuP0/q
sQUrSxAuxZjpGvX1y74PhZOm2SxmM3MsyH3rG7aItp0=
`protect end_protected