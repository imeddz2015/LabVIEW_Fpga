`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 672 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/59UwEX+aE7FohaWu0/8IpTj7mav863zUNIsgIH2BWb
Uw34kZl5aMhQsSK68elNYGdHF2f9w9SHbeqxdIQlC6wOPXgxrOV96INP1Cv7nDv8
NftU1zrGwP0BJbKLPXpm7vszusvHROnPdbv9gRztTz+dL+GRs76kjxnmC9X8UAsn
FEexjWNq4qi8/T6AhkPRnnXklp6BMgExhbZy8+wOXfv7Ss7CpMXm2YksGP/H1tIF
dfBHn8tl7cUsppQ0jghOTosqIunWxs7yxkXyuatdXjzKFY/CQGijlhGlunc1vOnE
VwvzF6uEPm6arBb6HBfBjuRyfXPQPYnjk+4pOGy/x6nps/TC0fhnBbmQJXWiMhG0
nxyF7P6iUErnBmwiSZP5eWjuEe7x7O04E5JVOJsOA+qiBV6E3yCzwd440GqjzYMQ
/1Yr7v6hwdv83JwEee58j+CxkFVzC1a7GACVTcveR7ZsbPcXNFaSDgRSrvt5Vck0
OS6Cacyn+xxwm0tQZoo+f5xVynz8RU4eqTfBqNSCjahN0zhQjbci0l71IQKQW0rU
Vo6ZQbpxLZSutDuu+tQ3hFuLINrdAUAzQVt0mTy2Iz3q3K1pUQ/grhNOpxFpGym3
VuNT/TC1xRjwPEluL8icDaTJoNnT41qyy6BqP37J9Dw6MqMVWm4u1ugi8cyz8WIf
bruyUzMlXJ3FhIlhTyZb56mXUNsW2TJEL1B1WVF6VN0rNraN6TanuutmzymiGEXe
5dgPGAu3psx6VGHCwdeXjSRpBcmlNEmo/z4203qjY6/l44lOo/ajGpTplARHlWKk
dZqLiqugtlGltRPvu5df+kaveOsj9KRRbMrJRxWB0uASXo3ZNjrOMFbIC6u4P+Ow
`protect end_protected