`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 17648 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/9huKRhRMtvnNqb3Z+UU7TahEoHV+T8U3P3ufru7l1O
3DlgtZzb9QxCbOjthp9+wDkjygH0eUfDrEl1ovhZG63gz3sDLQL57y2AJa3NOe4o
Uut6fRNTWYHn5OENSfhnnhvB7Zx1OKiyvqNhBENS3D8iFTdP6BDkAxaUWg8xGcKJ
JXYQgzBd/2VVMh5/ItMtSHSiUCSXF+PiKdyYk6qfURTnXnzm5EWcNzTXsCLZMwqq
pP29OsW2+R2G6SGOdGoD7ect9Pz+WsXfC+Yp1a149ZXeSC+8HMZbwi+MIcM/xVbP
cvL+7bVys9GlUNk10PQLaiIaITHXkxLxCyCVK8MsWipNZuF4bs4+HWxHD9gYIq/9
aWaz0ePuhhItybE9vbQAUnbKGUsseoFCoXO1p3Rba2WNOzrJulMDCj68200hhAh0
tZHf93WiAp98jXv80Hy0lfE06J9jREDhnV+Z8H9uFLMxiGHBmEhyG7NpTdh0n6ix
F2FQHTOV8A2mgpSR4jS4vOlJOGRFXdkk/Kl7R2NOfEK480ITYfABwIdq9gXAkl+P
ZRaDBwddQ2Hd+LwlmIVQ+T2Zafg4sP0xC5LtDUIaq8+w2DTyYWFBqL/6Jh5+yFbH
j9UpeNUljZHdb774Q8u0Xl+TEzJbs/TpgV6vU0Tl20S7IkR9Nk3JCPhhoBFHCmL+
4oG0o8FbByQ6FoZZ2E4tNF92972N9xxNBq3Nn0139GxSkJB6yDcAxbLeL85Yb5xu
oY9Poh7haefG/z6MALgdmcSye40ZXvrUKiIve6/WaUlFsP6T/iaJUw42hpI640rb
4myvQGcdz5clcVJvAgMGLNVuzptP27TwOqKwGck09VYKHoTndonFR7VbK7l/CJZh
mITs9zLAhyrIADt+bNQMn1Iw7iCOapLUaCgnSVCCsc2vGpLKC6m7g44Paj+WCQQp
EYF/B8xkdKuTnn7dzWue4lkV4K0XVa5Jmi6poWzFYhU/CnZ7BbcAz3hzNg48W7Gn
bu/sRwkjMLIO1UO9rZzwwNOp+Ou4QZ3psJFze3ftm6OsxfwblXXjsB2VsVqP7ZKy
qX8qfTORQSS2CfSPmqT9LFK0x2hsjQVbgB1QOojuzJ/G0O6QmUBLj0Vpj6NiY+Kn
ujJxty1rw2qDH2uS2Iljk+w3DXCa9F6QWh7nCAHkNpI/hzyC8Fr3F+lIcl+F8cL2
trPxS9QNZyLlErCWz4qKuMxHHHoXwibsTIJ0e05J8D+nwnlblgJNifoBq6joEUG3
xXcPVBCHtrdkOIhXHjioFehdElIiagHPXOD8m3SRfwYuQe7pYc5/8hQdH2ssI1rF
Oea3qzI5wk+/igS1uxRjpQtM1plyPan2udI/nTKpy/HcU6/f1mDynvi0DKuVA2tT
txLlkOEAbO5S/pXz9VFAqtrny08b33vITBvlaADdRV3du3KPOes4za7IruK5GLWh
YZh5DQjXehVnyGukHnPgSXNAQIKCC66Xz2lmyLTmUGkFn2nKH2iBlYgXi/w5557A
o37YZHiYH19/JBOOj9E+wZrijdaMWhfwBapqZdoGIK5o2i8Er5YEq0yjRGi38krT
TkcIzTcGrjQJQochRYZ9en+jz/mLE/+GqlIkuK5kUtfj6HzK9E+Z2loTsSMNsXyQ
/Cjq8yf+kTEr3RewXHlhPQDFhkg+a6tjMs72oAWjpOA+vX0AHYoUKqO70j1xbwAS
I3Hh3p8gbB3i9FFkrP9CvqW8U8xaLwG5+H6jQNrxgiwpX1SY3uidbAZORrSo+eR/
x1X7Wt3oTIbxRqISbC2DiC9OLee/8ALg5le0qbJO/td2+D7vOKwtV+UHbh6zoSlY
cnkBU2iPzwuXWASK/mShTc9PUzKBbVoKzYMWBCnIhBqT2+CjZdnaVOcLa+5hshCA
HxSW0QyX133V9kpn/12JKi8afnw35VKDxwJumx5Kl+zKCt5f1R77elIoOPU9iSlB
+aBICqQtu3jNzEnslIKE+aDCXi7Sxx5sXuHNKuDsjJ7vvgkml88IInkWlG7otvxM
XOmh2aMFYzWAzrioAz92D/dwWj7TAv5ZavceyB1p+9qzcXb3rCd23sq+dlBAuUeO
92LdvsDBBJ/9nwm0yxvG4Fzt9Q4mfeyV0H+AJcrKm99ohG7pzpcIkGttJef1Bscy
BK3Y7PNslusjaQXButDWTCsIwkVJU2GzjmOe+0MRg2Vv6eg3iMaZ8MXIal+cPpsY
peJyJjMGRUypy4wXyOmsT5dIciFcuRFnMmSlq/B5NEDcNQMOSnVYASlv0I21liFi
NabfoXA9DiJcU81bYDXXXy6rZHWEhm6QYXnH4apk8OMY4ri0a9bVl92um7jx+R+v
NegsTIzNfVlZSZSm6l3/V1z/9zVoxV0aJHCzt7tigKSaVJWWWx0qd5JNkU2Fa9Gc
7sJ+JE1nw+MLSwDJoySnC6K0q7sG8gHKPY0uWWM/1Rgf5WT8SV+t3WdBM7odA0Qo
IqMrCImSMCKj8nTaDXvRTE8gd8sW9Gdng3s4TGJh6Qxn1NK6ZlBG+jFN3lvZo9gq
MMeeXwc9CPH3qFyQRdYG5q85Xk6PurN97b/SfMsNE2UsCK2GqTUWbLFje1QHfpXN
0626+6q99zECayA1fuQhG2Awh42Vk0zIZs+2wVFhcWuhYcWf7wp0yfZSsCUW7nBh
jP70OYEfi7p8ZTbMuYMaC2dK5izbyKHOu5dQTGcW3ZA8fpNeqGT6vHtoDRSw+dOy
XaCSKs13PGLNOgtq7buoFByfdpt/0nC9DxBH/3+2EoWz+gI/eu9i2dgTPbi3d5Ol
G1YBtHN3OwlTf/rSNBepu9kilmkNE9KE7tZga7Ft3Ie+buqydS0Q5T8w1Kym3AuX
5P3/nh2z7deB/oc9A1fjVBTzMazsYYfsBufvUSeQgzc71hXnytkssArz8QyTXjmo
VtvGYCixAqGBfpkhNyPO2ofJblqOQXojm6Qth3APmHC9M1iVv5uWJ7hXFbmYAtAY
ofSr0ooZA8VzEDqC0Aat0kj9hpOUJcT1Cv6X6ER7qnse+vKLH3amj7FfI1qeUL89
FhDwGXyWjW9pY0ucM6gdi2PqdUBfwLTKn9ebsARKXVE3yYRWsQYzYjswDZdkY/fi
GLRaCwP/Hku79WIjb+BU611B9RJdYaJ4WKGTVae5xhgysDeLpmub8MM/aO2IOONu
gwadj1/LWUoeRXDnD668dvLw41OhWQvccek19a/faNIzQtB5jKGLyelNe/bGFY/P
Vu0lxaPSpPoTgm23hsKRqgOhneMM11oGSqVLZGLZD9m5Y/D4Lmx9NBfOpwYAozBq
kNeTTlOA7AUM5ZA3FVdYTE5TYb90OxqzSTpil5H9+AHyZ3lk4IMVNfVNc/kE8Nx4
JPku38e7tP18V2RmolNdctw7V7ZpVMcZYVbLzfb6KksQdR0QFY6jlt7aJEDTDW0z
Xrq8ZuWJihJyceHeHLkoOXl09gNhI1f81PA1d9DAfpNe9e+Of2O6btQBR2RsXw+V
J2wFkYDhatxoGyItjR1zTbRy+3QK5hrcZl5zFjzFBmVJsbWu3BY5BN3+E1EC+rcQ
evvu9Bba6YiDi4W0VPbUdKRSH4OJqu4T1wOj6pFTWhxZqMuBfLvlxY1YQCPOBjgx
mNq5Qos1RaA3ijiBEWt3sAMiOawRgyjxWPNsiqWYjol5dl+dO8ODxTwZBBLlYE02
vsv7+LmFHO1gjnHBS7CqNgN4ttNHjsr1oz4/n9162QIR9FEgESuraYIxHMOKWztx
4D7THx/q/Kzbix85Xykeq0JoXHasp+jhvZ1GOIKikc8uydMOuD4FZT/spX7SnSkl
yLXFYNVbvAhYR3sbrTfXSCSJwtY2YofsSwpU1S7G7yjHlY4M/ILPDwKjEcanHbXX
R3EEVU4PQ+jDnJ6vlsg47B5/Khk8qGfKSNzpuze6LwbRm7s2CEdpjJJyC3om9Dlk
ORFO1f8Gqa/7HT0b/wfrU+mm/ToRhLknW63+KmQ+28k+i7BUgR1RyT6wDmrP/Pw8
rFmzcH1Wk6CJJOxzTgbbbTwyYO6agbF0h1G95LYU99yg+5/Yydf6Z0SxcLbdR+qq
9Dz2+sAt5IhWdnX9ypPyuJIlGjYPw0WaY0rGK74Z/dJ3bFq44z72BRRPDZ5Mds5T
P7DO/ZmFPA3V9np/crtner05uMT2b1Zyc9pPetIFHMekHvdUjAR//RI/c6gG8tk7
yP1nHWrSWuBdHHVPVQDgd8KnpUhAuR1PRSjUtY/++ukYmkmBwLfLOKcyB0ch2krk
ZUVIve37jvV2EOSH5jWMaGjnbc3tdgNfONc6cKv4gW5BZJTgclmUawrX9yC4VL4z
YN9HTdhIeQsVFgKY1UYk+zCdlbRZ9IL+zunwhYsvw50Iu4AE+pgYcd9XdSP6djaz
KBAmsT/U/1sFiosNBRM72otpQ1MAlI2aLB3dyX5ePpqQyatg7usMFz8aSBjS9eq8
Iv302b5zhfsogVBMYP6JZCFJjWW4mrBs402qTDjn7ghCJWYHFdHtw8tVJyO1Ay+r
1iKTVWoYS+PbY+ycgAzd2vUIUgYfLvRO9l+vI4f9MkxmbjDnk/hXhnLgG1Rj8+pD
sjYMpUfeHx05VJlqDH914PGyIDog8+CYlvB7FgBrPibQttc2xtqu1Iow9MIHbJ4/
ZhQ5+zlpsFU5Zgm9e464P2157du7ktdYJBrzfDLEBkt7TCeQg1lWwW36reywAy7+
5DZV7nJmsSeG+2ZrP+z3d9P27g9pQaR2/Taffto/1lwModuKuduL0zV1sUSV8lmE
BUuwCjRTW4Up88avr6mGxriZ36LB07L26wCQfQMky7DI9BjDWiJ4LbhjUd2lZw5v
LVsoRfaYyxmkXXh3ZHTaOeoOOMmEOEJeO4s/y5OyBQ7OqUJFbHxi0rk2+LqfqY8K
8YgRvVTT8Ta6981u4zuCe5fs8Uki+da4dXrVyNJpz98E+Fu1Z23/JMHaRLNYRYDx
Z1zzTshmH5ybEAna4F79AckX4iXHJYOd0Mn0+EvEFg7IPokxDsCzG/IGbTqXTF4V
7/Mwrd/NIuSFRM7+TSRTEHCInGTO7lazRiZzQtN2gnzjT+lrNGIQplaJbh3DqNzG
8qLTSUUE2TnDxoDOkcz3RIONpX+L4Qpc3p0gSClafK82SNis0jB5X0du43bTrz47
dHfb4AWLGNSFX41cu5li3BiQbmyhl9HY/wIsqwF+t5g9y/eCQae4DMDp1+rHHSlF
mRPh3is1ZlSA8IYJn6iSz7vNLKcoxpt7/QmOtyvUrM4EWNf1xuwMbeTqUIda4JNo
Q3WT/10MdxVNhSTiy+cmDFnUfcBRkxGoBY3E7qaaj5I2uBfN1ZNGe9qa5wC8yQcL
NmeiQQJAmszBWaVMaWYNfiamVZuzDc1tYOwWh7iXjfx2Q2/36cp5/3ZhF7Lakyjl
2I4S6be+b+dHsnSjlDtjUEdc040ws0qxWxOINrfwBTG0O2Puq7v8wzg1FQ08Pb2z
wpB9x9QZPBytHT72P90/oMPUe0+MDRZPPYQ2L2tSSMRJHVZAl7bw6lRk51M2HCB4
YlTTJ/qXLYi+dfgXQSoTM2VBPArfHiN1dCgSONJNtVLc+mp39cuJXjGt2oqFwtpY
N1vrXoPH+g6n3l2JezRBAj4RlXbCniDwF105UNvoNMcA+ATpG9WGtvU6dWV+6Akx
ZTiKXf7fWSjNU/N/EWG02+8kyxP5F1I67BC0xlZqvWYcCEe3doCkh9kQUnrco/Zd
EIY8ztJ+Vxp3zTHUg7UOqLBQNCcMj/hsz6RU5cfA+feNnm8XZPt7v3+Gj+xy2apr
HkBv4gjhTqHtgCP212lsfbBk29P8CERrhYVelFK1xaUtVzjl3huh3644uNeT6bL4
nNi3TaEXzqOWnHn0RsPLm+aJR6mt275aDNUm8gwefYtcFkiEYI8llMVkibLhS9FP
twGfbNJpolHgrJFYoeoqmL3cxBwkaxUkL2OiN8CSN70X7TKMvh1mKmCde/zRDGJC
/ahqOsOFY2e1OLrxMIPdfkTwSKjmXKSloS/b1Mb4i2QRViKaqgcJ0vqXBGLifeKM
dcuF+plqUVDDTrJqj9zN3DeCSgl0+Kt9gpuer73Y+g/Edr5cJr4XfAk1w5nA+0aj
MR0r7fLJ3pHR/g4KTo5uE6xrjciyNTmonGDJHcqggw2W4q9izlOWWnZffIcbHtE2
a/NrNd2QUzwDRGIA4XpsP+w5qNDA1EMuGW2XXlU+VYixn13fuj/um3CMAxpo86zS
JATwP4EPE4BVdQiYkWRLVHhwU1zlF+emBNOvEAjCeCo50R3Ft/2N4v8aqYfwr6Z8
bxbMms6Lg/meIPsFtMswlKXuzqnh5fGeswpbwP+NKAja+o8+dkVgbXBbbno9ErDJ
spSrB1w+sDBaytTCI/BbgLzUBMCVj0r7okSdcCKt+H3MEjMu/7W+UM+Y0DyRusAb
legTyOFGY+qSPorriczdkHK/0mmRNOMs7G3oSdlpely5dG5MVZKdlsDwhtN925i5
uKDqK+On2U71KLtGRlbpNVNNl4xdhJa8sqECd7Jiyj3TitMuPqpBGBBzSC81vUwi
LF13MWkCrRUt9YCjYeM2pBI3+bfZr9tnzVN0JY1z4E5QkCiF4o4iZW19v4FbZj5k
kXfbRMVz2flLr1tezjZ+oTuJb+h0wVQQkAAKZL1QeMwT1kxLli/vLZHkZI/T98bL
X0s0DevEA0jrnocXs9sWljofe+eR/+HMnUOsFVul1K0rtdTmBMpv1B5aKX0QRztT
ad5NyfkoTVvglE9I1ZesLlseDY4i386w3/cnbFSMvgkxfRDPa4cwyCdRSz1gksug
U00GOfBgS7acdCIVeY/UVaAd4R9HkCWpIWQaWWMauc3ILFHYlt5TNYn6WNrDrDt9
yPNAH9P/gvQt5N65dSEuA6NKIweq4nbDMCKrBRHL7J5MisxL3IiK33CrhzHnt1vG
7uUJukqlbegrl/ES2OkpV9jM4shpAGerytHdlCsbHEKYxh4rraw7i4gKbJ1FGG9V
M7T29olNcjEFCkaaRdqryqeuqV0ydMonGaQT8whQxVdDWRgwgkMSj+6NmbioO7Zj
G9jQAaiCiCbt1FpgZEGQtMjDtwBR7c1IfQUA9kzigfs2Ol6MoF4S8lWtHYjmihES
3A6rVGvuuNf566IjY6Q6PLJUpDWjxsdX5XI83SM8HEYcdLipBbONY6YDjMWfGhQd
DG1kGwOd2mzDUZH0hGsxogBs28S76+gO7CasBIWMr/Gd8T79vx5KW91f/X2krKkl
APbPo95BvTbIwRviHrXW8r9FdN4lL/lDhlLJfAiISH0+lfyZoAknOM4p5LwpuCzN
vME6E9j+0htZgbWnqsfhgwhH0D5SqYWXNhu0la/1Hdj1P/tdb3zFcz8LfEm9EnDO
4/7IgGUL2JheQhBZ62tVk0z+4waMcmv5rCiAoJ0MGa5PA1QQe9Dyanlp6u5PvmLO
1eNI1LQEy9YzFllZgtotvSfxVlPM4qcWMWvgltAIBl9AY+9K1cN8QGaU3IIlWaRX
0/OG05YCvVKg2acwheGPKjmRcZNFg5P7+CCe6TnGpuU4xv21dWxAV6EhVaD6CAHj
uzgUheO01VdNzJRfwzC+iWnKgkP6dFRIrlJYOiEY5cbmYfAyABHVxTnj4UE3+qji
iE7lRA4+YoiNNMkxBNxUEy5pwiM+a38r944Tx/ofHyXYHJocNnCghikm/v74VuVv
r8QacK++UGgNQ8PCC9AAskWf5r3an3zCKPDB8ioyWesZGboHO/ZVsANeaTTZjydJ
2cYUS6S5JK9+/Dw1eXFNQevVrw6ti5rKCF3QKf63X/ypKPqSPCAzwTy9hRl+4DoN
hGfvjHlVic3uwc5hq8Jurq+Fxf281XImMaZuY/Eekuo1cBJukInmWGMdQBe7zN7g
yduib+fmquC3eI3WTecDyzKjLc0p4bGaq1FjGUjONUMSLFtec9kTAhHF3mnMUYZ/
TGxsBccC9QuKK47WuSk+jpqaFJFez3Bd339r6q08ydLL9AXtEPD5CZe4R+01nGyn
V+z/hMFD/YujrUVVBZeFlKVYoa+2dHKRg+H2HBOCX+GSl4R1Ji7ze6JRDp0shjHr
c1zovnu8JCviKtyOeWidIir/RZVBCEb3HnuJmiwvbVaIuDQ2go/e6IGffb9esSdC
QEKNc1oeKbD/Om1EDxdU4VCs5/BL99W3ewd6TauHiz1NfngezBbTCySpnVgW9sMz
yhx+PZvcG9Yr3/NHT2SPngU8icivKOilP8dAhS6zEUea3WKVMIRKXcUOWsupp/0y
hZX/e48lf8Kdak8Z6XhGYjWb3u67DF9McCZowQiSIZs+xUEroM4qTLRNFjWCwN5k
ToEHEc2CwNkH1VYaeYTQgUysKIVUBXPwbxuh6Ao26Rv/FuOFRPwqkLfZqSGc9CYo
JDSj+WNvaOLFRG31G9Uk1eP4XqKUWjdqrRAxctb3tNXeM+O/SnLG5MfFJOmjcoSE
McBoZABbnPyQ6qm3hNJiT/V4mRllPeK2KxKb1exrEpYWvVLZijOb7qovbudh4BiH
g8Q8Ni67leHZ/XYm6m2s0Z2FshSINZY8tR8iG78J7oD+hzaY/JxPnv74vb7Q/vcK
UsgiGrnGyhJvdlf4xO4LDSdqvHRPSngNDkC4LHGEqug3fx5GuJvGKUjhX76jYcx2
FbVtK8DyX5T9l22U+Wi5FV0SqmEAwJcNMQNWfs0DAfIxgIxVeHi0cTz37ea2i5AO
NgPRtvLrQy56IHAWcRsMrFW1bfyNPh6bwwPO3sQNzXzxmdhdDYidvHQzW/uu5W5k
7vaem94ArI/n/eAk0wEcSs9PthdkMEUiaYzLRKRqAxvFJM4FdojqnqyOZ9raDhs4
Ly+1SIfHqTzapew2hL2XsJhxLg4roAbzNrQ01ewWCHF6FgH+/vcjZlwotqd3JWCE
NyBlZLLvscGh+8rvkfRf7HyPi53fmY19AhOK5BroO/kfEx8kDjtzHQo/zQDxvSrp
09a1iWYyEprt0IiPeRIssU1gENsBWj4GoWQv1qnXp10fVWJlLrjbyT8RbBhqptJ7
I2QXobCVzg5rbfSYWBUtVxySrBm7VU91Ug80DgbSPwQRzNyPJH473qYc7jeay+l7
7Lxv00MBtVDmbh6PYbLBcNmaCHFMGapYtMvXbM5fQoEJePsy/4Y8pMOVhwDFlD4o
SCuFgQuVGN4sDGmBuCrLQ/Z1q1AkjdXBzY1Gu+4M/SvjtxiAHtf0ifdyfuce47T6
21vkTOyjtkvn3MPS2P8U3ZfATKTSFphTkr+ZS274GjQHRU53WLNiaRNMZgfqucwz
V3ulNT5uKRisT+/7IRU9Q0B05BIsAhcWLVvkV0q6cpNknfngQxi7kGb1rH8W6Dk0
aahHT8lkgO845NujGT/++q0KWKUBJSyzGuGZYuLWAMTHnu8cBosc2O43EjVjjyDp
8x/RePQ0o7F5CMGTS2t1ooAfBfxD1UBIDsFM1PV/x0S4W6c6CwAaBsCr7/zM6+yx
+BNfPDnrHXmV0TUs+daxGWXWxln/sWuyJjH8sODqah4Fo3Js2CnXDXQ5yqxzBwOX
SSYLOStL/jMRoKDONUZi5uRu9B1KpDM5rin+i4tiq9wpPy7MG47ipML2XXzXi7Pi
vbJaM4UIIqzxWvSgjXme/tuzZEv/ULsasckqBGiVA+C074la3yztRT9veUHnLVxk
/67lNpNGDXILC4M1ktFxDE+m4xZrlV9/94Eg4xqsvYQMAbMInMjtoJe8TLMIy6hH
q+x6s5JXENySxbx7TSyR5JLzFpKyyDsOTc62O+QVUV+IR4ntbnRuWQqK8Yo+j0KO
nG8OjBQrn0UZabZVu4yB6r2REQtWF6pIgXtC9lVcvvtm/XtNDO+xHFcUaIlmgUSZ
NwD02/C9rX2HCDOTzMTewRbuVsfOA5ed3ouDUSWeZga6aeyKyOOjCr+cMTVTr7AE
rKUDNKMZG0IbGPawTihFOqk68IcHDyj8qdJVrnFZDwzGrRI3boLafWPKr15Vtf90
iPnCh5KjRhSYPT83MlN8FZ3h9Uy0z8WtRsG0jHztgw41dd/mITYfRVDNUrgr4KKO
5X24yusHZMvQvGlE5LzAmMM48a4YtLfc2kUUaajPyHiy3Q4ZQvNAAOUb3sbqaBAU
gZ+FAghDOXzshs4y5eyeFse5qkG/upLvxqqt6rgeTrFG092numRasjaK+JwvRPZr
Xdf0rBqFXQ0lTai41CPppl4hOi4fmg5B+MNvjPXnXAzIF8965w1EFX8wsy5m5qal
X0IO/DohhwzgN/N9lTc7KDAu0cXka812rJcJifg1Rb/zRGC0JnJFjQCaN1mAwZUm
x9ioQt76qxdahbD6tp/P5zCPn0Eh43cEefIaNgwGbN2Tu2JJcSunkAiAopLSG8Fe
ST+grWGKPTCMTaDK/3bKpn9idzddMiDtoBliyh33J38yhwI2UqmEBeYjGw5ttvaT
rp76Ek5citR3XBiKrybk2XpWzvLrunjFnCxtldiMlnLnAMkyzCkM5UPlV69IryOh
ZhgU3FERyr5aNrqQ+HTJvrWhe/rsIArEQZyRIxffmognJu7IC3edBmzu2A4yKSAJ
h3+9PQMrJrULyDNGpUj0L0rLkdD0iFkg/0vnT/sQfEWX+b0IctARZDP8d1awdMOs
/y7BAJLmJIIQqSkK+LoEQNsTtX/4w1TjCite5miPH61LAO52PgiCVRo54Hz/IEj7
gwmQGEq2cSs9TTuD5cT6kDYKXQGQFebkFZK2XMeDGXhKPMqvGepYenfC3Oe8cAih
fqzn5scJVrnW2fESlfJ+8x+bmFUVZe0TLS9bwIAXCfnzj38RLSE6GJtqXZk1LvW/
NfE2HOFm0LTJyZ4lvsibx6ZmQip7LiwRLh5eEPbAxM3SelsfQCWLWv/rxWUGirvj
3SJ74oK0JPVLIJbHohQJWkZ8W8bOjwRQk08VPd1mS0Y1djE5NjjeLixD+3eW3H0l
OFMYsvSnL5wbAudx/Q4wpTGmlRw5fUiONpgLmOBTNYX5/Pb7DYzEbcyzYicE7e6W
L2BLB+NqwpZ4QWlZvJVzBxySMOOO06x5s+To7F+a2Q3emfmMIjRT93kY5GnrMOHO
T9hqd31WUSubxmkgRME6C4PWtWhjYN4+sE3ZKQC8SerCwJI3rYiBymjDTp2sUmrM
TYNOQKdRrhNfwHKRaQNwq2KT/E0sdSyEtbgAx/TAKID0I3Nk5xFVEYuf6OP77npp
O2ErB2AOAqkkZhshmKxFr5GzOsPZc+WHEmXH1k68BJvbtIPMEsfd7j7ND/JTV92I
SgP8UcKBcaiTMmIMXiS0DW6M3udRsQcSaBoxAKyV7OjCdEvzVK9o2o2TsVKsVCba
zVDj1gK3FkpgTxOHrPayeRUpItYM9Iv+6SI+v0ZASRzaqfun8dHSftSQY4xjk4vu
iFQQxr+ZzZykwZNGA5yqDB5axfy6kINDdhSRfN8gHCg5cqh9w6x1DyRHOa1AvSR4
qqIe3B0n9IZS1rNUQ7xvYDJGc5kJty64lif84KLviPT4EMfb02UnhSmGtllQiccy
OYJd+Lic3F1poKDNpuv2i0azRL+LuNFsatcoieP4l6Nve5DrrbGbwVCErrzI4QZP
+XXBOdrhBEKORgldNkQJLsInXjX6IMw8XA1A8TOfqak4x9j45okgp3qgpHuhhOZQ
3CKapjSLtmDXDrBYJ3Suaitac24TWdXos5p6l/U8iMdL0UXH262KaQvly2y68bDF
QF133xaAsSZdriWhH5W8TkljcHIS9vZhOUO0oZjeLC79HF95OUEGU3cbKUCVtiqX
i+m9HL5tl3oDbtqPRz3vt8/cbI6wCNIJDJz7Abik5zbuDGDD8PjecWbH/N+ObYvb
3NQzBBvw4vH4peQwS/ziO2RqzuKDlxrg1l5zGsQrzOQfq+h+EpiGC4+X75bxIe91
+Np9qIJx9IUegALy9UHONoKuqEpYl2CtwElqi5zPS1NB1q2gGmBAxDpsQOlAt7UY
X2ljD04gh8YFVa/G1PT+ALVyvIVslzusSnesjGltHL7HftdnF9oUZDdEPS5HoLyY
gsL0ElsoA/mavX2uiuU06QgKAKrcoSaM1Xb+T7vwuZgGEjeJOmtV1KuD5++uhUon
shoQbZXK+24EYwNIZl7CkCRjECL3medMl2cV+QZuFDZJvmZBScOXJgKY76db4mTG
H11FNzsENEgz4KHCBKlOjDfF1Qd2ohz4jRPAvgfk5N4DWY8JuqLgVNDFOISa7whN
yhNwvGuy9UMVjBvHmXLkqd4ylwJ2F4vlliTV/urWBkrDWZxR+8j+l9vR7jKx2muN
4jpBU1bsmlzCXe4A28pcf5UifoITufvTvZn0g0JqiXHhB7xVAnTG0JJ5um226u54
yCFCPkdT+ecg7/a3rRHW3ESpMIF9MG1xSuJujm/ndKWmcOEAPuDzv3u7bxYabR++
lWUjUGCgLb3kxO5g3CCkAmSeAVr9RIx5z/9rVqrEasZERt6UKFiq+2Ftpl/RYpZw
Fb2TIVnaQzGYTexIj0VWrNTOMo5eWjOQMkgWJg/fTHmzv5TtTM/j9rZMWvMAHJGf
QIEExvLc/WIOWxTT9IVyECuB5yWu3wwG0y2xK8ilneqQZ9EXlYrLOn4Fi1B/02rC
tDoTFSSvkXgO2Vbft/hFzxTWs0MLrspp7/bovv0K1fWvWSlAxjqU8KRP0rt+zsS4
pG8dxmnqajC6dvvgUmpOIn/nae1XY2nLkc8DKCmYf+VrQ3ABD66MUoFt0Kk+FLAA
N5qjNKHcO7/RHRONDOtLPEYBTh8BJJ4PK5gUu9sul7Wky826HyiLktgNfXp1EPCC
gOmmRwRfxaIfkAAtzr0pf2hSM6BGYohLBFqS9W0X6lnRE5HxZZIto2ob0h+1Zz4y
htSe/nHCT4ImNlyPiJTaR10oc7tMKDiX7dbkjyCdzctE1jEqecU6FK97UzKqimoO
bLO/oM1T5XSf930guETfCey41icKoYeIcTMzNlNfiUfbUUd0Ui07ItfnKkf3PSE1
iiixky9nYTBk0tJk5m9j56KfzuIembSqguzug6U73gso8QcnFuZtK4fB62xxnjAt
Yj7aarh5P8+s+aHP3wAjNwN0ww7DdatGN/sVYXDJ8wPK88TjyUvL5f2PCMXXQVIK
gzaSq/ubZH22jcSJRasPsFRTSGcmXtwQnK7yEU+aVNvASZURGg04zh/AvHVFeSzV
/qwJPjn2QmoyebEQ4YVuMmiRyDop7WlWvQtW6n7uU851MTAvRLuuwENfjAcxrMh0
8Uso2wj1p1b0Xer+UTNEuShMPlVE5IH6RuSZeQETXkeho8L9GcfGgZiKd37/GJTL
d/8A4/KXdYDMr0zCFn0jDmIXg4/dZ29xyRPTXRH3qzSd5pFPYOnfx7qo0BHBCdqT
wXSpgjtNQ48lT4Y8fcP6QybkclYG+pO6ce3VRDJjKj2bAK3al4dsSh8o9qX6GMBP
qtsjXGYpUWme9XKnh9RecWVVZ+/3wnSZkOfN5PG0hkc5ABOyNE4UoGMNI/CStfZ+
WCmuB/8T6dbu9+2UoHOheyUaXGhjUx3h++G69SgbvXlwIufJsK5+Mt41jaE0IGcc
g0Qqt0VENJJgLFkQ1yji+33yT9u3WvwrcJ9oOfR8jYidrIH145B0JtvnsrQSZEIb
+oflC5Jjpxwhf7nsS5khtXlVNhoy1U63O7HSa8iQaBf1ciVuG86wOtfHxtfPbcis
oYAUvop7871ncIRa7aQuM7ys1dNU8T5+rTLnrNxiN1fgouC9e4TmXVoFgoAbE6yW
MuXZAxAJBOHNHN2r94iPki60XyEX+m2Wb3gBApqA26y8iVIel8DqROuPlnVkulQr
Es5reSt2aqXWnuhjGGFUFtxbQ9sAPK++SUvyDBPJl40LN5BAY9NB4PRXztM02R1v
k0ZM63VctqvgdCQqWx6ZGOy8UPcTfz2dGk+Ucz/exEBfvzipLRA9XkSjvCyFxdOQ
aUqyoygXek9FE1Qmy0lvrDaPy/D1MTZYUZQeWOMAhqkNq5JUG0+SXbPDQuqIscQE
ARwnMKjwjSmv0+ed0QbvK75bYZmRD8GqnEPMuPyPD8i7AQfnwtZ6WMDIHYhSzauu
LPGB5OtUFH5+KhCb2ousFi0E7Rrfh/2cmg2QraHNeQWaumfW48RAJGz3RKw/GyEg
dRvru04x/FbirjOe8anOSM3FgJDichsyiJoJbKZKK0LeTPE8GjOJOpklH7vZMcwu
09O6+vG78l2UZkoVP4EAZT9jlF4R35vn1RSf2HLQKvW6c6bx1+2G0xHt6/+78ohy
nSo3kJYasJvvIsi/RlJ2B0HVr1BzrI+5b2yTqTjBaniFjAMQiJMBshjC5zNJHx5G
0GfIofjKM3iGx249P9L6+FhIcrs4FzkjopvB1mHekAueNURLkwgS4TNteOM8TlWJ
Y3KhgL6vLZoYugjYMRPhC5zeoCqTMn0H8GIX5ckqcKRARYzYCumSZdpICtUJzRDp
+XNMtnN5QEzoHy9Zht46TQT1+bra8s992s0/c8dwwJKdByu6obNeefCtV4IoPcFd
kgqOIkLldO3BLlbT+dvwrERJVhqEC6rfM8ZsSllltOH+OLh0IgKBBONgdu9KdZrr
9lNrr+XnXhuMdcvRbzmpfhK9ynTxF1UBv1dz2Uqcp7ZfAGz0pkt9RATQOLZRTmGg
wqLZvk8Y7pt91IqEXXL+pKSdQN+iLeOmXo+zPG7yprD9q+siz8i80c0OxmoM4DeU
JJdLimP6Cu1KUIpD/cqLHV5AdNhgWqGRFhPooSDuy9y2GjiNsI0yDGf6AScPeR8q
35NBXW8JK4u2Pm/GKa+0+dhtSB89CKxcpkH1jIHRP+L+emuCS0n8xBbNjAb+wpaV
1yREjH3Y3WG2aspb7Wug7EmRwzBXxTeusHPYSrPXE1lyhuadi/FqFHQ8yi4MIgO5
2+BPSrirZqfDORGxftQqctC55GYjpfdMBNTX8jgYugMMGNChH9TbXeAIW9BGi4EO
Gf9bV43q0kpJ/qehBc5fF9WJ5eYO2G0a9El5LncbsBeQJ2jaGsfmB5HfCWaj3qng
E5nGQ7h5xp/HhcNDe2WUfOnXU4/xROJEFUv9Wk1fQ3GLWOA26ixFtwjastgheWT+
dlly+cpqPyR3hcp0nURUJWmRQFqVsGoW5l9Cf8GrBeEgYqK8YT8C5EhAc9A/4U/v
oOlbPI4pUSCpL8XmSbiPxktwfD/yAdOazv2fthclOcJUIN0zzrmmMQoB7f6j0EHA
i244w/NWM+N/v++4QNppL1JeleRi7oTMwhjEWhIrC2RU4nHRw0VqOuXFSlewgkm4
Hwi+IIHDOs9FupK6pUfur4Nd061a3UsrumG9EHTxAut/88dPP3zyx3sV6Ad6t+bl
oa+TnESNvkj9i3Fd5DsgMXwWgHrm2yJN0CWl0GqdX0ELXEjwpk65ARaHSZpUPrwL
VIg5n+MgPKzrfoyBeEIveUUvcFywUtFNA1IfnQN56Bhyg2mD5wPSR64r2rSovsj4
oI/oDQ6+MM7a8QtLgpYtaWp9aa8pDgRIHSgQsOlEBdmEOT3tSMqL/LSL3Wv2j09u
yeBlFhnpk+n9NOLNdaKd8e7cOBRU6i5c35mMoKjhGDLZwXBhFb0ddDqCzq9mpPvn
PcrUVlBrU1Sbs2rsSQTHTX4RDOnuXfAPK/GBi3bBcOvymgBnpyE2OPw9IfMe5isI
co6ocwNWqLi/XVj5BhdfSipA53r34pxHBDk0TnapuajtFmAtulLblpLTjyRlo7p4
RiUGc2AQUWia/gs6ok0xCXwcmxmyDwebTcASUq9X3w30esuk9EtUAlQNFv7+6NBH
gpjLhZIZMbmNnesw45IpihjkF/Z8y9iA7jOXCrX69ISJ0gYPl1qs4oN2TuWkdkmt
FbTZfcoIRe8icm8qCdbhr431lMtEB+zVYQluw9C718PDnTvSa7KvyEIisZWGn7n4
Ok/davcVkcR5xPe5rkZYD+0TUoHaqibaAFFwOp98OAe996o1scy27jmjX8Ta7t1Y
qbPaxERbbyvx+p/bhlRyUd8k0CwdyUKVbbVU6sXX0WnVmdxTGfXYE2hgeCgVY4PR
KpSuOo5QZ9MOreCFKYRmuzGY0ah9gSbcnIIXzaVVryj0tcAOGj8iiyhaM+sO4Vfo
aeZ2oJlbJZO7ftzCfHzz3GSO+8Hwgm8TgFcuHQi4JZ/7qTICIBOMZQ/1Oo4YZDnL
cen3a4+Bs/qMGQXgERrTAVDfyaYN1tMbbWXeXnheX+qE0P0Cw547vS09Yyqt1hka
snxLtxXmSmdgAohAb3MUsTIJZtAiSK6/voBIuuMxUIPraOuABgR/khNgQBxnro7r
VoDwjG8ig9fLd9goWM/UQTke2S84V0UKoVYnpfS+vIu7i7YOTFMcJ+oc0CCAMR4p
p65qEBYzH+3MCl5S4dCOh4Da1k7YKIwB7n0kp6qtFvxkkH4FOwBMRf35dUavxtAB
XCT7tUMA22h2Zq6h/b1BvykWJ0xtIHjPOiDTTDg5tniMGhvkTCM7qSHgt7QY3Ftp
DWv74Wzt/Scs9El8Q206rXVUXcABq4N7Ltsi+2BPzALg/mpDm1yEnNGly1fvgqIV
7oyifTpYaTW6oIAC9tu56VQlq9JBXwj6TNvq5zZcoKUymvNnKoR/+8UwhSN1WnAO
d01BqF7EUSOAM4A6/j4RrEQdEkNet+NhVr4C1Wopj1lsFq8L/CAKfQSEHnIqDQoC
5XetbUOqlVfMHnfZRp67dqO5JNN2EBjaIV+BsuXkJ0DdCFtZTAA9ahQDLdrCgh7f
tNMQhbtRCNNUphiOcbHPT2kxvwhJrShp5nI5saxuEHaFf3p3GfRJcIRnUBiKrHYG
xvb+KRk6KFaDlF5QSX8+0ubqTa0txyceYwKV+z3JzpC7C8al7O7z8Czh/1DrbZHJ
efw1gOHo5EwAEs4X5CnBpjKwVDzJWgVkA2TQDFKbU1A/wboZgmNAs2xht7BiGDjY
xXB2Cb6lI9VbPRs/9/AegVJog4VSo/i5FZO7QROnGSYQoZZ2od2eTxFa0DAxDrAM
mS8eV+Nsao0RouyFDDxOeaXGkB33BU3AiJl0ORHTBhiyqixPuj6uSjhw3juHPRET
u76bv7q981ZwQz65pP++kGKjEk+L3B1SQGXrRUT1J+FCaenGzhy5vZSEwGNWEmqG
nOTppZdK04U6GAeqezLKgC3+z8CyhvrvtfPJgD6dNDItNEv463iLuCQ/exh28joD
BbmhkCuqvMJm2Ei8i30QJKq3EphDMraKJxHMxn2D2wugfDqn4forGSWo+rcieCo4
NA4mn+5/1dkdStLdnAQpf0YvhZNa3Pl8An5oEsSw3rK079/xaMCducDyQ3UKVj5C
swd5LmuPKihYMydifipwCaB83BDt00i9nLt1MKCqVq+uNOGBL8rG8jnIRkuKVZSn
CGQdf9tIR08dFq5G0slEUWY9fnG8rnupf6hXjLjQaTi49H2/O+3LRtauNXws9hEP
IEBJPp0NFw64zcvQS5Ds4a96oBtB7PlUn/q6jAyi2RP2PM5sLrrN7LRpBMBSbvTB
B9Bq6XIn5+blzo2AjKTnQsjZ2jw5elfWr3xfLe2NdrjDSx1nYQUsrUgkZuM37WBH
+3oPNb7KtLogf1O6G9NySM4UVtHnZbtNA+HSBidJHrmZPt9PFIWwkL39d33n3o7u
xYlFC6AQjYPRrhRzSQt6S4Y5vISorJY1wg35oKmSn+D/n5pPozPb2/qlH5MMWjgz
Pw1asnMla5erMzxEVIwymO5ZkmwqMe6VqsbRht9J3Og7QPLIJ78dmi0FjcSkPKid
qnGZiVzdkHJDhDKkzRTIJmqadTCf9fNlujz6ZPYAPmdDICkFlT3pY6IIziVi4p/j
FZmtSC2mOLzYlneykJq5Aq1Nt3rXZSgwZXC+hyPgbLFhqIC59Akwe5VDfwLiW4KD
HJ5pYY9LgaJlFlzIjfSzJTa3x189mdW8EusFDx0KFE9irqWff84l+y29OWClD4pz
FSbSQqclri5PFRsfMZ9SbdKc5EOe2SrjP8ZrxZtvRl7RgzyWVrWlhXl0wDTSieqH
QhJ9vsqw9C15kdFq0NMkwJ4BGLXK6ISK8Xo89DKnuZ9KlF7YKFBJDE+daK/AcSIM
NfSbPN6DzA2pN3HacpW7o9ZGKLIm09c0yPiJ+enVQipDIMs/4Zeg0IgwpIQBLf/W
6CKLJcsOUVfQIAO1HCVNXvqpMgqTU62yobYIufboENNqVbtocGxgghSwJU75dWYA
Cl2QGBcXcGVS2J+rlv6O1LCwvAa1lelHrZLI2LmJAbeZSY8sKSUAyVy9YIWtxhRZ
qC6Zg2PS8dEteKvr/+DA6eT4KoJLCE6esXebntQ0z+EFZLT2OodoxP9u7R6fVcP9
C8it0Bm+/6RWJb+e1hm+GLbBHnegeb2BJXWp4+MKgrlBqfXw6s175vg1QUXojoov
ykPqFh19J5VqCFTuNOrPfGeJcsXKL/w6dnv88S7asQU64BxeB95SsvIlMzkjvNgq
1BrAqaUrFHoB2JV3L/EM3dVpnIyfO/S2bIBNtWKT5+VHFaxPsLViHgCxoVRQqU35
awy8b7P23Ze/gNeZf+e23H/GMHGplY75uo88Hfdg8e4USxuLtaTxncfE+aUoxDon
OaPmjH3dML9JQ2VNCd7TKZe3WUMn4rRl3T9jkiouLLQNW1rNmDor9o3i6kqW8BuJ
XnZa9c8VUIqrKWnRd11CDIXrBoytQDC0eg0E+XoyxEt2kbGtUxnziQcVNXuIs9tg
ftym2cAozzcV3rap7si4fHNb6MqtJU0Y0actpKgp9k/XzwofTSaTs8ORhFCObURE
NJ/GBVZXX3MTaDoykOSSXL6fYhK2TYPJzijCdy/FVEmIJbGilVW+3pMKx77kYbat
LC2ZpgZl0n4rTTzqy2F3MbOCYjJ4i4rnDv2JulWNM+NA0NM2DiXbmguDBcLMYHpd
Uje7DfolDa+UA3NMJkpk0Emo3F+++q4y5P0SV6vCQ93OG+W5Th9ANpERZzya/dCn
8W7mHysWwXx4vUKx1RQBac+iMBx1yW8Qq1r38v6PLYlceEgdNKqnCd0K3OBv1Oqn
/8uGY+Mp5O171ycfdeKtFyGgAuoTTQf7UoRasB/cyQGGxVvrAtyE6BszbkgGNfuc
3UX+zFO6l16nXbjnl+fXHNeaa8r1/gk6WAe7CLjdN1AudXgW0VHtvsS/CrrA8Tkx
c2xdZnZPcQGQOKnJuLE8GGZRmu9/v9Xpqnz8TZWiftFrntFlDBeWE66zVaogD08k
GQ8EOu649F+ZxMqnD6lEIk130strbH55AmQlwab3tfyC3Y8kNN215mzxEk/lrEdT
2P+J796fc5NH8J7lm9WXymr4D9IOL8d7bRL8+K8WCmD/rff6jARm9soMLx40f1x2
dGXONC6dSZxejBl9tIkVUEK3uKODpsITNBZDupbMbbi37HDYR7rJYzsfhnj/6RX5
XYCBL/D3k3T5Mn2rQim+eNNpXHwyMUWMPHI/DlwWDyYVM8AU8xX9Q9q0sZRqy26K
0552767XQv9K9HgqdDE5agSBvyAAxwb3m8Le79LCALYAXGYUxSALGzRcb9p9jJzy
CIwznP6X6guioclToQzaFOGVeslplDoFNf/8e0EpbPDlJ8N1btZZSivcD8eLuPaL
9yIlQHDhmELlt7xhI7MT5HTmOGX+sGTlcfRuEwffmMAZP3LJk/0MKQHq278v280i
gFvBpLZ0gTzoywtQFDa38NJc2gpE/vaT0AzKKYeLY7PAcyb/mnys9uETwBlKzPhf
e7Tg1kpYSFencDWF4KGg/SZOF+I4/olwHJfi558wFn/zp64D8/CHKgHXIilVbbJ3
MD0wGkBoUTRwf5vTFkVQEN85ZYhKjHqJHtkqc40bYSA3dD4OPYApERqmJ003BZyp
qnWwV6KekBMNKR2HEawpMg81Ojm8Zi5LdlfETWpkXfelaPY+XRYpLq2phxk0Xap8
+uaTxS9YqHAIR4uyWmSAErGl+h5qvBWA5e2YrTbH+udO2ChbeTBPLKv0aK+A84Jq
TFWxUumxS31VnZE2W2euQB89aPiQvo8wjGRCp2L3fPOqPGMPz7fx8j6sI16J16MY
XKtVKfhQ5pGkezRTEmJOHetNL7vfO5XmnkP4OK2baBP9BZy7It1YtbgUTmj7/LBY
N46R/WnWPOOwpXPi9/vlxGIUmzS7RdrqU4QUR0uKmtAZQ/wOm2jH9XNgReo0G1G9
F8ZYJi3VOoSqJn41SE/5N2/5dKAIVQSIuy7rmanctgk0CwrruGc40oVfUequ8muj
2V3vLfWvj4J7PBcRmF89VExOc5EcRmpVjvd3Adh//3dwRBaoLy+muGGLj7I9KrVe
pmtJBTfQvykieBg8fS6cvdmeHRBO+MQGbNSvkwiuNb41qi+EPrx71f834ebLc4Le
1Tn9i4wzooA/feKmkb1zZofdf6kwUDkYR25UxZi9GTHQ0byM5GQJt0Fj4JFPzKyl
Xzo/XzwNlhpbXGWDe5kQHexPCvw3jmA313NeGt4Yws1ynN5UTQRh08m43FrTnH4x
FWIWCSr2XJGcwhrkqU06zPTySrff8j9JenGl5LgqYqSgibzV36iTtxjiztu6kDat
qOpP45ncqsRgSYymMtkIUuQDMi/Dn+ZWMHWZS+wse87AzobY2AJN3xs8IyK5fuFV
kU0z4HKwQKR8KLgRYXzycQ+NymOScSraz7nf9wknQhIbB6Y24a0agf12KDgnHT4d
j8gac8WFfROYcOZQD688v/1SLOm6yxJp3qb1QA3dE4cSYzCnW4j6i60UQR4kzeIM
F3YXpvvKrhuAGMD/upDqQogf/lUGPpwghqP9YfMs5ZBAfzcSWWRNLJp14kdlSbUp
76JHPELNOcgEzw3b+k8h/KIImu1r2FZbY/dfInUWSLWQjCag0Zp+D6SiPdBBk1KW
EITeynpVlo/Q+TBK6iTqDEyG223CLK0FTkcmcv+T9/bHgs5sC8MHCUDAjVOg3QZN
kqazKtooOv6854isZZDuIdpH1B5VKsLb4I/8d2cJcZl9q6KVXsyExAsU59Mbb5oO
ExTxOUsBcuwPJtjOKORUg5k2eUStGVhRb9Rn0brzOG+kCnTI9mdRUKg/YMx+/5N2
30GA4RcpvkVkwaCuRFQe4171cX0ux1niXAaiteEg6mV4r6pT/jKUTewb/6ml6DXd
fj5wgLt2mDbwukWvMZbin6RlqjWKR0jLdO4wn9kjC4ydttFtAHBjnPsOztZcufjt
UmoIgzNTuw+ITT9jGxOxku3PDBVX+h+YWdyKnuxs4jF4oRLcJickGs3Co8PZSSjl
w2lRHLuVoy2b0YnWm7MJ/M2SlVgFT6QltNDNmqYMG/Ahrt5eR4E1mQxvdBdG0uk+
LgR0gOHPz9fX2hn2tKrX3nnWEhAm9gn7eAbqFUfTjkgFN6yHhpRDl+H5EuT/eRHB
cqe6hVClkg/3a7EsKdywAF6T2jWS2fYiR8CheDkM7m3cuqhmWV8d4ZrzdocRt/2Y
0BFkEDrX6FAXsL7IWXZJmtjptXj5yip+ntt3kSgZgwT0zWNggAdyTkLkCcVu9pPt
qaa4CNm1TSL01Es5nKWDY6fWQj7kX9ReovuuvrWN6sWWx+AtTPruDBOSkTfK7Zt6
V8LD2MkNMH9xeSBY8CTSFOHsMRLKFUhyhHUdT8Ne5fbINNyTGwZ9Y6MWhU6rqm16
FbrVB4ASKuYHnjUWmRzgC8whgW6vHp9/NwxEdwIXMzfs1Lk6gJe4j7ozOalDrL66
Xnu4N5W9sePk2vp8PSQLv+So7ts1SG2M4z4lYJZ25ls1PCo5M5N+BMK4VJr+70Hi
ysOsztvwGqqcI3Ghw+pqzVlGm0kJKrNT02BqPgsOhkhsQo2kRoLsnYw/saYVY5Nx
DuaIkDqnbQLCV736qG9tH4Xen++2GiAyrR+dPPaQuFqP8EaN/lKZu9FRa82KdpRF
Xmi16h+qUTz6GXpNxe5/QGcwuKSJHUUWpBVigbpPy/3cYgBNzDr8em+sUpI24m4G
kxBvOJG1c2GrhMyUT+uzaXxOoOv9iAyy9dcu8qc3fPPvR6XLZcsnz5MvN8wZupGJ
VSdpgfXcHNihgzMZt9b8/zOJjhBX0D0n/X/bpfMVEml0UrACUk5uOfrjem+89Dz4
bAIPiYmrLE7FXuSwhO2h+HQOC0RoQt72eL1f/g8VtTRvxgm2KxQfarU+Zcin9Ais
8+cJVWxsh2AyxkKyNBjKN83zhCtfTaWm2xPyGlirMtH+w7Gezp6P1un/glScK5xF
o0HeAcJKM8+T1uL3gMlxbiLtrYr+aoz9u84JSv0eqSGwtl7W2RYh5KXnthScO+up
q1hseCI1bgF9w9MM3WOf9spQ36BUqZGdv5huy7rqNexyRqBmaBZGI2pTm3tZhlWo
I8W8GxPFW2TWQusheSpI4NS3mBQoisNAPME6EQD+6uAbfBoxcvy8EsLDYvuWqCfz
cqm2bxpQdIP18qmB3fLWCNXMZcKkmFCyPZP9Jb0CkyvaAnKqTM5nNrbC2YfHAc8R
67uyfeHmcFpJhgG0WX/jHvAs2eawqCBsxyb3DdLMtSqNEQY2a0vlBj+H8aCvcXiO
2+CJYnDWLFjwQhqvM/TpVLKUOj31l0MgZIsnALufm6g+nhTgmsfj9DJdTNsEAyDD
xchO/DqzkWmLvFGJZnwM0je3cy+8V2w6dIOop3fr9ry1SyKPIcDZzwrq3T7CRWaI
K3LZBjZ20pGjfkLY9i0IOmUKVPrXFu6QSq0zEtdYyHd9No5ED7KZN3WpGbym2Y3G
xcZWgEl1+MjSyUZbBis7mL4ZhjaUg+pwpdWMfmP4Ya1q1DH+rPAu4AR6/eneJgiQ
m1HY1QxuNObL60h/rgLMV4tyHenjkRg/W82cFWPzbOSwyY/7H4w/CysswqwZkR1K
63mmK96j6Ohmql14R82OLWRyeKQpTTbk6oiVy5NsELMbyoLhT6nrCWhLkOFURFl2
WlOmy8LxoaZbRgp4ItgBUjRPc0OOpqV6fJYxTIMQVH1OKgM1X6EFWMqgvXi074ez
EWOzCd70C96FbTSlfA7sxLsbMBLaXTGJEdEbuSDiT3fQajioWjN6Wcvqcyax9IhD
zu6V8RG1JqfaLbGwCzNSODIqavtN7fqLa/CFBzHicAt9hU8mgJriu4E56hnT+qsC
vUujtY0gd8vsxl4HW+OXKo5p0F05EVj/ibWgfq9SlWPxsvUyeEF9iDnGzgp48acf
q7AvHr9JwhjiXekMUZr+NTperkYNU0bUC7fwQNGytCyNuk4rLBnikR31Q4UY+I1+
kubifTw5D4n4L9O5iAAPUZLGL8Y0gVA0fTDiA/dK2vLLeqwtBOhENehEV2LVX+3j
KU7zDljY6qTgl1Zg8Op81VpqeS0Q0gailX6G7rjSC6cGTo2lyHIDQb474j+bTvix
dQk09dbKyQBJiLb/rKNNlV1eB0W3F13ckgGQJQCfIpw=
`protect end_protected