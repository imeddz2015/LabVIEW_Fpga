`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 1824 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/9huKRhRMtvnNqb3Z+UU7TahEoHV+T8U3P3ufru7l1O
3DlgtZzb9QxCbOjthp9+wDkjygH0eUfDrEl1ovhZG62HvmJg4YFiQxxW/Yim5dCf
8f8okLngF97E+3fIE3+1wFgyHlD890dgbWUZS/F5gSfnaETetpU9Z49y99TTNInq
NqpeZulD12mO+L9w7XCTGWxSe3T51UQPNGWYjn+VvMh+98V/bbgcv4YaVsZTINEb
X9u+dMXmSIrMf+jE0M/8IOJ1VITp3sqhQm5cHEHrlgWb9BwcfXLMrYuW2uACWyIt
Ft2LsfjuTsgLsdQoJ6/TexqniKxBLeV39d5kvAzR1pTDOG8guklCPTUqix8vpPW3
Bby/iWgN/B8b2vBRifeXzSAWgLZH/qmRHJbwMTE+wsZ38h01VVwoBBFkEDy+ZMGy
ECo3PhwMgOTIJsjHsjikfTETxnmlYupGC4u6dhdtuZEm6kAFtS5FvqDAuwezaOf7
zmrx1t6k0uo9VpTvBTIiMJMucjJhG3Z4GMZ+FMKGUXkoB8BpLckIfKolubzOSTRd
R8HFkaLC96s+oJWlYUUa/YJKVuDnmFE/yeSCwthqmeEPdIkDIN/grW2QrgC0qEym
4KOciFjxZdth2AwrOinxQnY9GawDyCgH+4PHuD4eM5FjTwf29NEwaLhVaFRt97f+
CY/5Gd0g4GUg8rcfpUidj5cWNmd6LpQrFnLzPk6Rwzm5VQqlVEIhvUsfs/t0vA3B
6VvSR0edyXUyb4oClXdYddx4qFGigXpQa+SUm6n62nXSAwwyKYkcXP4YiJkd/QGX
OdZxt9zbHf/BLNw4wJa9Ozt/uqIv2H/TFL6YQTunmA+Nfc2FmW/56Flqxi+cIIW0
svuQH5IAEmeQS5l4OiZbMr8X2ZMeSllikeHj/0EFDzR0SKvwDF2ezadp2xaFPYlV
5EWiJiu6JDat6sRIswRsJW1zIPrH3NGQeaAmr0eSnBsVy3ehR3zexTEIhuDT9cAm
QybzboyVsGgNvi0pNht/uv7OVph28nV0UbnyeqKevkal1U3tuUO9fzxbzJlMuGrG
Ya2pBXBqM/q9hiYn/GP3/ZnmPBigPvE0DmuzYVmhMz2uKk2JLe/HroNmboV8ECx9
Vgg6fK/8saPEmNrG7hPAUMqC8swOkT+OP+NHAcX8uunUdXsUNdggElTnE5rJZUAW
rPIkrCkYubK4JJSVbQRmfyCBs4vAtJ71V55welZnR5LMa9aT3P9CIxNNxyQwZLT1
bM+HKLqZ9zCYS7ABIREoW3SVK9JD37D0CXwFuBWcEhWk6y5zCLkKm1rk8o/yFbOo
rgJmlB+VD1nKWFT7RykgreIOeGFSG4t01uXzc3LlF/lEqpVasgNSbEjCzHQdcB1O
vVvZSAPpNbDYFZd26jnkthOHX1cXrN44DAVs9KXr8JuCzJTWAomWOc5dFsS5bsgv
7yyCKUEgi2GJAStkOqAGMQTTByXhtX9irsP2MLb8OJB6quNEcO3l+eyYgaK+3ibl
sgymjiXdKX6frbEo7fWV0PpmRxnOCgk9/NeFLI5t6skNJuao6TQ1QU2v3M2//HrT
z2lVrrpQPg4e4MYmqMFo1vk9lyfbnhtFF7h336Dm4n4ZwaINGbfi1JHu6IcGCzvt
GbFUOmPLEEd8YLAVhK6Hkx/o2ZtAaZ+pqenYEdGEsITx7j6O+WzSsEBc7pX9EzJ8
0tGFg2jmYxqJ8yXHiLSpew6RISCNH/KPWicpyf7v713fnpypb3pCdOQcDLL6EciD
EFoqfyPeNcEn8gFEV/m2i7rZtnGPIEGsa7FCut0V/9wTE3kPG5v55K7lO+1KuzjX
MqR4xORrGOOq9E9G5BoTEP9kN2nge5hYW/jyZp2x1S7QPvaAB8NLDLsIQJl5C0rt
ZYNjGFY1xJqTxEyFdtHLFKKnrfpvHNI4dwyOP2WXYuJeVHeSvOQQI6s9M2wtlzp7
lxAL8ZcRb7Qbrtj3/0KRwrUXmbMsH6CnjxopKQeER2vJfQwcxbD1OASGt7Y98mNE
ZldlXT0XVl3lW1RaKWMEAg07y08ojl7brra9lOIKWgqIotw2ot0eZj4TbiX4ASP8
7kh933D22oJCrecQneUTBm+U4lNKmu1ylOcOG37TM3EOP8ZTqLAgnendFu9BFSWQ
miZKzNo6SdNU4/CS/M9x58dmgi98RuRWDTAjc3hAzdD226pnhTub+F3KOUWjZ63r
r9cLQx74eDwIEdI56ztgUyuY2u18cBHtgQxCg1ECOCsvNGhtD16K8WHAWXO2JFGw
fYN72VEcWP+0VS5H2CpeCTVmJzqQH1WcE2Cx0rbGTd6piES0kiJ3QTZLtSkf1vLQ
4Ejbxy/QWJfdwNveSChRkVmpZqOxlZxdGWpyflfc6pyLPPdxGnONQ81fiz5ojSQP
`protect end_protected