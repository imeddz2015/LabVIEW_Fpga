`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 26016 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/9huKRhRMtvnNqb3Z+UU7TahEoHV+T8U3P3ufru7l1O
3DlgtZzb9QxCbOjthp9+wDkjygH0eUfDrEl1ovhZG63Vsj1nmhyW8fk6WjiNTn9F
7CHx/T8/RKne6jHHRPWQmR5CQXqq6lWfx5/ujn5e2BeWvDAh/qQA4ORV2MwIhGwP
ulrH2gHyuohq/XKqpAaBEDyT9a9VtOu4heIYRc8MyggGH1bt97TMlxjEBxvawzrB
GxCaZy4549HMQEbLf5y6vPGtzw4AyzScdGxIt5TCknCd3LD53VWgiRp0xSPQ8RkQ
CMBfWUSugs33rIksSmBwyDhSYTKCmhT1vHBopZWlPIco7oEQBOEhKp20ie9zDNR2
D8k4W1iFzjhw1S/zuO5rAFT1rCfrKBOa8SZuOUzF9qrULI6Y90BqWbLTwiHwsV66
OSrgzUtMXE+pwInENALrx+zPUBmFRtYdbilrO5qGU99ziEsPn952f0lToeYloIYF
WnHEDf+y8wKhzbL35bFZLVhg9Jba0bkcfgCB77t4p3tNFvaQ5pNQZi2yo2z6Ee5l
VLVUF5AT+0gp4MDf7k5TMDHBjHo9X3lAJYL9IO2FAzWE2Eq1HktdCXgAuB+j7lo2
9/JLoMy5ZZ0dpW5BfFD9w6R9Z6iN3rRSBAS27FVUNQiVa12OgXD2wZqU2DYprXzm
1Qw0MOaQVOSYvQs5p6rvspCxFs87crJwQIfb651kh4Wh9Ru2+27x/7YHLxhB5+W7
T8L1Pnnq8kQkTbltKzTIFZOhlFFtMZR5gAIPYor/ppXUuaUTdN3dB8Ywiwc/Ge2c
A2fso0/xl5cjfzndr6fB/KcQmp0mu1/GxtAxmiYA+iytSkEM6iPXFOea0eDWe4pg
ozHNWq+hVoBJiYwpTEczn9239VD8mnpS5PVC985H/d7kVtOP4hPFTy8rR/MPd8Sf
s1R2baxV/uzaYilXMOq+pjF3tbfLttwgeZNQBvnG8k2biwOAaHSRPN9N2E53P/Rf
jeAtpu46gDV+l9o81Z/zN3VgrMW4W6mrzNhSzjUM3HbKjkTNs1rupM9OrBuDB2JF
c6JVzrKwNF9HCSdz/NBFf2DZmmy2NFnpSFr3VzLHSHS26yLRDiArre594+CDJkZx
Rpc4O9y6CIIICsFKQZdNWkLPqGpEHfwAXh/4WufmD+2S+r9cpFWTkzEBpAHp+SK3
Ec6flBheRJs4I4bWaNb0MnLxTWCEEC51GnwYO/RjBlz6WHJeJbj1SDPaMm0nFppU
JBs4Toeaf1RRFMhxLnUG+l8VtnZy52Ab29osUh6XArpHs5BwjQrI+jrS9azYNgOP
HrtJygGGr0GYlz/QILz6G3lhpd15O7Uhhlm8uSGhbOsbYCijlEexqG8hAH9wEUWn
YIfYkunk8WKKZC2l0YXXIz38ME9c/s4bbFcKeRFC5AyK4SUFu+pj8TuCRMObG+Ke
eXPnenxKUL3zGj/i12P6dC3pe9AwhZWqQegoyFqsKKUDLE9ikGZr7sK7otQZEAkm
DUqs6OmfLJF3W1Fh9OPrwqbGqfJlS8vN8oMbg+FZJmFFekMhqmaZXy7jNr9bJMfR
4H9CyH1LIAiScfqXMZagkyfT0EjXISn/FodEJw0h+c0RXQuDgjbP/L9zGk5hl/Tq
MD9laBP4/bu8/HoMHfgkGSIfUb/df1ouIcanrxM6HWr9FkeMmVyFARFYcH+smvl4
8Z//XSxcxGBuRn8SFmxtwZKFG0qFiRK1XkgJmwEFcJTds4BvwZ9eT5a3mPY5BDAS
3ObxrID42gkeiDZfXTJcUfGxUX38RxWUUPytyRwIKwS12AdsoDRf2zaCwcfPBixj
TuIuoXkz+C2ixBKNn0ujcY2F758Iru9mrAx+nXn6H2m4K3bXnzoWJQteyQY2geXp
m2Wq5jbRUCh4LQWtW2iYZkQ/xhX1LZhJoTh6pvkcaP8/ScfoxEucfyHCuU4nazIV
Zao1QBnyNA4H1jFBDz1Q2+Kdla0mtAktIW6h/mBqb5Ha5lkd993rf30eoi915s6s
k+CvzKIX0JxYtrllOYR29KfBaBurJrQ16POGPL5E/LWH84/S0fSiYY8pbD9+mTlg
AlsjjyZetWHoaHWDmN4kYdF9ZW/9wYo/xv4NSOycJgK3wivXu29awQXtXAYGAjeU
/N+yBnKjjRTfy+BaRAYxee1QCFKF3RsmaSpJo448kzd+yM5JM1ly3jvM3j6rV5VE
sBVgFfY4gfEvyeuKY5x3O7eNRrcOblAx+f4CL8QdrezYHvtt7Pgqe6jp+XlprQx/
GnH5f54sKX/NBXOzPAUQfqOdmzRPrh4V5unTS5hHTMTtqccSf4gVjwPn59SF0o6R
JkdX8w07ETsPBH6VP/1qDStqXBtkJ0+q/2niXvo06sFKMmUU7bcMgdSkekClnJU5
b13u1c+6bO2Q6VeGq8HjDTG7DFnV4utu06uqlXj75bpmGINvABv1RTFcPzB1WB3d
vavDYgLO0+Ee3ADKM++d3m93VJFpu+UE5Ky4jvvP7UT/kYTUniZcOtczCGyk4DSa
QCVy7JJslYT5QH6GoXaNksFVsSUfZ/1eGkaDGgmfT3nTvrMr+KCyqN+YLV/erZ71
DA6c36DIqGOOeJmd8sK4Gf93SFAdN3+7cDPanb1pQQWuPI1J/pvfzJz1edp1ksj+
Vc7acaqxrmU9cr+aZ3dVP+XbpvEG8cK5XPX4siP5OwQ03bTChFZXU/4zSqVIo410
kqo5vv/24LsVJ4h95IQC36Y9bba0NWvgywptqiMvl6qkryI3aq2BDcXH58o8ahuY
vLCe3euGJY4EwFW0itoDmMM2nceFEvUoviEDA6lFlb8sXRZsIoYBsXGCleDOfacr
oCI7jN1JEXyICJ67qhhlsJ0ii4fwiYr52xTvr3UH3MzoL6XOVUJuLrCbmVyPecLO
ysJI+XUHar2csuoiZPwfePqLDeI/vljGk0i9KBDvSvpXxk5sP+e//YlIYZwPPEj/
Qx9oZ8nvAffu9XJhjOVLyxLgFSDOzPiOZY7QKNgk58iFBsq3TpbJbZwunvlX4h7E
+1+BpmamrVKYoC20zkarZBgNeMJ+/Ih910cdjVF+OqHfscUnITUB/tJtX1e+Z48a
w7XwWMXa9iotEOGQG9SdqCacSLOs/MpFpEVXBlLc8tJ1LR91c73cyWVNKlAwp7Zb
5csymcIN2P+Q758jk6US9FuvJgHbIaUrSCkEjNsSnNX/MnhEjSQSWbosCC2lnCau
GrtaXfpO9BNIUO3oasQnurXpvj1DUnHgq/Ts/5OtkEBiIYH/e0iWNi9lu4IglT05
cJaDSmAsNtDWIgSksa54sEttFMCxu8Mr7y2rMbcQ1wiJO+BHF6+F/1LNXkIG1ywI
6WBzClKSub2H1ZgoIPVrZAKbZHlyl+SubW5iXVmfig6diDZfZmF0uCkDtUoMMzm/
85gEuqJE91+x93sZcT9Z53ihcxEk50Wt9Bf3tX6hNePfnnvrJ8UkTO9XGIYEqgT5
6Vqtm7t6of2LnLlqUDlCrKYQ+6oxsDmkbb9mo70sUu5dAxni02iVuXiLElJo9wcU
xsVFZPFothQxi9Yz3+0Omm3WtQiOOz2zYEtA9NDlSl4DDg/zbd6ic20vsp+RB7Tq
yph4YVUS1kXzCoxJ4wpLT+rJyzcao1DWKD2NZlLap7uy+7N5YflgJBt9WBAC9fsx
kTIg7k2nQeAivPtzL06/aSXlxi2qUalmaSkIuB0M2ns0tcFG+5hBfrAwUYbu2vU0
pN+kmK6BEkfdmb83f0wGd4BFwlZSQ7JWqTvrFlcSPAHbsCZdK+9/dYJxhWBv6Vid
uoSGeva7OfpqiZEWR4E9vRnb0EP9e8AmnzuZh+5w70zg4Vh3AYhbbGkFBw8thHhQ
gBxMbeG0AEiYsLtMCo5wyRYs0Jtr57djrBz8erjP9IVj03G25/zAzgLGUCrmya5G
4lmnuIRJzLYNEwqOCGnNSmC/XFDYBmktyS3/HLddRuPg9F3ENy7a2iL47Cwe+hD1
8alVl9XVURkdxLsHS6GP6FrIUVAobNj8wGOG5PG04kA6SQGIrJOv/Ncnp46U2GvM
pLKOIfYx8qITnUkAjOFnLTQCBEIw+/tVuKcu2XThq+kq/ywSyvZ4nAdfHhINgop8
Zponrt2SAMibiXdTSL7FewubxXzmjzEPGBCEPxvza58NeyekPTgj+DpigNVGXkr0
NVM4vtvRPSgjUYFvopU8BmDg+O1Tc/A9N9MdPIZ7FM0ECMvSkt/Bvnp9AgPz5ed4
RVioCWv13f/iMQ75Tiocyn6MmK0W8ApMuopXV6TIIsnQ4gP+FVEBoLTQLjwcLhjD
E9sD8/yqQGB0wXztd42hq/jnIXXd+iaprCKP2I0/+kB/X/lgL4d1vjbVOCQNVo4n
JpRua7SwGXy2r5jxp1A5fkWWeNngEYLlZIOxbprHc/J1Bys4kr4ps9uWg6oSA52o
Qgfl8UTzaUNr72o2HilvtnIgobDwhd4myTTgH0N8vUniGBTgBQ/1F6UmSI0se4l/
SztmbaGAElp7FfPFS6cvNue1aKNoTiExfcNEY3ZVzDlea9pIUx11Fmg2A+z/zz9g
YkCbZec22aYvjf7K6DwCLKlIhQuRk2rHaQa8Og5CtPNAFhJHCNG4f/bISxBnYXV+
QMJFE0JclDApmBDerqTWoW/SoclYlzSapx0LMzV2qChNuTOAM87VlIyL1dCOiIAA
QkDvOMhjLLXXZSRDdhIHO5CwqbXIdFhuAPx2Zb4Zy25DqYgtE5gRrNg7YPb6yWpE
i25mk6vT5rUTXdPeR12gcm/lkUqZaoN2uJel8SnSWMTucw+B9GZeNnGOUZfrvz6B
FmpD7cog/+gRNW7m6vFzl1h5K4wDivrGiJ1iaaZ/U4BAbnT/OB1NhX+SnNcJeEHI
H7NLWTtcvPYg1P92i//U3XNhhkioqqCaeDks1IZfIWLO89zqId55GI8LKR9ZFYq6
6CF9Xq24dKaAVfa64p5RDinrYat4BTivBr2ermakg5E+dee2yS3xkN/q9hHc1rgH
4Vs+IYBiFUjdkuc3+HRriHWB2asH2kLCOZ3od5cmQAObEMU02Ou74ULOBVhaS1o1
NNkU9UURXV7FjpNQgv/ZKnOyyrJR5QV+J3B4I9PulixarEIIiR/tA1OG8VZS+oH7
nQugVgt23vSY0OJbaYyYQjQZM9yo6K45Bef8C8b861YH0tEQGs3N/lJgcnKMyJNg
tkuG8gdJMx9GQ6WDcaP5XHNWYRbdeiHiCiRsLdbXNRzHZ8cDfDOqUleHLwRyHyQ6
rqx/EDCsaIS0MpxNIxdT+pojWS4dkoAs/KXsbkzegPD7Xr8g54dim29lBCEO7hPJ
IInuKyVvF6p7VdqOkJNKyrwN4H84S1cjPjoPJTlxCYp0fEkACy2HzwGQSuJ4VjOV
ssQd40KgzwC+7aAtnL+3/dLd+aLJp5QC+8fNJepHbBiIcJBCgbT19sEMZ97RA8At
AHSby7uU861REn8ZBEKVimBdBz8DRiK8WkSjpkMSeJ9R2CSc/WInn3hZt+2258vF
RwX9WWpB1JGhZGOyVWPn1Sd9TznKcWYNdKQWcb97thQvR8nTvD7d05Lt3YBwQn52
dcfsAv/ggVLJa2ke7Xsx+E2dIjf5VlG8nLxzYOViWPfnmCejjxHx+fHxxG5eatNG
oesRR8DdejCuhGULKtD0Tc10et47c4jgPrcOwx2NilKW2f8VxNb0GzywsQXe/djd
uXeHfLsKuq90vUmergHYL+g1C4zsh5s+JQrjThEzIOfNA16DjO9JeyqaF6qJqRUl
4RsPj3y6ez5zhOgcwDrABDHGjH9DOLGXQu+sfnkk823J+5rZ8yTmt1R/vmuuUtae
TKR5Q9a6vT1iDFB9vLjpkOWBilurJxHFllu2S+2wGGkRgj/aJ9/WrPy62JFbsqi5
AzzVueertyHyNc0nHCHC0++D2jPfGmzfUXF6JWuImIBhauey4Nai15HWvhboevFJ
9H3cxG1U6p0bScZY2KfRlRUFP70sD7SPzxzYZUxU/OAI6UmhIQmYsoWzAtXW0rXF
MieBk8VTb+ebCXndeJhYAjqRIhBHCr4IFjRGIDntsFQ0go5GvqZOglO0T1zWn4sP
WMjiSPoNLMblW0oToQeTS7ZF5yTXr8qR+S+zhcnjpk61GWCoRM3skQchycSx971+
WtS7NHFJt0U4fjH+c1hJZxIWLbLELirNm/gjwG/RBUPnwK6+8xE+YO6GVEtiKCm2
NptweP5GHQooqRIsuqe5T5lILOvECWfPXiq1KgK5/iQPFVPmFKvrLh/k6ytUzP0R
6430Fi76IbDRWNJGtqOEV7/oCHsjr9kJNfH3enF6JuKT/VpYaJMmlHYfxpM1HFba
aagBzpT1DoZDOY2zjki/i8doRS9QnJsYvLchU8f99CZ6nQIqNDp7nnKX0NJAQXRk
sdA46fA4Iog0wxkqEH+qTQmirNH6Olh3sozHg9NWxSgxbm2Bz4Zs8LHrk4ybBLWL
lkBMtZ/8IrU/GtZa9qunkTk7N6PAz9+woCgE/QwDUqlJmrdjCJP0cWH0yxKaGi3L
LSBfWp4Hyn1ylIi95yQzOG2Ig/kAZdN5c4g5wZ6/V7CmoSYFf3z6BiHtXAyWOAj5
0D1pRoF473cywAURd9TilQaf2N5sreVQNK6XelqI6GN6rjTpBExywARr19xXay8A
bBw9OGCoDTbpOrMw7bwSnClRUAsA3CcPfYHwuhTbMv2oMVnvdvjoD0CvRl5QoqNl
aiLkWpElUAwD2VuvFKVVzGYI3mVh5pK8oywSscV+ZnrjJ40SObNd0H3qkCDMNaIQ
c0B4xJnUF1s2wA/9B8oxM/QcDDW87Czlh9lHm/0LBLaHNplCQy3ADTYct1sVSR7Q
WKHifHOl3tCWNDUV9oJATeulghKfkEV/cmIKwaAyKvUapV4bBiSFe0/xxddlPK52
7FLV8nvHN3ouxzVebf4/+QnZDwCURzmxgcIXrfRgM1T8PkQJZgqHAmrkWKKJiBUR
2R9pmQsatFLFWI2dcP4yDXKzzYRs5cAJDcj4VLB+uy3LrYWEfPxA1jiQ3R+0MNfQ
fv0/vpK4NF3zpQAbN/MPND1LKE6IGTAEFd+QwtP0+R4dcfs97k8NLNx69/l7CnfL
W9f0BzaOEdo6sur1CrvDtgfsM0CgyI1YgRSOjjkALO2VgfZa43mxq0EC4iT5Ffdx
PtBtGf0cegm51Lpu8MWdhMIxgXBGsy0yVlOTgDDmYRGThyjIlsFze6NAoLFYCrKx
itj0tfyY7ow7VvtlmHj/NiL+X+LHhCxvvbYAg31POZQIqi1KxRjKbhjpyz21rAMQ
pduREaTPdFs+VEPNFr4FD8gdotXt82iuHILJcLxHwVcur3yYXNGqTqTOulGMyV5U
kUycpx7VPYnlBORgHPNpoI1RkE5uxStTNZJjW+P4G1njrHiqRsL7VqsDQq45j+Kq
7416bg196Z05dMYTu8szRK2VW4O38CDWBIN/qLpIxD1s6KN2+ABDUy74/HrdvZKD
qPvnUzD0y8Olu896CfPmnWuwcbcHdgO0XYjcy/xH029tMniweYtXlXj8hWyglh7E
fW1V9EPL9R24mcI+JQj7Fl7tlefU4gYyeo2TwP39QnG4oSiEaoNE2V22Yu2mW3Vd
5ueSaA+isVUSt+0HHHP88WyYxxss0+uBWunNTXnqfCX9nWYt++pgbs/1vHIaVonk
N5BfJTBUKh5n6VJzFDV+XY545EnrKILflSRKbmj/Lt277MdW/sZlAePVHzBxHSLt
NsezrZFBkMx07Z/h6S6pxzZw/RhhdUOPUYVkbXwlfxNzDG/we+ueFP1VSlvRDHTu
b1Q5rY6jd3PjhbPjMp1vdUded/mL6sFo9kR1sNbAA9pb676nl6zp3B7DD+WOzFOG
/YlfkHdwpMaKzkMFN7lx/tDoiV6eA2iq5NaVnJHCrpJnKTkkj5opY/fanZcwSfhc
ZlKtRQzrSHxzAcE2sJqdDqCZZ3SjsIYduHKyGvkykqLzFvJnsvX80Wxgy9oRBNu4
3HoWCAR9QJZcBzvawR2nrtxm35fA9Q0KnVUxYOBfkOw23iP3YGW4TOL05iDDUXWl
ybeHJRzQY2qyV/1Hk29xATTvuI1NNM2VNzDDlrxlhV7SledzZM5zBAMdlFVhVYna
qqPy0jj2Irkhzt5PqtZCdniBawVSQViEKok++tUClSYqJPUFZco3ryBpntlpXJun
2+0xb/XFYBwrfIauzX06O8W2SJwYWOdOrRsTIUuRGdU1LhU23F/37F3m3L5HLKjV
AK3ubSBwvik9/Dac9XjNCRw+66wkikN0a9/7oNbXVtng3hqxjTE9HLGYFJoINmnY
IzT4rTpG01K7DykJMTImIkz7C4sCFF/Sv5j2HJu5YZV0q7oN/9+GNGvOz1qIndVk
6t92I8xA73a0U+MERqnMazq9vdYNUg/zGVIGpT/s5TvhxGHsyuhJT6E7NGuUHcH3
eILUXxjWJwu6tQU91wyk0USw0yg81sgAKRgGuZrJDwyn4aBtUwzJ1LAOJDA2QnXE
fyGFqXPZWAb+QtzX5y0tmxbMiXVNQvZS/NuuNeEtMakTnAy66IOgjLhrZyB03Huu
MQwbNUQV/k41oTZieD80fz/9mNCu+g33YS5bpGKiAFvHga2kjz728jB0RR66wt8j
9lLv6xX0p9JzlOVgtaBczbLr7H7FnBykT5g70cD2zQd4zGTLfU7OumQl0Bf27S/q
BXA4FzfDTqnER8keYmRNNrZHq5mNFaOP6CgE21FAa14x7kKCbXkK8+Om3+GmytlC
m7IXIC3YbLiE5IljRJVkNogkmdcYAcgGEzG4ubzkKk9fCOOReg8YGd0r0i6NoYf+
E9lquc9TMM4AcTEi6anrN8wzdQWEiW/2b26GgcpU/FqyxeNNtUl8BnFjeYPoOXdG
gML7DMk/r1xdDB+QmGenWtFJ4CCxbtFmomse8bqRAXUKx36e6epDp0YnyJxzZpN5
i/tZ2v8bmAQFT51h5Wd42IZbPwruTNBy1QXI39bQgDkNZLlqA991VYcTg406e9tu
GinC/3i1MaCYJ/M+Gbh1d7UiaWvswboB4yyyh6iNfEFwpX/ljqV3yZZswlIqbUrY
ofl/HbjCGCpy1U+UgAvnmoQZf+uRREsicPJLeYyI+adCJnK3wihuXds1XOtCqiHe
sch5Yz47gulpMECRMWW1SO65pDyZs6YMnZgxwbzf0Clwm03ElYsNYqy8ieuBa9N4
FQw/WLIiFtZxHDDChwCw1lVC+aSSCtIAcEEIkq5twx2CNDy+DqnWnYt8OSySH4Wn
fvRQgR+czXhUVFqxE168aD8sG69EMK8y55KM2Ng90ds5KmouVszrRhR3KtDB2/pS
SGDKvhRWR6yd28+ATADlmXHCk4HeIVjo98FB5o6wD0oJrq82HpH4xSXZ5uwgvXgd
V+fCvxy/OYyZN1aP4Yv8SaXeLvtNENj2k3jLwLdKIwheyYQbMoa4Qdd7h5tPOqJf
VOBuwVEfnZ4vrLcGzcjSdrIQAclyya1nnCq+hwVhU7fOEBSbxZ9/T/glQkKR0G34
Ehp0BLGJdwspGUTjv35OzVmWRDHXbsA89aqoX6bjo8muKQEC289N6e+z3oMCudmW
Fik+PfaFn/PT9BpGtjI8/2ihM5xcq08E0d0BghE+mP5XYsSlH5ZeodVb+hFJxMcK
c9uxUGuuD1QnPvSAGdkWmpZrunYUG5OKxvP3/VhkK99I42+9E/vwn5CcFl84AV8E
+Wj0xlKU8M8ILWOU/I6D850DlZm9XW+H0tGHlFmA544aHWas+FVQFW0QmqunnZzy
IcjAojjmbW5/aZx0+st0P36REPLL1uIKrpLaesTRUteQvFIO1jm7SW8Pu6xfjK0Z
4Lz5EHdzgXJq66g+dpqyt033/t443vgEdafB1+qtsceu3iILYHkjaEjSaVTNOxvM
87bi+eeG7i1oIOyoyasOLh7jTJZJybUSQSiKhQ91rxIbxudEtzqhVG7jLv7jyx1q
GiDtFku0IzUie8zzNwCjvnP76WMcIFwbHA+Q+0gAaoCW9alsh4UP0WkAALGa1YF5
VA9xL9T4a49CBmUr8G4VnU/50BUlGeKImL4e1mndDULrDe30L27rrRGHuQU160HC
vcC+lu/5vuFpDgd9YSjNhGqzz6SS5gjX9cjoySbKDg3xoz+ZlHgY9seOjUYvQu0s
WNOJbqrKFhW3jEKisPE1u/mqzSiM558omuKJXigZgtS9OEZmLL7YR/gtKAoJ7UTp
VPZUBU3KCdrFg/l0Juk7ETA1fWOuegSFVsXmVNFKYtT8xwYHGoP9RGV+TKpzkI4d
9qTBfv7h52+HxcnrMKLLiir8Xsl0p/s3/O2JRK3blIZWdXCLIVnhV/MIgFEsbtgy
7HtsXKTQKMHW6X2pJfXiZc7PNWReslBglYmO7uamyaLII5NXi39/R5fswQXU3HsQ
Lwv2EHI8W1doxdaRxceHlPNTPm7RlTI2jhLMJ6Ak7PLtcLn1TIfiDpSDDhcfOyb4
nJtu3gCjsW36w8MnWfGD+CP3LIWYHjBLDLo3/nPsIcQdMKcZetZypHY1ijs9tgRc
AjEdz25l+pJKuwFr/jOM9xvlMAldxA1VKbIGK0f47Ojaw/ZW2oHddZhBn0DVccPS
2jmujWHiCAV4kx0GD+Q32NsLSbZbfqaKVbA/QdLH5CZrJFNsxQU2ZutH4pDnc0GT
CbO71mDZ/oguD6xHth9N/rtWW0wXj80UVrn2pAsg6tcCEvyD3/9bS0y/H2CCA0Ew
KjSYrH6EZE8SFOnx5GJOYxYoUrAqAFKQ+oz9AXFs1/wWLvxUQ6KhiByHGMdwomc/
hauLP6m3lgM5nVII99OcpIy7LAfiRYlbgkPNtyOQSWGSo7/eK6KqtGDbuQfurupY
2aSREUk98LXvYKy5nI0Zg0u/6xPFK8WHTkZ6S4JP+jG0mJZ9FhBlbp67QuRZu+hw
jynJDrGXkcbCsEBfCj3eYzjz73JibtaB7Z8tRjlybQxIrc4wNuJH8X5D/PXyI8w3
kCdn2NR7px7PkFIJ7/raiaBTVK+z5MXoVuqbbsk87sbOslYbSqoypCr9wcUjJ/kB
q6eeGVXdx7zmY9Cx/1OVkROgd9oKCfzNOQEoahmL7fDPKealuUuCSSFSjterHqFW
bBAkpj/CVL4aUJt7HIocL4Pgjkw3679cfLA3w9TPgyVX1Fy873iL/T4OXESnJFqa
RBhfKzJg+s62C5VeKncIik4KiQcqX0o5tejItYherVS2ZJt1M//gPYWCG9JLjc9t
AlDE00t3zieTFDVFNiy0JgUJxO24+BrluPmpthvQgmnqjWK+XeOuXLFyIqZPDj3P
qp44/elYSUOJ+ikg+zQSUSqR4Aw1+Acy5nVmWixBPuFScLryWLDsjClUPB5w//lq
LGMqnaVKVpvwrkxaLdRLARrr10LCCmMV9WNJIxpPZ9NM76VnV5HqM7NHf9q0WSRh
UW1jYdPXM9OhFayUPi/lpyd7Ek7q5lUb4sRaMLu3i8rwi2h/P5f6SMLJ8kDICdZ3
qV/Cp9pa9HlcvooxdFBCUgsOoAns3MJtdIFqMe9hY1cMXxIgqKDCJS6szjdcj1sX
93PW8eL8VgY1EqXpIiWtuO/I0VEPvTkEiFd92zCTY+tSsfYfIOELQMXVhe85bO7e
DluOKHwbb3l7CnPjWXX45kkY+054B6fEAySHXBqncrvxn8x4t7o2T6H1GDC8yYEV
rTDr/3xw9H7ZhDAEXck9uYYiHnYcJe77pl7T7gxdHTRh4DocZFPCsCbdzqaEeUMC
Zpgll5LT5XuUEXKOKIbjvIst3wezaw0Z5bRgiwRlQmyXUzyA9lgRWpIwqe10N7i4
TI2MoS456O2qML0oWmNnLshNGOZVfht3wGP0wtAA4YO2KK6yiCMPTwv2vmU6yrlm
CF8Qk8/u0YPsSLKBO0g5+0Voh4RraOfsb+Icy6fo4o8Yn9mt0yB6M9h0rzuqjwk8
QM3OMdMC+hjVsHUFnwibMvxLR/c9wgCUSnGZk+t0vK9GGrHBxXaMPf9M/IKchyHU
5xggqpv34Sz7OHFU1DRfjojk25Ub6Nv0FajyQroUGBOb4OVQjgtDrbTmbMM3fbjf
Od9fjcdnI4LnwGhlHLoNjkkYdaWpG6erARN5uJp3/B/o6GdcHKpy8pWzvJbjats5
43LHfBv0mgj07jYtncyOYlW2TPbJDKLpKNSMQsXJSVVN+4cUPKDTneccLSwnTXWj
OKbgKSUBGF6e5XxF8/YbzheEv71QMYNr0krB6SiHvH/Qt80hgv1lYhuus7FfExix
awLNRJzw5m6MW1wasXl4kOfshsu2kESWC2j8bAwVA5imB/otSU3d2o7t0UKtUuRO
TmzsdMckvY5jKUW851PYf9iJMSvULP7YnNuScuI9SrLLyAsghnDxHlukI57ZrlJp
D6oYVdq7vwX5I7KY+HOoj+7gbfuAax13emfAn31EjIfFWRh4cTuwW6BsCGfOd02o
CKtmiQdq7HH+kA1pD9NMHFZuvXeL2U6XsPJNyX6vbA6Y6Rpy4nYtai5pkpdNaBQP
ojYSxRG34zmvFclczv++pCJxcJ6snDDW45el1os7Avje3j4sX+XoPERsfThFGV8i
3GIe2q47gW9TWXV7b8l+5MnUVtTZaWCJft9pTGv6r+ic1wh0vC4a/tst1wDAV2Pi
yYZh24nj6KMYJwCjSv5tncXP+MV/054crfam0MgKau15ZW3N00yNA2lBp4mgElNI
VXlrYY91G5qHnw8FwEo3d7NHmn6U2eL+0H7ajHhgL15aBO9b26xtBvo6WQFW45U9
BZ90bzIceO/x2DxtfooZEPlKua8FG7xlnsWF39jRp1LIcjuzw4R9ALpgfxNJwAo2
n4EH51YsvKYz1sDOPFhp8TJSpva6zFTCDilG64k0Cj1kwpQbLlrXbkSa6BnTCBfC
reqU6PeMP2PPOeD3Cp7GCWfrKUOKQ/b05c2uemcnaijlrF747f7a1nFwykyjMuB+
TKqP9x4H02+ksAzDczp2gjwVc5wJMoDYJLgIBnmwqQa7GbnpQV/Qe4PB4kZwYWbG
gJa8t0iIItoUwmNAPLHMMxTyCLrEVONbcwsQVy3KatTk5+gn1/ioaw0qioxRx7P2
4n6oMoEtrMf6hGaBC1sS+N6YwaZpGVxt4IsPkSUzjjJ99jGavVtJT71V94uCwLeo
Ocr4z810g/rIOqUYBzyXvdiRXLlU+bmYZ5SPQOFJXxIbSWsO417xUoUJuVssIuS2
OPTDI82PH1z7GpSmPgp1AUY7a5tFPZfMUjdPnXAxGdsmsX65Ct0QGnXkJM8ir/d7
0BMN/YMsJiOA1VF7zjd41uQEclUIAI+aj2B6CActaKyTQUOkthf8wol5VgU1mybq
gaNZppWYy7ejkfNclzWmTzYuJR3GxgR7rFBPxx2Uieo0O3KHLRiUEMulWqqXIAry
DCZSVGXhiydQuwYIxUie3qB02YFO6+y62uIE8azwDKaqfiG2DnTktuY2Uhc9vDCU
r8NGx8d3bt8NtVelzPLPw6dRvY9k/+HurFe3ENv0glgOhI8Xf44EC/e16Pyd9zSN
g4e+tqNx5Lbu1ExRaEpWCmcyAmH/75FUIbir+kFbZCa3Y/og/CRv74nseHww9umE
PGfTYI+bLCcZSIZBre48tdlP0cDgKdQKj8yL0che6RucWZQzh3w+GySUgzhEfxBP
UJNY3trX5YN5IAZlApiXppA0lLu3PJEom48V43FSdl9fUmiEvo0UrB8n6oW7QpTL
3Lvjk2ITZ5L5xRR8v5looh3UqXegKtK0k3SpeGMrwMa18NbEnPIUxRfSAi/UUqvp
9EqqtVpB2vKscsjOmwHFV1/ObQMqj6/HDieQdcTfGqBDfSAq7DaKeuJ6XWxqOloT
rOX6VgTqRcLjWSS4d0ZXLHg+Yx8ry9udxjrVIRUBnSi5P3L9+RD227B3YrKKTrve
jYEvQjRCPEcrleVKbaDrPm77b9sjFFxGGq4K80hCc0SZdaBw51lR0uOA6YARwy9c
4NeFXifZlioV/xJOVQGXUixKRCV5I/em6XfxfAkUFQF6cIMN1TVag84fsONIJaP7
NhSamjYx98QpTf8Pw2E2s1J6AEDML35dPTRPkhkvZrcsl2gDgI3cyDONqv4nzOM7
XejooaSTYb3weIa2jtlckqmBXcvMYgHq+/UCG0dvbsK45ac8QY0q7X3X9pRy7Pyi
nZxc5vIEmzgbo/OH03sLf87klxvH/6KBAfFDQAI4hOKT0ljNIGYtimKMOC0YHf+q
2ouEWvDw1mPz5+WziLzEMXWncta5Y82e6WWtaHBfn8rnLsBpu/r83cYaOcOmErWP
I0nzDMm0odvbmPGdmH8AVy5IXvXo9UVVvelUw/2xNR0FpTlwph4nMF37GNhKPcyC
sUVBycMrUeSZurmhynsXNt+6L/gdLTV34Oz8A1sqFbFFbKp9xnCIxhLGCXJAFhpU
UNgJPNwv+lb1Vqgt7sSaSxa2VKAkgz/VqTukeq3Tv5Ob4fkPMqxpWhRr3mCghIG/
NYqQ+Z/hphAA789ie+e3cnxcCCroImogw3VKyVYNFqA/FGVNggk/7/OJ6LWkoBox
uvnA2T2fCIwxfr5Eo049X11ioGMzCs7MfNWBFvafHgRn9RruM7waLy4fAPRHOYmG
Gl6Gf3mRVaYG9CTaTRd15SaH3ogqFeynkH3kgzv5BsekF8E16lbNyq9Gg9xoJhtL
nxkLV3JXReBQlRSPqLwivynYDS5F9GFEVkqcWtxGA+ZOXDp7QIkvcDMy7ELPVZrc
M++A/Ze01JzudXsJhHOcrxB0oguzGxr+qUkMNNiCrQq0d+2esy3mDwVWVJ6d6Z2V
XJ2sxw0MTVZGI0MgGttiYODFtHQ1IuwZT1G4jOpnJhNMFPi+IxUba50uTnq94VIF
4lH8ZZ21CawGWN9DXhAARpI2m4cZSHGY2fF2B3ew+AShgESakBVszcExiDV7KrQj
a5BMDDi09uQBJhP+yFrjHVfX8g2uJsD2w3tCxOwwQpOeGph2miHYTUMYfmx9ev9v
OdGtTDk6cPK6lYeoF6AdcfObpOvXv8SwEw85LBlYn0hVyUdH6JV6X42p/vWV8lGF
/25rZ16ENpPy0/GMpkne2a03Y2PoVTv9ZfVfNYbJejVYEIHzu63a0X4dPCTrlL2v
6nX/1WQHTlEOO3hd5I/sjbfGTM3+0LB6wxbqpoFWT3jA1iz9eQ1VVHJB/I7KGaYL
tlueznkijJTkUwSaudht6JvGXb/8ZXvgVbOMFB3oXU4JihyOohIGChu8CwvHqJyp
+h0a2a3uW+OiKfDoTQO6u1vLy+8uxRj8bNJulYRjB2jI56rDXatacFnwNe2R8S6/
fM71bEYFq/v1wh32odo8Xcj1EafKd2albxnqcCBwRcSjgHOM56LzD6UU7AKGYd71
T87BRBoM2InrYFui/jVNQet20+7YhFmYEW0uqrAeiO9xgr9wiZdSLnaEPvbF/Sns
SBYIFFEUMjfqlUwV8DaAfm1nuu55i+zaaPt9fHTe+ZIF4MhfLiWcgKXRq5EzbiUr
FKicXdk/sfEHo2V9em4ilSuR3O7C0V3CNjPrdWuVTAxLgfBQteT8dHsjOgvnUr2p
U+sTnF/g1Wh9SaYmVs50BYHbLi+gd/HT/pmM6Zic6DG6IA429w5w+SLFMYJDHnmC
MbsmLOYRK08+Xpqb/R5KPcPp2Rl3DUGvzOAQiuv3WvMbSDXur8xKQcP+zNuHW/mW
LuOl5pglhBCCiolwxX5qPYFvmt0NbicpZqaH+kV+et9pAKb7ZXrB1F5NLpcb/QHZ
bkeCMMdDR8TGAehz7KH0VdPgxTjZyiyKccopVPRo9GaclG8EYaOxn4NevGN5PfRD
b/iqRgcXo75OeIGfUxg9omG6i6N8C9qExppDZ6cpxBWXUHheUSnA7fJcfzg+QQK8
o0ceK+eAnxxFHDsHWCbLoXS4hs0McB70gA9+mbECtkjs/XUGGRP9aoOMuK/xeKAF
ZfVy0RjwCCoklq+P7fcO/KaXwzM3DoQdqIEnCFreQ18Zh2Y1jbj8a3XYtakVjkvO
c/jpr1x0P8EaJGlWJGhu0Mg4dBtSYIIFvF3qSugBQNXKG9Ob0aL0ITUuLzIu8Nkz
Ugy0p590kZS6zzUlWmhy0Gs0kW67chzk6+3rxkpLD+8U0tGXU4fQN541+5XA86nX
5qgdA5X6X5e+B3oYSrgFNdH/LwLQAEzkavhewnxcyz6S+zgc54XkirgST6sRWJt8
qtA0sk455XO4UHXnymvKkWNZDUoJj7V5Q6/00nrLNNSd1vmyoarRNn08xOkx1V5t
dOg3i9KclkDbKBbwDtjdDXJWboVCsGk/jYHtkJIrgRg3xs7B1iV/AaWOzIE76+5Q
xRbZWVYsw2c/XFQZmoUa9ffu8fUugMcVvtCrNrnfW+woEzWXAoC3VtxHSZxB84Do
QIN/dAuJXjkxRsLR/jQ0atVbnS9OtrMsv09Nc54g8O580QBl6ywhafGWt1UM1G/n
+459vynY5WNJQXqvzofd/kePVLw80ru8ffMTsxBSl7PfXO4UKrxdSwiosJMDrGRF
rywg7SIUaKH/heMp8VWy9EU0Dhd6rkOvLkFEWqMN6NI0Z3nI+apJmez5+MSOReSK
OEpY74XqsF4Ld2GIWLwMQiZ1OrUuYijLK5EUI6F3S9Y5GyXkcJusX7BdmcCwBRl2
2t0m4k6e0w7H7z1OZDC2ifxLh3NtHLgmaGh/WgTaC0pWZ6/H4hpGaVNyHz2az5X6
NZwjojk4LtWf+6HYsZhgvYCEnWwz6U1obI3bVBpCG8/V3D6OcnGeV94Z7wbRRV6G
1TFOErpFTlqATW4PxpDKWcdDC7B86MkRxFTu2i1ZnI8HRU7cwC/gu7ieCq649Fna
7cKzuLWljDQw9mAeFDkyoLwpB4hoDpRMaV+xAW/mkIYdyn4UBW4+HibCCIhAwLJm
6y5hN+oRs6QA5iyDDnPEtBcOLuhviP5YHu2nKG+URKQFgjWKTH25qldnp5qtxPYN
rn0HknbCDt3q/EAvBx8eTKGdvLUxdw2na0skqDgKviWfuMPrM68fTAw+w26K1jGb
NBYS1NZEXZSKThUwQq9q/b7VR+v3reZSAXRIJPzbjCjjpkf4ZU2r2FZIkFoNLtbu
e3vbgR8aG+9O/v/9YRLnj0rHa1I8VJj7YCC1Qg6MOrJYxcDucjDOy0IAR/aB/lGk
JKg6Ib5itdMmyVX09k51B/Yo1GTUrRWIxoG58ZNBvvMBVtJJmkAVpJpdus+iA/8Q
LtwnuyBNWVnhbdWEMcTjvSYQpe6WANNPGVKIKbzzp5Mn9yJcwuATxEQOVWkTYrza
IU2lo1u6R7m978FEt79ch9Bq/r4ZA0XCoVBAIDSpSFpS9W9m9mdxsa2hxi6/3RiK
fMN/J4ZxLzPPJ+mSHxIr2SnqRhhvJ90aHcZbOCI409sHo1RZPQRHS0i2WVJ/gNfS
uRMDn5wxYWtfdhTX28xYwAF/kCXKNlUZayNFbf18gt2eYa3X1eTu7d1iRnU4k/5Y
t9LfpWOJ2YdTPiBh4vRY/s6rArhykpdacBcZ/yVpnAB16rrQFYBvX4Ryc9Q9TH/1
gd8sDv0Ahjrr3AZU+FZn4W9SXP8W5Z7cIh+NmpptcmAvXx3aYf9pODL66wqgiNj4
48baBBpMCFrRFs5AAFYvSQ/4j36VtJV9f6GXentwp6uYEL1JVnBP0O+bOgvJ/K6B
U3JabYjHLJT3s/NOPlJuxzbpdf+2QLP5srARWkUGARGuEPBfgBwEQFJ8odMH5k3O
MvCCOY44TtvI9GYFc9d9brSPYuL/MvngM0wJCvW7MZueRxwpCuiFs2UBvCJ+WR+w
QyRh6gVzyzezSAmkIpH6W94+dYjztq5Jk09HRF4VRjTpVgCsrTmSYUzMVpi56jMM
jngwUDsOjMwQtZD959kg6OHvFaENoSEuHfBSY4BSVHK3seC+ppIEkLR6KU06PrnF
a8+R1/179iGD0sG3TAeLtwrZ9mXxw+VzSeXjcYN94HquseOwItU20TF8H4Dejo/A
K3aqd/p9wPkyGZ4bXSyP/PHYnK26vZgcTCzBhzHGuIzvKPymfyG5r630zBlkfH6B
1qzKoZSa/rWhcbLFfA7r7c7jZA/9Vj9UADDMP1c/lSimHhk6y5L6XYtCbp973laT
dbNaeJ3TITX647fBytk92+Te4Ck8qLIswYCuuei53rt2c/EJAhAH1fyliEGcrmb7
hDZtmZD5Ip4yTUk8+7n1sLOQvr+YzL4lTYlzPU6TjAaCCn0TNzgqS3/INqDkGW+9
fBQCQ/rDbtJ73kn+SEHi9AoG+9PDHPotlTdV60VL0GqyvSW4SoSjtJdhaj+YaB9d
9G1Qg36ZGKkecEZDmzI6w36L1K8aNd+xDIOT+5+WOH3g2z7A5j+n8BN0m0lKKkGn
Blmlcips1/hZfXloq94e44cEnW9vlg/I3IESLj06YzBNcOi5HzjvKwJaeuTkLgui
S6v1Yqs+zHfWZnroqYcjLAIwIdeyfYut6W84ieu0ofuBKIxXXHN24DesdCR+iMGz
wA4XQTh54RNidrtyfkDYgAW8rWMcuFeu9UbYFfl1geEpsX63XXM/WdyFKDRVsIav
LPtRJQHFhNZTo/678GJlbbFoizkpRiVRwBFnbbIsZgFiTK6/ncx36ZmFOWfg5rEw
KlUBc7YQwos8aUynuI5rtCcP3rDZQnq/L2OkLFsP99IvJsfbKMwWzj3emTaKdG6x
e7v4BEJzO3sKA+gvUDH11YeV2fSelWJdoO6WfquG+t2BW7KkMVsP4FWkMvvxJuq4
j9GWO3SsQCznV2oV6LPm9rM7Y1lIAbrjivTjCO3xQbXQEAVUEY8beeaHmH3L+8Ws
5Ooznch3k4GUWwFK3F6DtdD9QUk9T+Fg8WzsRTG8pB04UNFMm4/YCXkisTdnC8Zc
5YKTGQ7JJYxrD9U0xKgEOO41OoKRom+CSUnkv3+fOvWqUJybuZGg4Z9MNTVC7FxD
xwX7gTeyX38uAj+kUP4vXHABElc3tO29ANbQlnLGrIqXjvzIVV+n0lUxxy8MTq4G
DLGStsk7wl6TT9j2RV6vcD0C+P84Cm522B0KbBiQ1XgcmbbsTWHpsrD2sGK4+J6V
0WeInrEm/N+UDWjM2sbzWjAqYprxN5/5aiFAuWvFWQbhnILuLAy1pZq8AkKXhG03
Qlhru1noDpFQODjE2HYuZOQVe5q3W2y/28q5IebMsxYkZFk6nPfEFmndxiRT578L
/6y5e7awoQUtQLTc/DQv4k9ZDQO6q72n+bPmIaszIFQcsvZ4Y9VWmwZQITb1HU12
rA1oQfE3lic1cYq5Wmmi06KX/Jt/d8ejyCCKmutG1c8CaYIeC7ZG220tg40YB4XG
Ms5N53KmAE1cX1qW90EteRnwuk5HfnDAy8itVBAKLJcRLlytzet9LD021zTygE0b
aTIklVcjgx5ITdGvFN2DAv/COXun1uQoDBg9AI7CeGpB1w+npl76yINrKlcF76ln
9GU+EGGMCfMPuK2fWgCRvrhFLpp0/0qOsktzpQvzHPOCjMrfOtLKPbwB07FgEvOB
+JP/MEEhK0vQm4pEZl1lryjfYRrKQCkGZrXHDOd6Ql9oeFLEkoTdKdMtZLU9Ty8F
IZxHjyGvctqfU7h70ADhqmv6epBStuOAY2eBKYN+GB5M4uS4ZrJUGJYttmZLoAc+
9+IjZ1dtFl+swTGH5Ol0nNKwNjnY9tOlJU5dTRbypeXnBZWkJKZSALMZOjCybX5y
gcoOUsA5zRgB7snyLqI9DJUxomyL4kTznBX/4tYuKUhegpr1lbN193+dns+z2mfp
CTsw06pKEgJZwMbpgSttWNrWS4V8Luqg3YPoGA45V/P7uOFt6dNp2ex1JEkslUd5
qhlPFZebWTzJlV8aS1CN9596INlAjRGUdxO9x7+HwQ6JMHV3eOLHCtS2YC5KHvvV
eS3IHxdD72PexPA9NaTYgMbekwPAciiLU1MOb0Q/copykkCpAtK2EN+DlqWF3DPN
riGkwLYTkPexkdRa/kw/+P/IHdddu6wgWUWTNk0FVyICfBKekw5shkC3x0LQ0C/7
jqbWAtl4rWPufGT5t27tS6V/RA4FW2yC9jdA9VZxgpvaqqL+8/8Ubls73me0GQor
AY/jY5csoGr33vSbvMzQe9ukyg5wjlqGzOIO5CTdMBDE3Gv2NRj2BPQ7TwUjYGDs
DMBJc0GGURW25ss2jSDhvX/G2bcM6EdQeWKvhNXk+TunPyipw2TXOt8VQtqrLQcV
s+tKOyvWHTg+iLWIQyzzY/IB3RjJf7WODsUWn5aKfFKG2ZONs9C3oHRR0ltABNch
BurGoLRhyjWqteyQsZIC6ZtAXGjQB0bd/BFWWa96F8CeMivdj/KluDqWpbd+spW/
nAeH5GNoCNxyB7nQjQOswH5FUx/DYc+LqGiqQPsbnoEmoNCktG0BmOccZfc+vuZp
eYN1vkcdpyYjyeo3O94RK2o0BnBuHnr5zumgCZaRY25ADLm04d0Z51BVtuIOXM97
46TshxeSgWR2cYWhx8n/eO6MC1jMfVu7Y510yxQ9Nga1N2lSeTYddI5l+PCTE6F2
rlmPqdyhZ/A511X3Wf5nUaDcWodK/oZ1vKsK5CycOy34ZlfW6QgjQEt3DyoKy0iK
HJmv0yehz4hVleiU4ysvwdfL7BIwsVXcibPZHsEQj2HCU1dELaMutV2KYChrMwoA
jf6aLcXfFzGMj2WWQQxwL4OmwrLcQG26xCJyYmpjdLbapbyw79+oHkweN93IqOF+
RRrq24K1Cpr3TlAWQGvewBpQH+YkHkzdT92fDenbBRBZccro7rGu8tTrRFkmLxS0
OQzKb2eIiRfV7QHfua/Nb029XmYKbl+eKpOs2eFc2K9nzsJ5tpvkooUH4J7KyQaO
mxMZYo3+MMOApZTZ/Q36uy5kbY1BrtmQd+nBICTI+Efwu44uIb+sUWauzWFXHyrT
FVRT4hyD/0MEdOhj6tBNyrYPP3PuOruXfMZksk9Zd39t6GXDX1LRPcjdrCKvgIpr
+NaPgQm+gOH8WC4JbY0InoCq2jwUuCGTANEPXv/aVnwiRhTrHV2eon+cjxxP3403
0njeg7wgAP+YTbNtR3MlQKbcz3OjMaOddOl9xZwuaoutw4PaHbzH2mvXalTrfuvb
fgM6IbWIwsY6JoHb40P5mPAtDkmGOgW4AERoQtWNjYKYNgYsUOqUyd6ET/PsX0ze
6IrfNJyuPrCv+hxOqwXv5BlppCBZvz27DSRC6ndSnnV6p/UoAW9LTEgUu4gtiyFO
tuBHi23dOn5JRaGnNwMGLGKlHrnfmi30U6zBJirg/yjiZfom7Pcht/I7iwJQ6OpW
lVpGUX/IYCTVOxKMeSx67bD/VMqDoCUMJ/JuctJAVZYH7afPGMNyFwseeVELt2j2
VZpt1uOkqhuW9m8yM04NYwJVVUZEkbsJCp/J8tC666q7B4d1UVTPb0yqhre6F5M/
zvt5QmwO1MPQz5FZxc1Q/kM8s3G+GCKdGAQE2IsJFHlxYdIByfxtv6HGu6+pPGLp
b6kAg2db1Sr0/XWRE+yaW653eXxZ1UUlhBiHuZEXmyr78igOXyR4dqY00UYSmIgZ
G3rGjzS45liBE4NlAPNPeZi0js/3ntCbRal7sv1kT0dgAHqQQ/wqDnY4Cdri040B
H0gftCtJu3jecGN1ki8rCFOrK1pmPpXX2Smxqdj1dGqISqMNEbO8Q6t46D0TzzZ4
EBWHYShnrBqR2c98grzynsPxzGWZvzxtfVxg4ABgQmheLVFkUeUi3DBMyLtZYMdx
nwF2NxfNArLH+q8RXdbqlQDXYW9NnI0VahNWzloEhWA8Yh5Nm0toTEgGwqiGrOiW
iD6UMGKFHsdxaWf+tMl9e/oQms1cfqg4o/lvxZ8QkNWdKFpoTaMEgQh2Qo4NNWV3
qQXcMBKCquK6KbEcsiJjRWiCC98yIWL1+64pxDjjU34XGiGE9FKwDK86jT9cWrhx
TR2fvzzI+1uHa0IQKfmpZ/llInSSfhC1cFGKZv+AVkoGgiYn7AsvD0+BD3JSIENl
K+XTdhXqQ+Cx1dOCYJ2ICGBEJYZTAY3382WmrX+JsDqAzQgezdV8Tv20MdoN0hVC
kheUKHbMFbcpnZVF/RNIVYClCD068M/zWusM6yXIc3862HUDDYoT4OCgAN4wk2P/
CXMfrEM668xtGz+9abVolNcmIVQK80MrUhMtZALaY6DXwxXMpXFYyuyvdbKp9pQE
W4wP0mCje4UNzp9YG3pZW97dvhkXUAg2FLU8aXnes64G5534o7BEYIQOT4gvPdVp
S7DPocZaMmfnjre/APbM6VM7zWahm8PbdAr7vXJu2XAEKXsaO9ef8fguTWmoznjN
XdlvhNzKDDknEdP530zMuRIN6CEn1lFMJbFjaz6wcH0GnLX8HIq6YZew96Nl7Jho
gsc5ksioqhNXhS96YXWQIaiF3C5J0bo9YgvRzuOVa1XbpB0SRj/ZZqhlhCVg85HE
Z3NB5f4surEJtFEfaXFaCf83h72ZR6qDzX/oKHpE60c64zixfoEiVnpMPiBLt4q6
LQovDOeg6rxoo0vEHhIl+EPys04Z49ZVGvqOIpSJgsIzMpUtJcRDcDtevHc6CUSE
j0ObFvPCjNQ3657qSvyeerNyT2rKnI1OA3fnWgagOy+/MiysYjLrErqkN2A3jVq6
GQfGS3bMGc5ewYQNBI3fkZxBCvFwSbTZn5S0ZNIfzG/E1NiLcDRDCaKXWPMK46k+
2/MBMFYOqSwNJD7N1Mr/VHc7pPE+v5w3DbqAOfW6kbOQ9toXqvZhMDeRUSM5jF+J
zao/CMFdJMBnY4x+i9CXlmsoEbWPOSmiAWN9SRdQWwBVSeb6S9eR6l9Xi0XfdQK8
pa5VJBclcbnYbpFisBBJjprpkJBfxalGZyYKFEzwJGREdepgPZxBJL8YhSQTc/MK
YRl3jLpDENTJALp81j118TlptQAQEUbrP832UVF2QtYsSNjj4LmQTut2ZRWz7T1U
jlhriKqKkT0XaC+zSWQJRcOflhQpTT0knhtwnm/LZrSfFF4qFjlTT9vbiGE2t38J
rxgCwak/LNCyV2WYXfJ34uueSouC319J2xrz1O6ckSy+s/5n5puVuwegAnd9A8Uo
ueTWTlYmMd33+28hrKbCRpkbB5MtWLAPBjQSj/7wEYEICH0UhqgiAtp4cveOCKPV
0wSN+gAvhiIMxFEi0RVY18LFKbcvVL1xVt3Zb5v0CWqq7Fn/jfD+aKLMPypVlihz
TSxURWXaZO6nWOBzKQeR9TJ4PfhVU5bt794BcM5L3bCDqpJR+7qmfErkKPNmwrQx
iKhFZdqnbWAQVl3wfcnSoyKqnPoGqaepsr91RGoRgSuGgVQ7eYso+kIC8I8H7DAX
u7djEopec7zbmJSSUruMdWl7ioDKt+yBkrwVrpz2g8ebx6WVlORNqtNpv2Ld9BgK
kgf6JIJH1asJtvgSvIP/HOfzs8S6woNMdlJIXltvEggeq9bTZtVH0+GplmEQ+Sqx
54/J4lngapVq9KgeVkj+oXXSggLNBEsyC4unKVfUtZG9qIxKllKtsivx9sFxTqQO
XolYHctBvqQNKkpzZt9r/Bv3GnvSKChzS/9P4akeUxs0m1U+M+Q6pZ8Ob0rgcz6F
Yjqvd36hXIEsxeEkU316yqHYy2O86Y5JDPWso2KfCY7vAkB5ohxm8dO6WDdozf/n
Eu+MESD0XNXerhCJVQlMQMVi+XYAXGGWc6QWbGj3hlJqrluUz89OYRcpRl4V9s5V
hos3jIAXQWQ1LVDpZAvIr3p7CxlBSQ8wRiFiw07XaL6sCzp0kRgMNI7VVVfoxRfG
bh0L1hgeirTge3B77ldjx3bAL97lfyxsQLa+wsYotjAUDtjxZ9vYm5akmmq9h0QL
8ZXntXtU6WCo2oO3OPQXyiWeS6c+o9F3I93FHkLzrZGbjd5GlhzIN2NQ0a4RVIec
Q8W90rhUI+FOFYLmVbH2VJy8lQJGbZWLDEtDb3VRCRvBtBgbn1VETea8AALGKdin
lc8c68ivH4sz7atqAIT35o5fJFKQeyb1EIro2Pbjlmu0Rgm4tAZpRk6zI2ClZUm8
WmlM0Ryfb44/Rx3VlMFJXSD/uHCn0A0mw2JXb9CPKxxZa6QWI5xehHDofG+QlENb
mAq66FAXWo1d9TJgURvIsYQsoykTFswkkhh3T3Umw7yxXPmV7v8iknjwtZkGiaeJ
xa4xWtc1KgMKP9GHiphLW1990Sx5odbrCT+IR96ZbnhzhpLv2RgsYbbPI57Jxp2r
gMMqGG3t3CPDYB4dMR4PPq/1uVzQXm0rN2YNfJuz5N8SOUYjrhOVmdf8VJT1LYMg
uuj8WrsbYAC6O0iU7zelstcI2/b9AvE5gB72roRuHV0NBX6OB08FeS4xFKV/7MNX
16mqmFpxVh+VsZV8rtas/Gu4YN/KFBRsr7HbnJ3UFuY8nDdRU6KxeTzjIhpkfqqn
JsXFgeRUgt6xj4MyMx1P4A0xjEEm8b0apwMTIkeF23x9vdxn9WH6lsNQmRIg5Z/a
6nfPC9mBmhyRVQuZJkNRTTOS5ahMTX8KQKcub4dC7G5eOppn+JBON1waGotUTSp5
2UeXTs6/jiXUgNtVPML2pH/BDacJ6t+4Y4fz0BeLdlE8+FXYBw7xuW/Nlqi5/7u4
sAL4+H0Oo3tDMaeoyX7W3VQ6geJfxMWbDLzOa2OUDTm4Ilw48jPh8doJT5AGq4p/
Afx0P93o6sZi8AEVT4/FU/aWlCF7/2DqUUNDRy0czbujz8uC78EUnJTKOPgIx3i3
/+1Bg/a0MUjOWJZVAy41kxbpGOhFrFlo3VeaMAuVeYlXaWOexWvHYF5JOQFiUGBw
SwJ62XsyFGGyMndfDozQkkIWo6VbBmyak9KR6PR1ZhC5xovkO1GNM3LoCbHW83tu
HeAfZBHhJtY9Ikchjde6D5tMhYhzDpp/OkXNFnZ4GKO+ZQG8J/Dibt63SWMDvhUn
JQyfby+i+tNVM5kGqKVsg6rTWKU9xsdSoE+4Dh7SGaLdOYdx6/oaPH6c+02kTNxt
ZdVbdNfsqUHLBkOe3htLljcHlBsnwGU+JtjM4nieIawTZ4KMtFRphPmdq0ZMbI04
gsqPX2oeq/Hc6tDSKamE1VAOeQ5Ng4OHdbmV6jWvJZW4pkcLeIXYZ+hAlE0odW7v
myuV5FfRoMSSxtVyZJDL6YlcfEYgDB6lTmTtkvTm8U0sqzKY6b1rmkxsGtZFf9N+
r2xGLUUVaFhZQI/p+0ryh8S0c+VAna697h7A8+fCLvfZmYuLjgYrduL09E7gAMkb
BHtwVDagx11Wil6bXFViaHqTr+H1OIW8RW0m8kO8gYeoK3FBlc4JM9OVN/tB4pqe
wlUElznCPqwLGTj7f+hS2PQnOtHeEJ4bhbHeTdPVRCdc9GBVEbXSAf5TTes8NRw2
QnZtEPECi0NTXb5JFBIgw4kkxnJQz2qGlaKNsRmVAmYaOWXJLyy4sBvvl6n42q1Q
xbqX5UgQ68THHSE2ns5uJ9hUUrkJKUG3Eel8DBk1hi8Y66Agq7S67v+xJDAIQkNA
440xwFYPnzgSe+qs1hX8onKfieVU+CMEFeEjxCWgPRYTK8jWvRB7nGBvtb2kdJBg
SCurpLAnR3c71BGnryyhsmzMXsCbTJorEN8YT5pgubYrH7iUdU3Vp9fA4mADSXDU
BxhALfOhtgJKiFqLjkHelW0z6Sel9LPJC4j+9J990rYj22FVKbdUG5l3MJh0FD5b
Qx/nRcyPM0xmP/p5vn7pqVm9V7bVHdsAfKaFquI3xqYD1wV8hJuq9RBzTc3Hj3ad
SBdFimOv+34/4O7j7Kr35ZfY2aQ+FbI6f1GnGJaJaksq4+AU88JVJjqfQuZMXTLt
Q75Dm/ZRirAEyV2EkTjE88m5310GdBNPWAF1qrCIME+R5aW3cFhN7s6/xeJIcfau
EoGKpuftYT6TLykZ5r4zZ/2WqHUCgS/xLPV5nhHM1TIJwGIR7tAwglaQ57IVIlRR
I1Drthe2PmCNWF5ZigkIzOStytsq83OGK3b3sRGRbnOp5w/kKMl7CxzPjTfuSPmn
1u9PyCe5HjEzBZCPhfs2No7+QoQ/qsmr+pLrQxXqqxUPEx/XyVJ497jhuKojgbko
DucCrxRj6k3XzVsRRiiVX++CKnt36qwvEZ6iOWmwHJwIVVkjAvtOE0ePaF6+RX7q
oZ6DxtZaxj+njMkIK40v3F/B8mezbyIBzvHqag8WPo3Y7dxSsqKcXFh6qTb+XPWu
YmxO4mUJQSXm68aHG2IzNzKbcR2uKdIbrv2Mz2v3vc0705IwpxDNbah0oozqLwUb
5muac5cYe8zRZeknfLTgpxaUdbi1zD6k3gYFgv0XgOLKla3gccOkR/PNNT5TLxdb
wMyQxdAXrK7qbBlrLxYzXcWZUJbqVBMaRwZx2/WTXNtPv34m6EwCAQWwqXA5uF83
6bQSzoX3HzKp5AndqrtoDleCNroXIwP/UiLG9nGEHtngNMDbJ6Q8MfnzueGmiO/Q
mOANa4LYPVx8wiH0vj+PYinuExQJKZ+m9+PIh0OqVYkEDPUZH45rdbx8lTdBCBih
hMbGDmT85V3ZqkAde4NqY8baYnyIssUxVe1YaoMg1obFYbn9357aVpXF1+PftrwQ
363uh3EPApvMYzHZgxGqIwGuuSz5+83ulnq6eWY8/FbMGMAC753viKrAWnAMJtLT
PkQIGPv6oEwIZwMCT478mJhBy96FRe8dP4sD3WkuDBo6bZ+GImh4oXh7Q5On0xdH
aeeaT3LnxL4pMrcVH0/95bPvz9XwEPG/HQ+wissr7c5ZjJ0MwXIlruR/E46jObpA
61XvufMpabIuH8O7W3ejBOR5vWu32ZZ2NpFslW9vxKbUhSVUg4fQmQgzS0X28HBU
sHFtMbt5/DeepzqvZT937k3iLwVBFDUN4yLf03Wged3vIKv+Xijh3ls75QSeWod5
vq8/YEc1LSLxFriy8VI2TOgMTaxve9IpgZv+AJTbaahIBvp/iPASl/yMxpTsRAEY
DNZAWsNJYfWKls/s0TNTjSRi4zdsNRBdFwUPnU6xEsBwtw1Q+BsKgzMzK3d44dla
jpob7BE+9TvUeKZfEB0VUxs0+PdvNlP5En4ifmqNgK07ssXBxjSl/4Ut+I7WMH+H
/vuJPeK30jQa3b8q8blGAjIvvoSBzwwKf1LHbEa23SsMGR+EGvK0q5VGA5LkmYsj
L6I4jmL/+VKWjV15Ct++CWHZwj+Fx8M6HpyoOmxODqDyAGJqURqrkYTxzJLkw3Et
eYq20aqdTbWZOIWtVG4oGiL/azwy5oJ2jLGNT0P1Aemtm5d6Dy3TEliSsReVpWI+
g2sFkxumQDnMAF9qpMiwzV5juM/ZPliXVKEFESUMumLy/Q8b5nx5ahCUp84pn/GK
wgjv4XK0urD59/9Zc7unB4Mrto2z1q7INRTTg+QlDvr0EHciR0KtoXNOrGUAztN6
PAhZb8I0hceSGMrDtNM7L3gcz2SsVDXCDRsgMZCIgq7Vy47aP7f+kBP5xTvy2Aca
gooAiKHgSypk5EVrnllnd2CTWIcBkswF4QT80IOa5AXTuPkjNnODPH1kpCXLCJho
n+OXBK+FAZjyonVtE7prd0/Xl05tGTSez4+SC+o2/7eK6nm4q05K5h/84B4A24Dv
hif4AAhyA4kZ8tH1/cLGaD30hP7RybYMmO2UBi/+nTraxS4bESNQccqhoxoir61C
hhbqpSXWPYmrYUEPtP8OJyrRB2C0NYW04aR0BU2vf+8U7uDXBE8qyXkrAJw9hSlv
S1F+hqcvG79cUhAPpyIWfLzhnEf+j+lgE7NwC3pUulsAXNYlFS6Cqps9cJmzQZ/D
snjb632Fh55wfm/dblYtYeHe9crtylA+EddZB8lq/x3+sb3R+Ew5PgEcF5ovV241
Q50R12wMVPuDMpIaKP8IsKCBBXY5T5VnJHcmNZhArDcq0gU4OUrdOCBttjR7jX1L
SZOur1eP11/SeUKfouC0j8HLu+DP30qDq7TnToibrML4sIbG++HKN01YAXHEW9b5
ZbPjHnz1IjC0605Q14wRgZ4uz/EM/yXRyk8yfmqmP269thR4dLQIEgh26RBjttpu
mlBHZU8SMd/WuCccpyE4R6NEf0Oiw+wzM8SkPpmvADe4vJQKgumqf/fdgPJKA7i3
M1RgCQmeMR34SxQwxPjdsfV+5cBsyV1Ja3j5Fv/18ZYcc30LbzWcdoIrAV5pZwgM
kpyctG95Zz1uN5T63sjH+Gwyb1zC8693zSloPUuzf76rQ7QLICHgazhrB455kTA2
6bB/0mNMslQbSUaiquKd1sBAqaSwEsP7wKphW108KjBvvrSAoZ//m7z30pW/C0Wk
/5AW4gHt14uXAwb4f/3ENCHkDG1mMSruKikYlX04oBkFofJt789JqopGGyDVG9w/
pc9/ambiziqECb6THTy0FmYLlBMveWwS532zL74/Dm3HUDVZwnmLdXYO3Kc45ZGs
AXl1yhSXsZ99sv1ZFH0Nv9j+2wAifgULLrRQBg9ous2tR/aOwTWiyiMzUw7YEuso
r4P9qlWHygCPH5qpaDvclBsg5zV0s2kEUjRFm3Km7XWceLrV+epQYamfPcMm0vMD
VY+PwG0E4sOxj3I4qzKfMJb39u1s5S5X3W7wOpBv6SqwPABylEIs2ODDN8kYZT6h
GK7FOFQZHDjRocE0lTboWf/pXb+4qnW3/zRib5FfWba9C9mz25Z61t+h7QaKsmz3
apHkhiHwaoQA3pocTkMYm0H794NhoTFViKGCubgZN7zXVuROPAHs87qAXSSHxT3z
U9fltZefYPTvdBedS0yIJ/6j+v9zJHE85SnziDy3MKIAeIML+jGsdkcmclZdlo1k
zhr+n74Nmk+2lXBRGlAzzl9s5wBbXIcWfRPo/ZDhTQcfDqMq7A4QC7EgiHrBf2Ac
1hIfu3QK/21328LiJBqnc4fjGh+o+KQUVvyQjcyB0iTQ52Hk1UpX8/EqAs37X8bs
iK9sT6apKCEIfjI9Qdkk1byI1rDFjrvNRTXL8q8OU4XWWGy/wgXm24zKAaM0wU55
e+yEL3DyipL1RYJof+mfTnWuLYOTbiH0flP97AUkW+hqySYVC3LprN4FFI4dFCcj
OB+DyH8MbSFqCVX5E0I0oKq5ISOOPX0VJs3UOcRwKoUQ06ePLbPkqyDfaUkGV1EG
YNCJX6g1XQ8A17+RK/fr/dPEOwBEX7qyXhpz3/t8Q3VEwNrEsKhE4EdhQ+JYOl+T
GNubY4CM1G+VwznNDFg9ePW/LIcjpq3i3tzeIrWlDa3nPvLAfvhI+omcdFdyzPDa
dvuRUcJm7vlKFvBYp4IU8cIfOv84XlOlLzkFFOYoZ8aOXuQhfcmCETGIWkKRyN6w
OboUZWY6UpIyuqWkeiGiekbgUYZUk9lAUfc01LHLxmNxCjyiUQk2DdcpIf13Nz0M
QnydP5CN9iEesOH1IAHCk1MIb5TCH2SQgBl/OKfnAcOZgAE51QqmE7dnNttfiQmm
fhjz22sbJx5IuVudpUOyDdgFykln6Xf29YnMLm/0g1upZ0jAu+xPV16olrSmAfjD
DqF5WT7PodbgTrwQ7adbxGNZkd+cjVEmuSkz0mXbFJqaO+F5VjRLIq1UZsz5nUoK
g1p3TNaxyzGNsgiWsWqBPf7r7KCWZIhvTrsjzGmDN4XxbkCpHwY43mUEXKHgNOkI
FpZw3gB0DdXPDZ0v6GNkMGZuv7Wy3520dc/RQ/oV/wfHupKASQUXOrtipE1T3ns8
NLOl+E3M0RmJx6U+xE6sbPnmE9bKhdumALZ7P2Tnl85pcfZzxHQ8OTtFYbn3q5B1
r8m9FymDrJlztZ06kIOIK1Lro7lEacs/Ofkfy+utvBh+mbkbUubTftd8QqinanuO
Q1yI6fkD3+OrI2JEk85AROoZM8fNomNb2d0eoHFl6euoaB77vpjmm32/BPUcCGsZ
g0pg7mRLKAfJqqtzbhMENVfT465WfMjgRdLkAfWfXO+nDvLZtokrrx29/n02nySO
MpuTZL3cOOgdLTMKZW3u9KWxtETSQDlyRALgwNj4uB2ceh8oJcvpKFgXPta0dfAX
MuEcKTMmiQc2jhY/dKfiedK63c7bmOqdUheFvZJ/ht4qOo+W7W7Yyb+WqEWIzicR
iqgAXHqhC/wCImHiqr1CSVnq4PO3S5xKrCKwJL+Y1iJyHhH1AKV3VCfiPJUFkMGn
O7xAdRqRHkL/pFOu2zA8NRt1CDOcs5sOUdyXchT19wUCUxj55BgHkwZkIvVQJN/X
H43DEITM2NdcVb2wnV8o+j03CT/bshWUwWqjLqCHzp/9Oz+FXn3Kpd7alGjkcWJ2
vIcZ5C/ExY0I27AhV+ud1Qmfum1ZNXkflU0IgwEvmNQqqmC3DvJ+2c1/dByZqwwQ
ovWTMAk2HPHSaqFfdiIwmfQtQeT5tHYCvtFRxNinflClVBZit5lucCcsMRj2bp30
xpPfHx3gATMmrQ5RgO6QV2W4M/xnyv4mOq6TVb7PQaE5mcs/eIlcfK9jqFdV+re9
RnkAkFNsHNenLkAQXyLg/Wj/4rFmcuqHS+G+hty54G5kEadjZY16ZhKLNgUmLwU5
cn9KyLIQ1c19a34zcIIdCD1LLLkW/K/SUR4NUh/QYoOtueiffiIuIhwKvD0L3viE
eQmRi6KyDiHehF4ZAl8qfkvYEspy3wPUZNN3ooMZzr93PE8ff+mdWb/zQ+X7IhtL
V4CtsbPOmqYuUtb9MZggylNb29Y0aEnQlr5EiX/f9jgaj/kUH+BLY56jw3vFkMs/
DL5mostg2W3P11QeUe0k1b7GSrpjXdhqX96xr1cqj92+6AueiNEJo+kdpJzYj+TM
hXGvfl1+AKcvmaPESHHjUj0cGYB339OrvUAFwK/nzl37CsQzJY7KyGAsnDouyNJw
ESRm2H81pBeQM8Z3bVio6HDmuaiNMO0CmhwDEoIqvzV5+LeqKeZzS/B0ZxxCKA4t
cR9Y7pYbb3n3Ug7r3xoXUGzVqfkJuswmmDcgnL/j2Inwt3Wj8FEAgcD+TMFDHRdO
/E6Gpn3ozH387Rq5tpac0ByJgwZqEAOfqc2rpLfNaTNzixjlYyhguXzkV9Z5oCFx
8DnwneAU4ysMd6MX9DgBR+aD2PzX9FCRKE0CupyeWSE5TM2n27lZX7FYwUZOxoKO
Z9vxgn4MQscxn1cP0kjN07BL/M35dA1m7gc59bVi0F/yaiJy1LEw9XObmhFLsKfk
7QwG9cR1N5218lCnrzmweGqGoxHte48xnGpC30CRtbGLWvCtbhUZNqTmFpXsVuVT
PEAZic3pZrD9VHUXOSJfWwixUWVPBa4Xps60I/FKi0maWAiUuUwnhwZqtR9f03zl
YhVkKwZtRF6Y2ja4zKRiroErXulNGNO5kJOtunWScWnRsx9+sAFGpKdW6EruWggU
x3oBnVmXJz4b2l3Xas46c9SO6WBIZslDQLYEFAYPksqY3Tx0ZtvRj4byOtOA7fR3
f9zfX8KvjP6+rT+ZSsd0ZEV9AroO44hM9awFhDsuzeSHQEGDORZVOALjWgU7GMH/
3ZRZt1/sVzywb1DGWpVe/dBaN4KWtbI0ptSdnukUXVshE3irmLE/3EuJTNKUnIe5
abIeAOJx0DAvNfQ4+45bHxgw+0eb2RCrbdTu6gZHBB8MRRh3+zUz6Dxum++gX6Um
0FMJzWS1/hgTCuMjF5nxLQOh9MAiZpe3r2AI7N++NBX9sicMTnql8CtF2Bsb4VOx
HbHx0gZDaJs6IxqsPpL9dvMq3dOaRXhxmoG5XvjiAsuu/gb+slSW9d7OmviwlZCT
8PDcL6XtkY9zGr2P/M8/H9yjQorvNRUZRDRh1v4xULJ13sCI8Q7AOVBEKebk9eMt
wudpomv1+nRan1oO6h6xLAeva01Fz7pIch4gD3IZaRyK6UhA1qY2n9CRkc2v3v/s
52q0ySCE2TqW9nxCAgStWl67RqBF+dGTH85vQJON/jop2D4mNljSjVwCGQ5DIcif
tFfvy/Nyk9Fwgopf58Jdj+4leii2GHoM4MB70o0uDrX0T4tKYUVBNHGWCOml63Lh
msxLA+cil1wKoQEaFbqa15mgyMFNcpLnZFzKOU8knsowVPF/b+XpfPAWvaz0Opcn
xQCdOFfgbYqZ0yQ1BI8BR9ycQ00GO48xCyhy8BycFG1dFUR78tmmdobEERycVkr+
boDfL9cGzXGZM+qzUI6pN3sj0In7zyKJFn0jhLr/C8Y0pZQgOlpz1n0IFQ79ZRJc
p5+wZX39TqeWbuYwIDnVjwXkpTSFOqCOOV7Qu5aSwTMZ4ces0M+Zc3vGsXFPVKfd
RTVEyBYJc0SwWGaiDl+zB8BsuIaWr6OMOEixgaHH61v6ubLuhi+hnJzUHoVad/Cx
smb61waRM5KzXe3HsUeh9XTKJfWydN605BysaU7fuB29fy5gnBoal2vOQ/2gj7kP
wbZA4f6wO+PpwXg5gvnQu7SKDT/KNu+mKcSiVIebDXIxSfITANa6YmymUgaWk9LU
mFPvZnCguznZNet+niIQQV16pu+yX0p98cm7/ePWAgMVRum4O7XjQKM79qQP2oOh
+cv423CAoHA5E4YpoCnLL/Tc2kfBbi3hWpyp0yz8izb56LTo4z38gUv0W8+ELnE/
M+XMNzM5Jq6Jza1MLfklCIZvYcK8XIOn/Wuaa0+1TSUdtXYaRYdbe7HVf0MmAqwx
cQQzXpdck0AQ0kfDSv90WsHTXH3x9EwuDYsNEMjXBel50aAM+Vv1xWSLX0q62GQb
/SpxVxLzvFuf8wMXkKVfnNMPpbgfQcbs7lDWddqmhDpOkxW60NtueCuLDloPhuDF
G+FP2+tecMBNpUEWsRErrh9jK2QJ00mnDQlXRfR71KS8ZFc2bT84bjSJ/4UrpsTr
BIluxm9t0HEoGRhqPqozRgtGfyMz9XCeVnmHKzhuGsz2Qno6tXoJ2nhUAZvAO66J
koG8UKIANFTl/7bnVX2LglUosS6s/jPaWi9RUlz+Qzd3QRS3dnt0a+eVRcNozlaC
9btW2JWtE3iSHhs6o87gl0UFWD0tJlOF+6X8AayGHjVnCoU5Z11unLlVoK4SnDrR
tGIrxU3GHFvFlgdnoF9XyB/rAB5MFZ1/tr/cPN7/yEs1HoLwbQqhlI3PK7XfL8RG
ARIICWFCGTT55HHQzqDuFApjqsNDqqU9rLlX2gAOI2s8lHNsP0dinDptLDAMku+E
CKpT61ziWZL2dJna9RH54AvNYfI5xDrLIOBTViFP79twGfFz5eLYLGJ2HJJ0Q5e8
CWSkP1oLA0UkdPyvsB4Og8E410utJ+g3MWeKUh+n1A6y6AUaxPCrs8C/KI12mAJw
yxCN89AwayLkmlNlPTSbMc/bvQMiv4XxQDsHE6s4sml7MO0wq+El+saOhcSZiZeC
HG8uCjYd++y3nPB1/9iN3k/T23FCUurgd2UXlud7Xqsn3GJe+JMpT4K+QSQbC6+q
DDOFH6PFf2NUtj2hGBmuzOi1t9pvbpQUpbN3N19HZcefbBhe6idqBz1tJrQK/zjI
LqGbio4KXKpvFMIEDDpAIRPcAakBdbnrBR2mrvkdLQkYlc4QsegunskfuMLKL1Ad
hkcbx2vJhs12V61JBalSqfd3nN/HySe0AulcFiTR7zyM5yPToUXzxsD00olEauNJ
A8ctvGErF4Wr3SikDxVwrLkj2UrUvDsMGsdD63p2WrESfF/7rKrjnW/LQZodEbYH
dYbCv80MBBA920PqC9auxGupamoIVhvR/WQM65TZm4TebDj9HrfnpDLGCFQ1qwP1
SAL17SrdEZLjQ5pY4EsMYvgsKvPt8T7w16bLyuZnsKK7LFTP8ChumedN2k67gh0C
tjkStlohSW2XZsAGTGbf7dzvQVh2yUQ8KjYJIPkFuNNeeMq/j6XrSxc1XKO90HoJ
PngtO9TzMwZR0yIXy3ZwYv01DAjPHaXSj0oouwPVvGvf6eC8UMGQE09ygwjlMh37
fVuB4GPJMabliWJidlrc20L/2pFVzNVZ/sLbAqGA7/qXi9IvBm7uaPtNyWynf5zw
sYQoZMRxRVdm3+JhsQMqgLwFigC7bSzphGJkaO9M9VKyMhFKBnbhosIP/XIuOK/2
0TLN1jP4UJO0u9ADTP7tDZmhfGYVP8efT7nRpDZ03m40PxFzQNDWeLGKxACd+qUc
apcCn7AXKZ5rMOnegOymBm1BmyJNj/vv9tqwN2eHpcxlz//V1IHKqBsXBlj4r/bM
5/nA6+fMGOA7iD8YoQkQrmRgB1mSQgLnXyKvnF4F9oDND/cGxncRVHIt/98G/q0o
M8+G2GoTVhLxKqr31kUfatswHOjlJhfDaDDeYySCbTxnO4KrYOEdH2tbkm1MKLO5
zmekLDZcI6GfrdlDkpk/qKRYoocQHCtIIIMMgaz/mW0//1rV/CobdpThqZLKaKZv
HGVn5OvzHQXFJotER2xkF2tnwnZUYAb1LMxAQ1nJy8dVuU2PCpmkVYZdTZmilsGw
ukaYthnJ9dNkgAL7MWrgUAZHbJQoJGLJEgdxcGqbY38Q+/vF1Btajpcy0wIRwJ9v
`protect end_protected