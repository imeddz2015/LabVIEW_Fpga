`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 5216 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/9huKRhRMtvnNqb3Z+UU7TahEoHV+T8U3P3ufru7l1O
3DlgtZzb9QxCbOjthp9+wDkjygH0eUfDrEl1ovhZG60wIGftgTfryTG27sjHqFpC
YKKtOuffz/ng6PLvqRkiPfp5zNz+YPeBz9C1G8QfBA90Y74kggHRYrl00UIG9td3
ynUhEWx5VVWNsXezrRFOLVc+m146lQ0GX1IwZnMyYm7pPPv6NtZHNKh1hUxQcTd+
8qgxqS34ZtXqpSjVTzxPS9XpL6R3llKHAipL7lDYG14LNUacbZrjjXax8n2/EfM1
FMhER7BR/dZUTQhydxt5QmEIfykGLCFZhCau0WD3Ky+2t+isnFUB4MsrQN0ocFLZ
eHe6Uo+w9rWEagi+NtQcXncEn2Ey5i7HdyEX704CYcpKitjXFYYyGm/PRC4zPHGl
Iiyv8j5vvinREcPcnywbncudecE5NHjZjkU5xxupNzNtFJ+rWJl+U5NbOD/N/GMc
bN9bevZxSW7OQtH0qsGbNuARlItYREwwGjQOVEeIpzVDk3OQJtt3zh24fnTLBgm5
LWkoSuy9n3/573kRRddj4B6y30k3jLhR86b/7LI0S2eKApx/9NQr2ktj3omPFgGp
C24Px0fze9y0k13pkeDWk+XQ82MZmEAQPnXz4ZS1Yx12Q+MYIZvGrfuEDLllNi+J
rK3+joH8c9GdUfo/XLtqSmsqNQO1nWf3EguJSf6sNkZMHe9C7Z1l1uSE0HhP8Xlh
3toZwklQpxxctPYxktLaK7jxNBZHljeSGZ1Lxf3FEYL+p8XELJTzm3NpWNCVs3pO
zOtecD+KVxlkMiKApzkUV9uYU6Cwn0ydONSxHK6+wo7mVrykJLKJ7YScb4zRpT8S
LsLMmjnDV5kjSESyQwlNT20FbX5yz/tPQVt3l3ptNFp+7rxjzFMVW91NNzQPBWQI
tKoVBT6FtZIXvGN0RBKHfyRqHbIjiqqkq2FX8L2Ch5Kxn1G8A0XaMYQ7sFD0NEky
pfBqHECbc84XoG0lHcj8kh5jTGVfO9oNP6hnruddV9V1bQpzhOX6Fm2ZV3/K9dSi
YDF5pJrPLFVevMUdaoeNZ8lvKTdPKherYjtjjKh5aeZvtVwwKlKzknvjKEoZ88+J
LwN8rbLIqsO0H18ZTtu9FTnM+cX41bMM5yBG9UceATzd9Mw4hxC0+Jm2Zi3Wxqvc
XalK9z165r+8OfmGscCqM7Ocd1catlrLzF4Wq84fdfRR7nW5N8j9HJ6cockDXshk
yRS8QsiK7XeHHtZvVkJGdT6xykTOGrcP5w6YM4hQsianjubnq9eMWq7NI6Mp3l7t
NL1pyxAvHTN4PBbzx26Q0PigKx6spe9zPAF1Kn9s+D4bOrlGuxNhtsfchMsc6mhJ
vnasC95Jeg+YOo8Phgqjk/LcLqu746NvGgzQLah8hthmdwccw6+Z+UsJ1y+5mHDO
TQGNtZ/oAvIMIy5tXcBJXWO31SE0aMmZ4kYvt59W1n0axwyboT6wFgzrKc1NDAfu
hUSUle+ZWtH1Ff3PA5pKxsu/PId33n3KUJgAYi5kY8/KpD+WAoBdf3ODoCr7OvWJ
hFXuDVHa2v3yahAo5FZo9nukDRUvP2orqQ2JC83krIKp6kao93DC3cgM3YNTrOmD
+VGZqeu6nX+FLWXcGGsYgmAr3uAfkQn8OrgRHYiJ8I1pA8I6tTgEBuhMWe03x1rb
KjOkwxmWOcCnXdJ3h0eTjgdaL8UxrMlEY7dYHJH2KChO4f42yP8dQyJDuSnrWne0
gB6eV323yQCJSiQZzcB8X0yNKp1d2cXK2GiFjF5jFDW3MASvZahl6OBYKkUSWR+K
Fh9/zY7sHnsywtEX519WC2bv6DZEjmeiltNDX7ulvW8UPh1WGQysfK/8RwiSSDof
Y1SVttklAKRwwqNo4ZA+GF/r6IW6kNRGNVmI1ue2II0cWmmNukYECC4rdiD6d7Hc
vz5qZCt+BljaRLmeFqYlZDRBS1T3UQ1qSOVOAW02fUctO5toYLSNgvOaHboL2Sbg
rshopOQzn4cGhALLYrZ91p6ATQY4xomYkzFTRuInOeXO6K1SLB7j1chxTRzzKlZv
8NCGNnq3AXNq2WxnuHiBy4iFjL5Z1AEhhlCMHQRzEsAytMRSFbV04izSlq0cMuFF
5vut3cnCrJL4iY5CjIOqqTQ4PmPE4AvJZ3n2U0fGaOyNbjyQqo9i0ZlrR8gcfvHs
TytES+qeDgbt7VnD76HZqEx7iuhxla33Qt0mLBJ7sIy571CGuMOuOKIUq+8WRAws
0N2P/pLY9xT2ol7hlgWhQhlZ0k5655juxs1aFK56wokEjQXOLBz1e21xLoxBFq12
DDayvhToB2HGQeTPvAS8KxQr+VxilxWr6T+6xkm77k+29il9o1MHrkg1dCkiLP8W
5cKR6zAPHZieFbhXS5M7krX9jj+jY6rUyTo5KVUWGqh3XnQc23necAcO1y2vyNtC
Ydc1yUYbHe7HVNHjT1Ppf7Bpf4Jr7NAhnxTSQqAl+vuEIamf3Djw22+cU46NCfID
75yWXoBeEAMOf/20tCcB0ecwJVA1JM5HF0/fng/PsRdBSejOqtSkalMY5MbAh+vq
CseGxuIxRrCLyhFsnzaaCJlk4UPQApgoYVOGWbAigqK5ZBcKXVa3lJmhMqL8iFM5
TIPvdZqLZxmbuBZsssbJZ214R5J8IN9co0Y/T5LsKzDZ0Y6cC/J2yNH9MhmrFP0r
6FVNJiSFcg9yWFEgBLu0LLKKI9j51n44uHbRAW0Tb+VjwOYsZkS5j8XuDEKsp9LY
R/UqePVas+RBJYVYisgF5noN/YadevmTalEOquSPsOZSVaUQczt0GNKDMcnM+U09
4N1DHALde/4eKFsEPvNjHURbGOwWRajEZLsiIUE+Ks2aRO2CA3nDCRNkBIq7L2lV
Y9Qw87qu25XahV/580LZBVYV2lZSJWR6kcYh+JbRMvL4Xd6o8YbWcPyobOBB5DUc
evKT9Z8Eup3ngneCV3QVHW7AtYcQDLKv0uxM+SeKCv6fs7MVE0JvytZf21eDV+7v
dgbllZrBKaBzstHQiKcNKaxj3j3b8a4U+BsuObVXKSIo1BQcbaJ57dZnkIuskKgS
YZKTdn+FY4YbjI3vOSnMKERjpEoytwuvsOVWGV+GIL78/EZnr0l3gJEWySNe71H4
TlukGUx5cyu+Fvkv43D0EotEhZfCH4JHGleQV8L7xsuORyz3kAPxZlcZlErGdmWd
DNb001RnrfeJAKjD9tzD07Uk7SKdteIB+REyGizpkH0JcvdOEyXVNyAXqDqkUTGn
JO0N5bLqIDP+GfX7NOS699ecaXdXm2NMdoaFL/iUrK4srUYttAfDowXM7RxwKroO
8BHotmRhZMJBEqPtJiJbhG6gDdKZSpS/0UxPOa8uI4vC9w3oBpG+swtMHvRZtSuO
Uakr5W6GgIQcblLLei203690MGZSe2jgnEQ6dL2P/+nMrbdcMhWOW71jztu1XJXe
gjkoNck60abt51gfN6oKfjTv2BHWBbxCmH0++J3whppGwInemro7GQv32SOJ/4vg
Nw1SZSCa0dxS67B1TqPskDzDzbu9q7ld9cXE3sU11AeTf5jxJVVd05Kbeovx+GHU
UhjLDsEXObaaR71GV/AXKc94mml3/QDXMrj91XLmBg6pooRXX0zHN19i8xD6EQGX
s9aYOowp8TvrXoJYUAECg7sVw3S+seyBh7X0MFyS0khHncPHZMUL8Z8+K6dOY0/1
95mw0soddf1EaqcvpFB/Vvcobs8q7BEwyQFZKy6mS755M8yQ4M7CYNL9NXU03Cxk
gUCgARgnFECsrf9Oh1PidrxPhW7fPmYRSL1YgBk0XyP8/hBFO+7zPIs22oIWlTr/
Bm9cu33EjIKeR4AzEjDdbVX7AOS2IIxETBEy8NjSuA4EQgKPo9WlVz6d22Ejfbfv
+zyidLkGCwqmpnXRgKie2yo+5UvdQgjr5MYnT5XrxHJriZ972l09ZxQu6BiOrdDc
QnIrM9XTxr0h4qFakCiiSrrhG/+gdFA6HxW3SNFnk4Fx8oU5mDkExYgu9fM2rD8k
17Woa+xqodSFP2DOhltSh74z/C2ETT7MlfGSuIjzZOsKMrNBz1hvJ5r1Yl4zKj2Z
bijfOReeLPKdNRMPssqIAxyUmHbEjCUd+mD7u/d3nYKLSmoUMmpffSGJMZPRFo09
DXITIOTAOZq5IQKqWJ1A2EvU4TlpDSBIkxoq/3vVX4QeXIXXnDuDq+mIJbILCnYO
mdymE9VYULNEs916rP77TF55Jz5gN9p4XVZBizK7Y/WAN75HhzitpTv8+KeUadm2
VZksFXkdNwi2+IAYX1oRd/gcVdebJm0zYb3UcYnNt3DY9imkN7P3fp6AKojxdisn
tM2CY/eiJz2J/j+yM/447RHjTZUeMPCnXonJVY6vBDNnV8TwwVYpJ02ubZPYNu/a
IV97ddweObiUGUrlufaIQv6pi15KXeP5IWao9vVHNiSKlbNtNIItzHL2XVD2ozBX
A3i4nHfNDo/ODi9F5NNvLl3xQVcrwajpFAM0nGz6swQBOhOVVdHvi4S3QG1bReaY
IiyFzGRFDQx2kuHbR1cuZlnROp40fgU5pznH4tui2UuIXDIv0YrxJBCpv7XHf1hG
GynN0NIgly+ckDm/f8BlgmOOdUTBqLIRt1p0en9bUoM8J3S/oML9yGtRjO5VY8qq
llStAHjzMZMF1uC8XWVuDNKNPTNRePm7rAICI8dgpbjd5cT2JHQ4HcVEO4qZLr4A
u5JTxBAQ0fsx/U5bKIMimojBRpInjczeSR+xAaZ5Y0WFfa9xvkh7xibnfFjCvtMV
oKhGIooWucMEQoMJizaIktSRnbIVw+ao4ytFHff3eFW/Ld5CwR6CuU53wcnS5Cu2
Nxn5ADZd/aOPqrz1pDdWt/A4yDvcYLCYF7tVY8Ardys1ntSu32jFuFPcwalbju0c
AZQ+bLu/mdwEtD/o2sd6BRlAx4kJaBsHaDISObseT7mBQczw4x8ATPmbbTfMRUx9
aRXDbfoXUD1P1mYj8VQRMzoQx7KovSncyrsK7pNv/PmdcD9fNSukoI42x1Wp6TIn
kYptoDPAgslBhQsaFPpfkp3e29F9DKQ6KFlJ460HlRUeJMQTCaNMLdI+wihpaMnD
zpmS5q1tZgq6sg6yC0j189UTL8cvKef8Ze2ZsUMxQf0fRCYZbVcypfAHzg8z1crJ
0JWQQT/1Qygas8aAOwk/SqGymxfDmUU6sYkdx3bulXJnWQK+0tovskZs4TPq9Hk6
x1Qct4xvUTmFADug6zTSjapYMcIDHe0y7TsI4krZeRBxpWkp7NpPTPGFSrWcEMSg
Oz8F1LR3PcCJXLfFRvYMcqxWYs4Ds0srrKz32t6wpoYij0w1/uT2KDs/ZkWC7jOY
wW6yicXHQ4+8B7DF84yHFGaVnaTfDRnCqdOAgeb/kHhIGtcGkRTacG/djm3/Ja8K
xuQZx7c/z7ze1bxKvxn1yXMIT4vcytuc5zH0xQ9c6iYeSNAKeON71YzkcSIDMXAi
0oeqEIXAmpfKuBIL7V9W429dDt/PvBeexNlhxOL3nK0JQqHMOL60BBS1rqFs/1Nx
fkLIZ/jNPczhGvadjJr003QZ6EsAXJDAhZEE8T2WxhPibpwasqU5ZwnYuqaENX9/
ivvmOBT/FM5Z4tGzNgsYpchZvVQQWcd5sdjNNX0lwKHwEP4OdzdlZmV/YGe7lO8g
K9KCUDd4wxhjTlcuMHqTSgV0puF8EZETge5nFKGZCWWC//Dvb3UOkNm3523PqWoe
cYW+3W9W0egiMoB7cxK9HgOMPWht+58H/pTUUxZ8GBUXwQ3hPD8DWybxi4Nhb6eY
CS6SQ4GDLHOVlWtPb1kJLSFvz1yxJKRY6p+ymPctozizM4VIsriLB4v6nv1NWxRX
l5we8fUu3tObNLao8xcGxsS8mahNJZeN6mDza7Y2JFSwTtIfzRv7UEWZf5rIbwO3
k1jVYfVaxYdqndlKEGOJK6YGLIGcqfbQu0i5u2aVkZfYdplH1Ae2lURmP1XzmIJU
CYnEfJWlaIkrArNS+Cgf8DqkG6ZSUDUtKVzBSN8mF6xqgWekzYDiAbi66bV+rq3h
Kn+EnApQEYBUUQJV+AN7Y6h3Lsp1eO6cAgw8g12mf0fZdJvsRmL+wZbz5MvHA7XV
+C5/1KpehGbWYEXzegUZolPt8p/iJ9rjspReHk/ZHma1rXAw9/sd/OJXi0EpzE+b
p8FTnRjySLZlOhI+95+Z5Day2b463IkZ0p3i8Fag70vk6yOWsKUfQ8sRdIAaS6i4
oRsoiiC7zEr/4BnagmhKxH+8O2Pa5zssBgtdBdwKpUYmtGadE26PlzcEppvdMP6A
QYIXHhN3WVBESvq6UC1rPpEdBk2sr2xo99ZLLRAmwwPqUe7VP/ViaYP4rbRezaO/
L9/0sSxkIZsT53GmKQ5ekhvPImUF241hakCw2V+VPCjbEjqz1cjTPuMF0ZhGyPYf
RaAOquOM+u1ujI/osEcjhZT0+qzkLw5oxK9+zjXDlE7xDgbOk2/kRg9471wIyf81
cB/Yk2iWBOZIWvDRbvcM4hUfXiJNsxsLjFg01sP0wkMkHpsfa+/Gqs6AbmBZby0D
ZFT3w9t2zjX6GSU876wtJ74BTmpJHpJp8BwWnlMZtfAIithOcNRdbCbntf9DYDRA
0srsQWpskNQTBlKdd4lNw4KCmuVAJ9AilRu08g0qifW5azAg8Vei1e3sboMEvFmN
sClhGDlccumhG+t8USg1LsaKcqxH+DF/fXNu/2F6c7qHSrBMFeDfVTvHDLdP6Tl8
7GokVqJ7NNJahl8p5oolBAiZsRNBqQPeAJClNj1r+eXEtUmtIUjrwytYHiR9XUAZ
pML/OPh3DyH9pnExvRu4EvhQOguDd0P3zI41lcKc5OQ=
`protect end_protected