`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 26640 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/59UwEX+aE7FohaWu0/8IpTj7mav863zUNIsgIH2BWb
Abd9opeuBjbGF/waQMI2vMJTwD1ie1YueHc3nSNpEh4OXp8P5ybZFY89uyGz3ztU
W1EsuUnchJoQgbHZ/sLbgtGRgsrAFn+ZoIeGN1d6RAF2wAESJmYP8zw+p00RvjZ5
G2ATm2jrAjm+J6bPpiDE311fdk8/KRYbx4wKgzx8PBiSqToDqXb+EPALsiJO/m+m
VTWcg5DeFxuMbzdVR3PgxrPvKxpK7uPPa6Ww14Huz1q8ftSVuCHIA7YaYXIUWr/H
oa/RHiIklnA8SkRJa42g5HHN8CWQ2D1xfe6Pe77vkNjamS/kSi++TXnofJiAFx49
nD2dySQ7/ulLl5HnnTLbi+MMXeafRJTvIZWMrrV8EbWYcjRUuy/ZPJx3+2TVEmRd
s1nu5+OJG+kil/92IvzRcburRfBE3Ns9f6OOPxT3+R3CKwVCt6R/rhSFysTS1kUz
Iru9otDAffF+rKfpXzXx3Gl4UI3vxPKQSTe+gdPXwKxxA5pjeNFUiWz2lDCdY1vB
DraM6fjDB/sVlbd0uxNcughUU4nr8jHPYj2pXTkI3b6hXAcQC3ZBGL3Ly1PDA2zK
FNkGNLn6ZJONY3dRBzu/mvCLt2kfZXpTj/8PS5bNDoqP7XCnIdULpkIoPyMnVt/e
zrnZiZXjV/DhI2qlpdijAQn+drwRC1h3vMra8zfWSqcTYJvCHVmg07qGKQ6YCDj8
L/v1tOlQJLobF9MUCiTNtOEV1WZCKOWZD1s05Hr2smrP21OICrxYRMPmVRcJlsxS
Zm1sC0uyfq8vqCD+LpXdoAYU3MFt5CGSfFAeRUtoU3hJu+BcJalRTsXG53c4r/+1
J8fsSIUqmzvfpby+WtXYWMF3GtAW01Y2sGPHGYBs+3atb7nDEHoRasZIAtMVlxOy
hY2fMqFd6e6hDzHyj7bHuJ86slWb18CIzlBbW+xZJpaahWGCAcvzqDlOr6Lem0Ua
Q+5+XL/AXZ1j9wHhgJzMbUgDt0deYJMJrg/W9wGVtsQClX36iYEAUOCy9GXoAyWU
EBHft7yQNxuH8qF07gKZg+KzurRKtzMVb4EQfAiGyTfwHR9+8wFy2ktPNmlYEdxB
Q/rFpSS1y35Gj8pB7tMQx7Kex1Nmq3xr3uQDEqdRBfvcje8bH+02BYX7nGFd/7Un
nudxgyM5rl3xLAbYQKaJU4SbwH+3tpuIdPNM75yVxuzGfgZ7cMnCbpPntJfv6DRv
A9qbQPrHdJA5VG7/CU+sDf5GJc6+sj5TZwVCPziqf/2uU4msw9oPjpjUHbGI0dD2
Df1NrEHxSOYNwstdzgJqVN1nNCVyHPlJaX+TbcSn5+pAKAa8UfYZVeG8VWXuyjJR
/eCDiqzFNi7D4YQhUcsZc/Ra9VpwAqv7MYUxY6b6rneeMmJf2ilA4iiEcLlSaJTP
TJtSfH8tmpAxpPAtLVv8gZhe8uUMdmWJ0ku5VSyc4M1hyI9HN9UuBU1c6bRV9t/E
jDFtdLCB+DT4RItorAFgrzZ6EQr9+GmGOtUyhZuQauFAmjtyTGQ+i+2DOESzM5iS
lNQnlOLUQeaZfUWGJZyJ/Lt7aQ8kbQv+/4EEimHsBIcHUCwuq/S6GUQtQd+Ju/h7
UI2tDtIyJRgCKh+p6nv0WA/qRRsF4qTlcqbm0hHMAGP6OAanlvB1msLLb3ZLmEAy
WUd1nYitTD4KK74UXq896r53eTraiAW9H8jsnucPI2TdmsHQs2H0QAjqe0j3QZxo
nSn78OmXBxdpeXJSNh6667jwVojuuqrJMotnaY7sCHWL1FlfanA8xNaXgJjuMYIe
5XsljzGnEK/P/ehgwMWjJ+kHf5hLkfJIBR3oruoSfLbAqIRgYF2jEJl0wphno/w9
C95/j6TWC64qIfVDVsSt3iQcbcf+MqzDbvX8IyzcGB6gpEVSHPgDKUyMe94RQmsw
/9xgi1xGL4W7Zfx9VCKeqzPmyduDN1HpQz3DDcQ7PwNlfLjGMTcyZzgNjqQFJbeg
DawrrivTnjO0CtrpUrfB79HniB+ed3LD5hF9HWyQqS5WmZN2SHzxydCK3s3Ed9yC
MN4qH5WPhQA63rutJ49smv0fNDhF1qFduzhvBCnII2nIMZI1FC8DbWM8G8ybHqnT
Sj1T1SSAn9SAJznsezJRKHDJDSubNY53YQ1L9ZdFMwieYFX57UKNdd8ehR9j6xsL
nuRjyq+3bNRSF1VQGBNhm910nUyII2wTzNPzGkDSljqJhWO3x0LISTxfn05T9bCV
PRieYnuJh/QSVjdJcrBLw+zNSQitGWvVeeSknxtNTvtNyfcb6f1J/zE++Yc0mEaM
4uaYMr0yn+KW3Y6enL3rYdJKlckW0gWEkHH5quNX82ZALB+Gb6lvKkEWR8ToQeW4
eEP+NVpfEUg9GQ01nm881xJ+gfwUokLUpoMJKoH+rp0Btv9QENDNkCOBPq+2cUuN
whQYQ9yvA4puQntm49P0HY/zvCc44qHxrPNnKeY0Nj0IR7+A+YoqXjq+glwM6R7W
Fh7dkHEDRAqvwjNNbppbVSP0jS40ZpVxqTV6rINX0Uwx074agUqnrjPwQHfcvVIM
kVMpRkE0rf7VHNN9y7cVLg9ArdOc8LmC8XlaHOA+oJOhQ1KBqnhbqD9wKmp7dbtn
s7gquZjMWpDEhgKs3oQ9eOzaR7mv26XDYlVnXojbt4rs2x2xmyAt/NrBl26lBjaN
CxNI1LiyhGp/Xjwxsp5LwwcKhKmIdB6MCT/5aVXC7QcdcQontRRh8OK1wJjlHacS
oXuV8+zFCEhcIOSOqGAXb0iJucR1x+sRLxO8kodJqiiufRg3f/qGo/aWUfKQImjw
EbLrN6TV2Ixs0x5NHM1a06I1Wb9RnS30wFIgNiZwGl3sVgGowcEjsFU5VCOJcbWp
e2SSR+f4D/In+qHLHOcKRTK4BNR+aP7CiOu508zO+OvqhtMdotV5imXPTxBV08dT
7zxU7MODQklYDl2xr7yAT2pAIF5E+XqTqjrBhmSQ12D7vnMlJEVTAI7QRXPsy7BL
J1lsLPXE+WOWBrWEBuzBnSJy+Hh0qcSY1P9AVlJYbUJigueI42DS9oaW1lkgDqzt
4pfT51hjtHf+YNA7/W1T6xSN9jHectyQ+eK/eFOYqvovl+5QOLoiEZFWF7bFsB30
zrGow1kqj32LXTyDPbl1ENJ7BMTI0JAeevrnFVocBezUq18BUL7j6dFrSGVn9ng3
ce3h849/sFaxJhiEsz9qMyIOJxfUH6TjOF3UR56jlGZSTf+dEavFfy+NVpByOKbd
XYVG00KwqeLYvB/Wo86i2S0c5UAAbdMZxDHdgtg/FOEDG59zdpUVrAkU6h1yg2Ab
bwQVB75iK/izbMghiAs2KHeoPcvaJxaNSGV3Y6bY/o3Ruj6fOCzAwGxQYGLlKT4D
4xWlpl1/lPmp1OVoQEBABtpFjsXK9JiVkWr/ZiffnfCYUvAZHMA2uz3mM77x8356
7WM410oFkSMkvsRd7PtH+hnqboaYRGaDDJ2Z4By1zeR5Ts4f9i5m1AbECp3BAKjb
AS0sR2fe8w8yYdoULa+0591g4M7nJK9GR+tmiXf4XvdC58knQlDOaeVwiAxPJGEe
izl0JQOXcCbNxQ1FiFptRFRaP9jRVybPCpYU2Pq+sTbs1wdNCGL7ronYfiZxI/dy
Ya5kH4SW7/EKgXFYmpUgIomg2nLzwxEtxt+6mYhTk46DNHRUI4/gRVczZQvQQ1BH
/TWFRbrlHrtnrF4pZMedLODhHr78DTA3H/gzpNmT5AuT07D/PaiToOuGTM2C7klC
5V0tSBYJXS4XybBB+eQG0G2q00LxPLJtl/AIP1EY3lAlak3NZtoVU/zhYRlckSFp
fAmlr7mWzCyZqq6FvRv5ZKnLoqUGtPI8h3IBxhWcuhjzQ5Oydk5vZtJkNYmrXYJB
LeOm7i4I30S5G/xifB7paMy4aXMsnERX35zF4D0IBUuTLPJYHW9yW0WYcv45Y3ws
JT6ESGJQzPSTwgTbyJ1fSSczpWqwpoys52QNvMUhP0UfSFFGKmi4IFWBOaKPJUYZ
lhz8XJc9hnRogAZ5vssECOh5lQYR+c+Wd6BW6XctV1wZN+FHaMLhyvE57jxQ8k26
NIe2ZgG3H8zyigvgADVqrtDyZ4Y8aMxlkuVEL6Vx6kJQiFmPCOZet1KrJ6mCCWoC
/SaMuKPN7hXv38VcfVUeS+rZEomd8O0xmo4nusT7Y5NToG+e4iPrNi6rypJcbK11
Yprq8LqrmNt+FBJ/R+do0IYazoKmyzSwcbEseF58UKMv7Jma5J6YSetKZV0Ybss3
aZM14U/7LNxEq9/Debuq8HjxUq5oQ5IDwlvIrXR+heXdjxEDNjGlINzqB/5Sn43z
GxBhMOi6tQetVHO8aDQIS4suDjw+nK8FJ+ptp3lGgmL35kj4DcEVsU6j4jWXWnV2
gHlkPGbxZpvr7bhu/j8DoNmbr0Upzz/LPT2sWSm4SaKziy1SxLVGMbYVlGE2JwYE
NXiY4cy29wCPDMLnoBfW7AloABhYnsC1er8YLZRd+pDfIQ15xiA7MGyFIG0yadJt
k2rE4s/IVghwJSgqjI6LDyxBZiYeE7ayzteFHMAgAhRxs7na/YXyA00hyubKuk16
/G7BmarrN5AdqsQ/O+48p1bNWGzGJhjNLN+9uoCKY4w5gQX0a4Y4pz4DnPECG99H
78m5ArSTWJ4BLZV8ohj9l176chicNxPbicUDwpkAl6klkMiThRXqEZ0rIeItxsyU
2OkWnk4up0X7rR17DQOya/baCBXtitg+OTorzdXX0sCPJE4ayw9YGeVXYPURXkVz
GQx2gqGiOmBDHb65ZxlertrQUlmzNcRTpcIiSNMA8q4TXzFX5PZyUO5jF2aq/4KG
fFFLVVyCFuN9s01e2HUCRhvpNKxTlev78VgbnCE4ZsaaRMh2yWwQYDsRXYpH3knA
HbBWyzbm5OTiYbDQa9MUsDVy3gOHe8LEPJHVsWPaXv4shA2YetRcz55/qbX86P3j
QSXX4pUxlVHXrB7tcmEPTfFmoQVkeyUFxn7tfR7VuX0DYJM8n0ZryMrJXh2Dnb3H
RlY/hSidrk8ad0QDQCmrC1uGCueBWsQokHGZM+Bax8LPIaVXDbIdhZkyAy4SKpLG
Rg7Hg0234g2Iu/g+9AWhKjkFHI90HJo6rXxhi/xgiu4J0jECj9jyYaWEUNFu5MRJ
nX45+yL/Sici5ILOUJtdH9K4jMuTblSrXEPsuZmtN4H0NpI6QS1rJtNXpAmsiRTX
AlB6nnqI4dl9n7IQt2Mt+teovZ2ngDy2n+csWhX71tnL/RnKG3D9n0QsRzKJdEVi
laTB7UsZvTmnvrDaPHWIul3Yv+gQ5ZVqBfiqtuLVdHr0z+c1QVhHXkstEQNRclQD
WxqRHBdgOIIOTlSDQ/FMlD3tPLUvNRulmn6ZTkBsX/mgS/gbfmYnSXxKzs6OjRn1
vnh2MN/iUEHAFjLs7gI3r5uXY2Vgscpoyq6zpZAigejmprsJVcm34Un4ApBnwZY3
cwHHMzLcTwzdQ/f79BhahjuxJcc5UlI2n8+Ywa2rovSBCbZ6iVWJVZ1EbkendB9C
eDcNcxyEprdZn5CFDF4u9cer9lkWFvnNKYRBRbC+sdqFKh4gmsFC3/tAJqA5f/WP
HZuGTgGEkWSgSWv2NmFmv7Y02fSEXTMA96mcOGRaWaiggcK5NHVkfglZ9wpJsfll
n7m8bEECwXVR4nXUny94BXKdDGQA6CS/wjuRjcqf9MTQG4q62w/HzAKd4tuLKCsu
EkT4T8JTX3ZJSsMv1mthJioklFCsL7580sJEb1mCffSutkQk+zzPT65XFGI6VQFz
hPZS1PjEx3vqdzmkW+MIu3kwp9ElDetD9AJ0Efu2awXpJ4Y1PC6F4uINGEZxdBxJ
nbnu46iHpJicwpKQYha6YYeaWtG/0BDlIBbqrEboEvP2ZC2n9BAD90/o9MxbzHPB
niAcFlr1BIOntdkckfD19km9dtN2t0/PwlF/KSvffjBxVOXzNxmqSwFrnihclnjn
yHT0cu1UM09zxjkSos/GYBDorJ6qRlXSjU84lbpLINiKqsDypqRUMrd8xpORcerf
T1/sPIPWU8PunNFPKyMbJ3nrO43QCilCL3fCQyJW1MSasjvyHY7ERGAKAkS4N6mA
HbYoqKyd37x9m3Qt+qMsp1L/IRtijlHoNLbN7n1/5O2cdJaHcBhHQdhSVpKmj43z
D3chGyIGRndc+pPyr36/b1EwlLlxPd2BiLlzEEQ+d1p9Vb7NfrKzaBM+3KYeDPu6
J19CXrfw1nbDydconjBuuH+J4VZHvNlhkQ/bxZlAx72nVtYANtbBBCwO9Ag6yxYz
7z0eQ2JjMuEjtgNhZzyvVCoDAJ/Z1yNJ6DSGw1Q0uoTQyb95hAwAv2u8EcmAOfmI
N9ZIMFJWCPwGGwg06VqGxfcONNOqcLzPPS702bZ5z1+11gK21VLnZuHMNM78fWWr
f9yNCepcNNYG54gQnAaJ1Vrr8CIjcZJVjH37+ExcAZMi+f23vivopNgR2ztd0sMR
gqkUTUXBCoHhYEgoRsqziqUc7eWikn5kQDT5/v3UkElTlNltxhJkrg1xkmALEE06
xO1k3q6weuTknksadxA0KWpOtpOQcplWhi3MDMa4F7WgixrX4PzEkjbAtZ1NoIz5
ERBNfahHRMOtExY1nLzQHp26+MZVlwRwqX6QwRe/WNgicSys2ZYl6OQSvMBCMKaY
vjXS9V1oGGgO5GhCM8CrsXedB7BI8iXw356o3SVj+YCr+2NG4tR7ppmCSEXO2qHs
p0BXM1E2whyJelj6KKtykzJSVO/UX/O8LgPyrddkpffy50LvCYm3JslTbcO0Q2R2
/ZnbYoDaoQS1UjObpRZUmXrI4oV5Tg3RhGa4hZ+THsVHMw04bYJdUcLD9cx5I+uW
VSd7osvvLuJdc+4p/RQshkeWFmd6kjMJVndsopcEPr+lJirj6daRX+vqGdaLR/hz
nNaWnIbNe24wS7fVxbZfGt0Lah8wMvFPmZLJs7Qh4Q8Kf+XrbMbN7k5Kvi5Ei/Xs
3/SQDt3Ld6eNZGcwOIKm/VcC0g9el1TkBj4J4PvLo2eWenokl2W1SI9iWxHR6P2M
5OdO/ogNtvnTqUl0XrQ9I29434ENwliRVq5aE8tYfBev/FobEvhW/ch0heehITm3
OjPJDu9dAArRg5+qtVAGxSu//5BaUM+wW0oQSYy/Dia5jRuIkSN5aWeEueZod2Bh
dYibO7VB3aLw8+J3CXREGTyw8LmG+nU1XCHzsN+/dYbEVCVA6yrMajiAkmwQL4ut
7BAA4rREZ2WTg+RjujdMmBZxnMxnxdDycZci8uamK9K+Zyrq7mMHRKLJ/bOW7MjV
wBIdgpICx/nuycojETTLJiMHb/7pzMYmT0Pig0NUYp6GA3jzEzTBzAboOCAyjMMj
LqVcz/tmls0TmIWSil9HgyNDqZ93P9ytHNuVNimZ5R33qoi/MXjaggBKairgV363
L0zou3mOLpi3siRWOsuMkR2ryQXWGx0RV6eikPKqtJCPBp77AvLEDwyn6OEwYia/
D9+XbSoBwA2R7aGBmjrxJxecyU4cz0JpdhXDElgmBNQYsIalohJbvbo+7DeN9RP0
XFr/+Bxc59iYWshZ5oI4y451yVGa3xiSSctfU6VxyTeX6lp6+BDXM8VYPEzqP449
p0Mo2Tsv/9bLlG8E3PXCgXjLDE3jOAgI1OFWD4XGhVe075DvSGdUfKif+3Fp8YIz
k7+NyFk6mPkxDvgk9IG8ab/hfiYc8rMtUIVUlJf1LQ0QkPFK9djuqCTf+OJkY/Bv
qVxg8Okf9sA8b3xU6y/B6cwO+BjUCohsVQ/bqL8vig7rFpnlrqoIjkKJ76Xn2koL
ZiNPAYF22lFdz16VCmct1w5X/4jq0TYYJDf1Duumw2BEgR31vyZQzjOHD+gmZgi8
OlHZpR3DwbDks86bJvM7xTrDobRSMUEJAUdTkH0JW2BZluJZRgCxdi5rqe/MJB9F
L4nCkHvzyHhy29rzLIjPanuahwaAsUxWBss0kpBZeF2j/urr6GxKWf4uPsz0X8em
4/830xiV2Kgdk7l2KZLbjMoHw77bIrzxPYrE+VjItHNJWYHzxDAnPRPJAaISRZZv
TL7KdymKhBzXWzGOQxNv8BAqAZyyIxN13FjNjO7qxaUHK+fsmx1+5maufg3pw6Es
WBfHwZmDyqa/P3KRzLVHmpejNlGNzjNtJAog/qJVb6HTbJSiJ1r8K+UWwoKdFjx4
E2X1/Sh8tNK49yZdStSSHO8cFOE4HsZF6cu/Z6ViLu9QLOZCY61/KdLx6wLbKAZE
1V3vh7Uo9y58sI+d7jhLmcPOYlpGUwFA41vlV5UWM6+D+of3e1inXQ3hgYapVfRh
nbIVJ8jtgzFeEQ4RsSdtcelk/6goJLcLhT2CDvl2CQBrAZ32rlFJqwdLjGoI+VBY
7ffMfYHoBli3LcQ1qhI34lLgOcy2E/UU5kf3h+1TI4tOJ1fSBUj+nlzVrVdWQnIj
tUdmlqNQY0GRBDIEF6374b01JziRgDM0YGigSFQiF3/dl0+V0oOFspd2UU4H/Jyr
paEbK2BgPEjjpoZmRlpCJTfuZCw5U+sjUBILiXozWV+waww+2adfqDu4/UF6ZDkl
Luy5Q41NsuZS0jMNhJReMLUj1onUpt99iSS4+oM846CKs0f/ffgOMmd2mfcAz58i
looMXE29hDgsre6owfidYzFyG3ONTnW/zXPfOXYCWUwoA/6F08IuJMWPQmrBAJmZ
vug1ldy/ajbZiXpO53qM2fSYndSTGCKD5lfr/jQR3s1oMOWh2SB+1fr3Ryk21NDs
9b6NulXdN9ecXMRT3O6w7wvIh2+NyebYNbr9A8AaKIBYSMSp5CGBUAYP9PufkTZZ
GhetzRn4FkZmAnsutjEQZVhSPi1L5d0RX/75uGWqQUTWzBeRj37i739L+BUpq6Kx
Q4BfRvGjYxdNgUTP0qIgzCQ14mqosAliQG+hN+pqmmbVrVJRBFbBAnWQkxqsoqZP
mJ7adWawb9zf3xiQov6BR7csZAXa2hbcvvFk0VICjG/8qvKZy5y2I1gYen+QoFum
1/4gHyR6X4MOiAL/nwUiKCJKqeblt8wx9zTw2/t3XfVb/bKrL9vo9Ec55rMKbp9N
vJkhT+J6WMwGrSlq5Q+x9lXB3Imon9uegF+G+HHWdLRjh2L/EDJbjTmR9mx2jjqC
s96yL1hvO6qkuBgZ3u2uIYXAHPtAXjX5TloEAKQr6tdgoU9iwsNo2IXhm4hkvP5l
0/ZHQ+GXpoVdECsXZPuZLtgof7tjSWgzXPfJLTus9T0ntvf0UbIdN1PpnWgQKqXk
vn/1+U+3VEw22Oebv5rL9n9SPPLShg7eJYvS9RAJmTNxzm3pb3uNUF6eTpm+Esj5
BjaunWa+f0VtOK2WIbtemyBjj9LtR5fADYVElRCDUzXOhPz7c0SY+mCXHqlPg06F
c9oUcewZhZUmHQ7aQ+O459MROSR7NIlUDZwcVR/H+a3yeRr7cmEtQe+b8FdqjawN
eteW5JbBPoS9JC4zSVgHQzRitEWlTY7jJL1LltqNCqbtQUP9R7MeU1FRhC7YpaZi
lK2DhycOG4zB9g6MhZDT6PHvu9XSlSbAe/LlL0MSGDXEQw9z1i/ljsDPO5tif/N5
8CSNiLtcXmFsJNyKwjK3rru+o9hw2DUcgsc7HMSdC20SFp+ftmh0CxE+G7mgksc6
G9XxmHw/E0IXqyMTNeBwN5CDNkJ11FpcdsvyINm6O6vPfM1jWmjt9BgFDN8W/Loa
kNjX5G5Hrf4dJsnL0J0ZzXLiAbH4SoBscb8sSEFmmbyLHGAXGBEH6JCMMg8/l2MN
chw8qwAGAUCrPRPJfslTG8CaGScl4G6i3NSkTT2HSVi9Cwp5Gthn0RsBwa6pXBHw
36ia/u5eEI2w4lHDAYZHx6gfn9PpnM9UDfo4ZRz914WtUiVVDZBE8/TURqSWohb+
iu7OVCPlYWVjYz5PI21tsJbMINhNjvD4YSvxg2REtkcqkbuO+HHSFa7WZmnCain3
7E6kIz/4Hn9Hob57+NhYTHGqaQ9zE0539ISK8ZzCX9Tdx/84PSZVN/9SgamBX0Sk
/aYeMkFplNcUGili2xzsCx1WrlQUKcrFCQDcZb8UDh25nkeGWMwzXeuiuKcHJmPf
1R635o4R7h6mjszqKXib7QXk+P1BLoJ86Y3pFaGIFEGqb2JVPF59k3RkzKuB/GUf
FNWago5JnMhgbq0rfAK6HfRSz1tQuV2GQTvaYmU/39Y+j2KjPq/loKVOkQQ5G8KZ
FYCePY7rEWMfAyZ/GO3A/VE710rAJc6hJwFaKVIpLyU7obzgSVpe9BwXuMyKl1W0
kxu90Hbcx0dlJZYxaQmVSMBgirVzWP0hg+5CIz2ruRAly0KO+4+i5cjSW5BtK4Mb
SQv7Pcyc+8cBwSULJBe8+xh4hlWHS9iDsLPqVJwoPKiBI1N6gZjxAjDkUGEoKyJf
Pz1SAn0O01YwrCb/Qf7C9En/Bs1+GbABy1FX2XXW6eef8wALt9Oyz92dWlQTWqFh
E74AKeZWRHvZvY9BEU0hJRaT+zDB0dxwbdVDVcsWX3lSBv87HlCe19f0NN/7KYBd
OPp1Mdjg9Q/eZwvyStr7FXMR05sVamdvsZxV1uKt0nwCfAz6/AWCV8bxrN660u33
kDMVa2W9aUMZJL+Y4HWolCRhOlA59H6MAritfLb6HTuuI7HaChhGIgMnjyCCYNFi
mxUHMKhJZQ8OUxAsh35h5vLRvDRo7rb7HhaItqOyyHDly2K5cfxdHbOMD9Hdjd9T
vf2EQau9nfzIysEFvNMruYA4YBS8acQMcx7pJuFZ+rLM+DdOfUpKE3uaqFSG6WYn
hmF1wiWXpqPv40c5ZyRbyWz1X8crwgutDUeMOpqD0qYa35dJc/CC5f66ttKqnDqh
3q+a0PKmcf3IykLGc+SGxwOfN/rgLhU7Geo0Ft52H+6BmSIwef1lR7eOLHZBXApy
6aTPXbU7GZj4uHMkvkOUFslgHWpKe9C5ZhMCS/hYouhPJIDlLsitWPaW6/Ftv8sL
SuNHGewfL3IeN20jqegqMsDN1YJFT8D+PsK9zQrNstE3DRmAo/bjLzV6HBmVeDf1
PDcqm/M/6TGwdLPrjK+063xc9LCuwtnsvcy9OB8PQb3GEM+zqw/qxp0REO4k5GZW
mUBU22OCMklxIYVSrdrPmffmup62xDwsUemgA2Vp6i9DekmKkeyhTXHyYjw2sNaF
OWuP3t23QcvRLEjwAADC/Qcjdy+5CV1tXYVLRB2DRuZX3Ox7kJTBCcOG3X7y+Ce3
Oo3PpARDRh80ZGT1BkplgHh+LOnyVkv+VxlcwSSCE8/HLz+NcXf96crvRWMVP+0I
tIFFrAOj/5LWcQMABlVy5xHEYCgtB8dmbqjYyjtMVLhf3SaCjZo8dyjdFk6N378+
aEASNNXD4HL9tkO4zCzV+MVUHcDHqOO9crO9NbBkY7BkdJuPNj1NDYWOHgM3o/Nf
bZWdkmjWbADOBnkbUoqOAG87IlqfZjLtnXrIBpm4UJlTbB71n8uL9NPpPktSbl5K
nXPsn4u+7oFzbz6oN44g41XqJuNIeBZ7kvIKHnC75KWesjZp1QBOcVSfVRWOUDMn
LcaiCWwVmKozEGFe95A9d7tvKOZBWJzZh4OX3+8YdIp+iBLKITCWkphDiYF5x6F9
CUY9H476rmy4wX/t4L/jcJLjB40ypR023UvLQdcW466ChabJnxl3jYzkaGdW9Mx3
HySYTtE0FvEL4VR+FnRUH1HHe3SXHkggEUMc3jq5utdevc5E8kdmVrfixl4SfiOE
VMw/Du4/l3ohasa1sScPn3OfNzteD8caqVpzLnlIV6hKQjhqr0rNQyFR3N7onYgc
/5X0mT7aLOsUIRmmO9p75g3z050cuFY21mXDX+J5UBWly9ES8t5liCh9q5CZ6xDK
GmutZRtYXKOTKdSBZ9K1AG9uzLbi/lCPFtiVriOe4g1WHci9gn2tvhZxz2Uzjxmy
XqyTAvK2oaNkf5hVArC8h/Ed59XR+ezHXrNf3noh/Mgt0DaxDiJbDuXYujA0z1R6
LjBGDwf9UtRACsVnKQ4+N1goxFmYvKfEsUHiGV4e8AO+bmDjnKdtxtw2LUJqzoTP
vvfFDwQx66XlZj5BCRnLTKSMrtS05YSfO4ztq5tmz4u+mpeykdhULmgYabAula4r
1f4h+PS74TaAqG6G7TvCWsWHy9fwO+sZhkcD5n9hsPta01hPNgmNWLdD8YI1Tx4Q
b9lOMFSU7Tm2dIO8RTwc+D9Tc+j8blt+cYO/CIZfRUySa46JGCxw6HjCHKQY7rpr
w6P1lXS2VVj4rcOKOucrXVBMMVmzMR3pFPynYw58frnv6o5wMW8UTBeI9b/kUXjO
vkNbGKaPpHsfmIPOzj0vwARZf7AmS4OZGAJyLibio8Mhe1zVKW/IEczllB/Ix/D9
cO4vhIeY6b3qIF8+1qC8Ro9hLeyWFa3zI7UN665enjswoHcd8PBpoSZefBDyzL3q
tFAWbXLzyBEmGm+iGLQQ73AVQDPLhCElqREq1meWyykDmXdk2/iLj+Sxbsrood6/
vkVe35nOH7xPtWCoG4O05UldJFuztZUPMHxiitpSjpVL959Q4UMLiFYsMX6w+YFS
GTmqeqEYQQiIiHuMJRvgop26pVxuiRq5KUVDOciT8/Cq5muk3fSajXhvY7HOfRak
G/7R2+posDV1vQ0Os20mcTmqfkPesNjQNmgKxDvcnbyPmQPFButxHWLnl5UQeWI6
HrQGZHo6Hz5whEy+Uc5tvWJY6kWE5VtavBRyE8Rlz3s5OI908Bcue3J3WLEd0BwG
WHUDSkAnPZTQFEp12L7B6sRBriQCSS9Q6PFNrF9bA39KOHqXmqHLPig6KG4t3n23
QXM6YEB2ldTmbxrhDca/2xwkzFSwlzyOT+uWq6GtuNrcMFgZ/0vxO3PgUHg0kXog
EuciluwSquzkvjxWMpqKp53/5xZesWb96dCThr/tNQtmHQaI8/IfdfbP59SVCa8D
U9mwHjIJOhP+UawDODQpPa7blhgrqdNORk55NxCgPgvmI7E5GTyCqF/U4fbpfPCd
BwYHPKlRdC+AipMR9uXRjAy9Om1wPb+EsKrM8r4QsVv6uDT429Pac/MJIx7N4foz
dTgLbiG6Q6EEzD5VNS53h+Z3wQ9HIcku/Qo1ZZmy4ypIKroAZZ0k8YcPB16UKrvv
j+Ews2AU7Xxgk1TpLZm6ovhyUzSrHvl9gd7Oxy5m7jIbk5Hqg6G621WhB4gpLKWa
Jw4lMfKWFYKR9prPy01OjwMO6iQ4dD0fA3STvaq/Wh6AbETuIgmvjUxilG5t/Jpk
8grLlNoTbogrlfl68/KYAtIJbdJ5iCbSTzFPjgteCvOhg5VnWjzLaa/T7pGBZe+a
ETGp45RbyLH+dPEhqHvb15dxzxjBsg5RX2QvTziivH/M/Gy/ZQd3qY52AXq0pD+a
bHkM2dxQhAUxiXYdW6o6oPIQWEoka6+CeqxnsMNOWnBY3lW8bPpooW0wH0fur5ar
kc62yOU86nAzVZ2CHW7SDwSSpCkda0WRoru7AXj9iTzUdMGJWXoOSXM6EIC0c+lL
KQXxs/IR7fLpY8cFTJe6a6gYNQjZ4gkb4GOsQyv9HoorRhA7P43NfBSdNq3/ojSp
txoJpnwS3ufh1uvjg9L1Gd+DLeBGX+kZlHa5F+jp0/ShyU0gWzmIqfA8dMQNKo5l
wYYhYJMqziEH4WD1y5cb5w0mBFsTDLrv11vb2cJPnfTyLSUC01nq6eD6BGXloGtm
bQ1+/oDWKHG0Fdb7pH+imknuWqpoNvi1/qyCYhIXCPG/wfIR87CyCEejrYA3A5MI
9MFIH+AxWKseFUj1c1ArEuY5gphkv0yfEhfwiAcLEZ71TUtV/4iePgh4DuWvSOjl
UvrJ6yx+yWRD3nAqnLUc4Q/XHyKp/wzOqw9T8KhiMuOc5d9U5WrN0mp8tz65Tj9H
zvx2w+EU2uhdVbsv4vP7J0d6gq2YIGNweV70Em4i1q7cLWu326ab+48SbATEE5TJ
IlQxS9C7z7W8l76UR557Bzs9y/dTDMUECzTFWtyBs+cxIcJzR6CTJV8kw9d4YIXV
foozLJPrQUJ3N3AjurnF4NqtJtg1bPTqcy77uDQndOuFdarqaYpqc2O4UjzlhSDr
JpWLEh+zJ23wOxnyZgLDtKsnAgQiyzWBbE/MZwMmW/kKezDezvk5hjYz6ZagtM6b
NBwAH8zTexkUMBo9c+bOgqt2q2wsXcFO184X9KnWxII6u5OTyqlBECgQN1teAD3t
YfgyT8vrnW70/O7WpD5aMDKK7YgbxJathGiD3/LZmPWUYfpZxJrLnKaoQB/VFDL3
aQvD4/0zJvIMdxsx+yDgVzqaRuc+AKNXP5PY/JHrMdNGOkOUcm6Hs/OPFmeI4C7/
LQ1TKYwH0I7/Ikkt5QfVtizf82Mcyz+Y8tkAA1o106RKC9c8vQ8B02CPr/2eSnxa
OJ0ElFZ93vMb2Jj3Gcy7/g1DnB1GpMB4N0UJBYd9sKT27F9JY9w+2OqoR44fbYHR
7MAiZhOmyLrbC92AeYQec5vHYSBlWdhCecAjkYY6UkZ24cFgrPPzT41yrRnRR5sc
PQKSXH1xDEG508BpfQ/GCHPfBk+/HNE/tBsYa9ouBLOR1VRz2UXnNjzuiCcY+sfq
UTA1lO9odDaWh2ngp+DDtfFptdy7lfBjlm9HsPIo0LpKSjZIJU4JY3nIPB9Qi3s2
MglEUShIDHp5DYbQY4sIpCR7M4o1t8iQ9rBzQM0FRfnPNy1eMFEz+vICAHy5qa7M
ytp+3knNm83SHJOlTb4nWezdLSZZu4a/LuH1vFBmyGu9Hbq3lhatv9yAPrXpWHmw
IfSwCWA/oFl8NM5PdnhcsDEC1ewKHLNhOwrTq9Rdqp171HkmQw4GmZZyIEk7FrqW
Bd5liLzDf2FSN4ILqme7vZxt9kN52CdjO7N36pdlvXoPJFTYowtJwvLw3HUySXXg
vzTHpXOnf4u4hXdVieL2cffHa/ToNhD5A3GgvurKmiGl8RgPiFb95/Lc2pxIqYY9
0e30wgQny1fQkPSNr94yASMIRp5qJZtb8piUFeectPQqHMr96MLIJi6KvW/4rsa5
i0V+dBCf14Bq/4HkgVBGQlvYD6NI3N8nnHqJlqj2Jznnks1J7hzTYjBrvsZ03x0c
8d5po8ZXoTK3z2KBE6+l1/hdhK8zuXeZ3iJTOKgrT8JL4bEssSnM4mVywwhOxb4R
7CqXxEJ8XV/vOTVVZdBqG8ZAZ5CZIjJTfF3iI0FD4Ez8b0WxmxLbfT32ac8KCtBg
q8YBqQBnxENNBnzhpeSTGQ9Jelrsj8PpRIMBDwWvA5oYQFHuYgiTFo1a9Ug0YOJo
YNgk7J7+IiMn4tgTwjESlMWoSLE31TZGNOXGGK8JAzbLfUHATnsxswMSkRgugEIz
RcAx6PiZT6GkmWddhB5kcXh+R9opUHtr4hk84PPMGPHJROsR7WfiZUOu9QKI/bQ+
pWlMfwSpUao0WKwU4sUjBR9qTHwSkqW7H6OYUeKnFoRDe2wf3E3FN3UNC1fSlHrP
QDBJbl2mE/KGmJe2FFH0aEkzE/jzJvCYyFhyKkEJHbxOyO5jFnBCVI3Dtwywi0ig
vqZrcoUwkdtY2FdE2HAZL0ilQV/6T56huyQM9OrxOUsvjd9mMV+/DZqG38174b1I
vrHnv1H4gMfaCTYD3+nR0LOSxVCH1n6e2ioDPEQ2iGHI9uZVxpHCPya6mOIHWWWN
TzvTBuDbOB1siMm1Oi8JaaM7iA9qCibZFm3hwKHLDa8sTsz3OGQLo1i5N+Xen345
xz32jj3L7fJGssWgidYnsq61HpEGujCYTc0jicIkQwuggF/ZrWSXwaFvHz26LbXV
3MZ7iO7AzFvm1PZ7rl5+3DakOk92GTpSeogxv8mYlIcy8Y/W5CPKoRONJbpIz/MJ
9r8/1+ZqrZfKLjRXYeEDa8833QvDR2ghqfJ6F+klfHDZggh9csBKC6CpeWxr5REp
KIm7w23W/Gnx4aUNvwk1L17zSvWn0ipjWrGslzZXyUd4CxkeO7IfgHPgUBw23a1s
3kigMzPqEL4zekfG+6NfIJ7TJ/mXuWS9fygiDCIzOkF5DuTcs0UeBdeZnljgtyNO
K8AvZ2WeH1lo1ybRDKS1Pzr3XlXJKq7JgKcIU0Hj1L3gLRWoj65nXuttvJc5ctwA
sfKPZ+sIEgQzbrMqKvbk5DCghuAMgZ99TGzF/+NJVR2tArpQmFGNllqY/hhG3hp+
aakAaJWit1HHb4SDZErjWebLUPnvntKtawgIDstkvOgAWrrzVg38nOMDY/GfLCgn
P8zHIzmPwtcVQyfj1NjGOuR89MBoh3JwWyM/5W/F/0+qROSfSUW9eq8OBbWZBA7o
I6LedpZk8ENcBL6ngTqbxENsB4dZ3kkpoeru3NG5JvWMz9bRKLL8kbqGQHFn6SCn
0yWrrNP05aXKtUikEmDdUjlTIIbibhDMHgLgRPaIc8ioO89f2loJAOvFAWlEPVzb
kK2NurwJOYIN4A+e+1+I61C5nr65uxIPvKhSOjQloUZoyj+vnzftymHPBKQ1JC+T
tkDU86+RX65Ik3S1/Ozueg8yF7/Yy9npcYinQnqx7+ezVTpPqOb8YKsC19sWr55J
8L+3MiJNQGoe11xp1ePlLKZAp6tTirv14UxcD6Bd4h0mYLkgfxbcTbKRAz95rTQI
PV3AxSkrXW/+nfa6Xk6zD0J5fTNgZMrJaL1nN/vJAmM2VJbqsoj9ztoFGtoEtv/O
vGIidqPVLw4TWXdWjRCW0QO51i7ZCznePKiHtlxCmWA8BfiyHIslHUESbCtMRzpS
VTyOFg137ywET1MaoGqzlN11lIZFEjiq6YkdiM7X2QHU5th5yajH99ythgJ22gjE
Pm9eAXOypjFDiNZSS8C5yx7s0p2mBIMVbzaEsTGkLY3yHRDZM25VF6/vqa1AeqsP
aUM0dK01k9MsiRDM5J6nERXtL8abvi2XtNZjeVkHM1biFeyc+sKZR88ClzuvB1Hj
Tqsb31yTeST+3WDC2VoP8WZRDTFRx/d0B4ZjmfANDvxUqc2l9yqQRICEFO65Eeej
DiqL/hMw3Znb2BC5rNCRSuKdqO9QypD08oVocc2H7dF3FhaldmwVMRN2MwVxr0p9
z8AEDeTr9e7N/wRehokAIpbRJ5ibPy9jtnaNQFR3ZWpbdP+RlD6baLCvaBpYgtzN
aW9m60++ASE4h0MArY256Kef3hQcG/kkyeqfof/Z0alLbB4r3hkJCGj8vMmQc3IV
G5UA2tNlG/0SucUSloKx6s2Y2yv439/xaWGD5HST+YjM/rjpiZmePdoLi5pqp5Dj
+XfCyJtx/QIEe6bP7a48rgv0h2WeFigvRtcBeOclXxEL9bk9KsU9MowyiQyf6Rno
oB32wOjMKW8SfJbejaUz1dOwx8YbKbBjE2MTuM2JDT11ccG8b8woWhN43FWVNDhw
ZWzKPtW/wD8SfPd67jkjrJ3ORhOgsiPfwq3ZCac3guW2mtqQ6u7BNJl7pDHBMdrl
a39xS2x+M3ol0GjNULcyen3o/Db+mLy0eN8f42IvGNUhlhvDzGZzYIkwlDoO6qhz
Iz9il6VtfHqmv+J8C16gexrgkAcfwtDu4n5I0r4NNVAtanuMzRDsyeoFJKdOjLzU
esubAlE+UCG5lhSZcWv5oCK1tj7Z099wmj7TwhNuI8smNRVQGoQNKidh/nhqYH65
QUFHcLTPxa38pzodUPDs5ehMGPrBTWELggr7Pky7sSpFSKV9vhRsFY3H8CW4jlEq
G+87okWJ7HHbu8yIFzQ5Bn1SrhJkEPW9wctmeTkBj5NdsZPRkbcQN+uMBiuTimkc
5ac5eUlzGPJ1YJzYaafE+3b6cbniAK0LW4GWf71miPmPgGMaqFEjHW1re9ll/z+M
zml8xtr8T0XysSO1PV7lC3CFhr39gF5NT7BpouleEGwFdlhwMdx1h5Sf47CdVwRz
2Qw8B8corF04h42tj5pF8ijzj81A582dfRxisA35pcQUVYtbpvxrHv0UTtxMmtHQ
2LFPVH1huhGDTZlaJgw11tYNrmZc9hx2sSBbTS1W0ZCtsodxyC85qJ7dNYd+P5lc
Whmso/Uk7jbpt6a8ZKDZod/S3e6rukfYWFKnift46M2hD/tK1ku6QRIwsu7U45Cz
RkdNEJQRXUiNdpzoAWH8EYrM8QMqpLqyRJY5psQQQlceoHiR+o5I0jtm7SIp+Yq+
ZSKJPKwnvkktnJbTDyQX7oV3u3VKClVKMep2tNQBO1ilH/OiRXVHiC49w0aZGkf/
v7OXm3dLF1pQTCITfp+/0eAGjeZpsT+EvGNwpchmsfQnnQVaeAY1b1NoQ8OJewjR
Yj/xqXU3WMqR76e8liBaUpzDG5O7NkUfDbHIm2WzoDUmQsc3E7cSURJ50q31BkeX
y0ZNHRNkxKOiXK/Hh+X2u1N746AEOgSo4/T8IKvvlIv4fbvNy9UL9TWi12atS6tB
Yo8lOOuHIMvje2ShcxeQxvYsBFltpwSTIpugPAyFvPMh7YSMCdsW7nx9Sn8iAmyk
b0G1xVp6xHleM5oS3x7JymIx3WjX9OAgcGtsVG1sDANc/HwOI+8SffdGDUVdA0Dv
EgiGvHT69tinGBGOe8bSiXkOOBMSNvVIeIZUkfU1Hr45GcS4vsjvWisca2yKqn2j
91LZqFYdBpmAv2+pXpJg/yjqvwInFc5f6wTF9aWvqF5MFuLpACe4HJ8qZBM0FPuH
2MqwK8mC8M8CxtghFF+Jqrz9gPdk70rUUCFVbZoJ5nF7yjnCHw4kJjkPI+t41yE5
D7ZXtSDp0PeWH+Vag7WUUqMx4cd+jACdtTSxH5WiJTN2gehh7gIdHR2IFlCsmMXH
D0xXjpgEHkRx1G/gBrGodf4e3XGhZcHmJ//OKbEeJYzE8gDn7jsar1p9fEtwfO21
Yqhy7cVvyyMzx06dxszT3Q5lDld+XKQ+wl43zOYwBryTTcxoPvHH3wGUqLO0s0qC
LjfyGmO16Lkh/olCNOPdNHmd6HPgXN2TQzXHkI9eB/NcrIXtEeHv5XZGS2Jn8P2S
uLBlASe46j9rSnbeCiiOaCmdW4nzUjd6Wqngccxbb4mSmdWJE9JUo5draN0R3tt6
zfQZMJ3ivoJujPq5dObO7OlhA6As70SGu/Ysc2psMhmNrNi6O1vY+l5MCn1JaSCw
zxAoa9gSDU5ix7qtUc6LvqhzCmBY5uRWBzUhl22smldsXFDRoVWHuCCCQDqVvCb+
syTRJZh8mP3d+8mUjIj7483PbRkf/AvCuBaSAmgH3BgLvq+JTj4wITuTO7E0CW9Y
w12RJ05INCvIykrB36/HsCUBPiKqfBSaBvG/E1w5jHV3pT8m0lUpi1gHGDn7CDbw
b6Qz+cmXDdZi3Wal0LWLieXp5ddW/fW9trUpZ0UeRP/5Q1baXqgLyCsOSX4ef5pw
+l8nknhFrQlppWcg7VqygwQCsrzjT3A+2aoeHMTcXGO3uZ3IHNb9u9TfvvhTRs7f
M4nPC5KCurqvWhifLdPH1nAYYlJUZjTrhhEgOv0X8yyxX8wpAFsFTe9xaKU8Sa3g
AX+jX0n/GzHXhyvgCV61sX3zrWTfAoTCkexiproWHcNdvwfjDLGxKNYJRcYaUEhx
Rof/dvvSt/E+UbItRmpSz1boYn+iF3b3FUSzLGtcKElA/vMwa18d5VplFJMQHI9Z
eC4OewiLTzTFVHaKnpLKqMSMR6otjrYDKoeCKJcKtcxoAOmnjVhrhuHB2aPT+MZ4
OVxSCBOnUdYPRAS8pBqOq0tO/s91shKUN/7GGypDc8TU8kOU36bJlHpVEEN5DTLJ
9+QU4EahaFihZHh734k8Kano8yf3Z9DAOxm8fHCTf60J8Gmc2jH14Bzszyd5nLF7
63wzgnBSPyEHVUmF2oAvT6hANg7rafNNuGglwbp6apb0lyrA16Twi2IxIwNupdyF
LFitpE8TlymTT+UlWYutfqAcEjvtnYntWPM5TdQuQzgHHQy45bv5VYksIx8LHcXV
W0olJaQRFuHfM+PpUOvG9+30d5xWapolEGm+6gjFBiIG5sG9jCD5cNe7dnTgAWc2
42PfMdO5xRB6vjA5yN6EAijCbQ9QlIzxNC3gxfA330KuvOo/MOL5VWWcBlHbj4VF
n+CHB8hOdE+k4gbRPeb13Dv2yuYtopjLeDqqERQ99H7n/7yrRDqSHTonzayKXZ1J
TgNVjDNO4YdTNS5gSCxQF13m0sv5+8UViAZcusyOMkxJKfuFVTXWRVCFb6fqXM/3
65AYlsJy23y/O1y0qVPHspdM5e7CAbo3dtPj5tOJzmg4zetOeO4R8255pH/7FP75
brO53LryxOTzHj3LXJbU4zmMxJvr9Q6vSdg1N3AhV9NNkkRnaaLLMNaggoc8CcUb
x2hXbeJlCxgj5yw5vSp8WFdMC/mmn7E6kj6OOv5qjBIgJSafaRQyLi1qLDDn7M2M
uJTClN4dlfLJSBxms7C3UBLPFBRjuBV4wvmxsTQyh3qKVynkRWLpeb2ECiuhaIYf
GInYgzZ52VNm2YJMAcgWV9nCRgz8H5PKYY/BCK7WFuCYFf3QQpjjQAiAZHKA+wnm
atr8XNhUjRqbEihC0AFnSedfT+u+mHE3OHitfC8vjt3wsRKWKcW6uYp48+CJN3Hp
R52IqUKG7uSvP602JsBVQ4evHOOKOXJIRuEVkVtODRIaO2XrhgUy6usClag98ylv
RqH7eOXdwZQ5nZaohTicRrHxNWlnhqeFLlQ38RyMHYjFU6sQYDJgug5GFPnFlrkg
+eqhsHW+xzQZ3WiHXdFxBfqbQuY8o48MjY5qQVKDxtxzxvKxmHq2+qg0j8lIoKUf
A1TBJ9huZE2YjL7alMsx/d9BucM4coiDImfuh1Sjy286FkDBoqlnOgowopM5JIMJ
8hQbmAMVU0yez1HFoWMBma/BDETlt2BZto3dudXwTVV8yZLDHnmCy/wiq8CWhBNC
mWzazYLDe24ics22y5TQiNXjyIatMC1ta2F6JfcCIj8b24PmfJVAKIE311Cvbyn5
hsh0ALV2nTX6jYztKdCeEmeeKWdWaMOePsvSSUzK4++FvbnB6tgXvvIkMnKb+wMr
n3RfB2sNHK6c+q3R2Pi8+TIOrpT+qK+5ZlOytxoRfjBhsgpdGZPXAUmLn4H4rOlQ
XGLgwlLt44fJOmWSRUlbcfNQkkgQWsUqSSlhWxAD3NWXoAd7/hnynTMkO+sD/JlF
ejw9QtRkP5VFrEZ3gqY+Dfv5u/udsY8U3bfDJWVNArl03JCJVTjL9HrWALGKo/ZC
fhMmqfnK0XqmkJcdRfetRDzQ4SZAPfkVowF9dKXrpH3gmIUUMHkdjezS37ZRF52z
m1HrJ+wbbCD6Mml4p+MuEfAO0IimsTOdmFdU3KecVzmW8Fbqjb6emd89pHA1UYJQ
cNmgdWu0qb8z3lCmY/aoy1C4Zbht3gUaOtd1G11yLGXXNrz2e2q7OgdEg8zPa7BJ
CoUJ3vXQuIw1cGddcI5+Wlk+q547F3S3Zq+3E92Qo3On5zyWkSO0CP/Wkr2sRH0U
tFJnStTtUoq5FWLcszCjbpZAyDtogbf5JO2i+duPzAduqDm4vGTYZamZLYm9m/3T
i3R4437gks9Ty1IjhkHUvzx5Q7TAZt61Ut4eaVv8ueDlvxOQKE9SXY9AFivvVPVS
E/MUbJFa32lztlhyu++JSGOFDxQNvh3X85yU1GOmkeWdVQHuVCVckkrceQHAstJz
XswNr7xuDDrn0PebjnxvdHRAp/5ip3quwy1czCHbSHkxAzmGDuyjv8b9ufUkgrZV
h8C9c3xiouVo5dnnOuRP1dWQUQ/gKudq4RZqeplyEDcatrFqePk90DROMpXl9L4h
I+D14wq/Pn4W8ombwDC8shiAzmMUKOYyo0BZm8j36WNY0aoFqB7UIqDOET0D5SIa
UcSk5sSII7UtxMHhW1Es81iy9LeNtvFHmSaaCNADngllyD5iCcmPbgRHHSBnkpwM
Rhrkoxw/tkrlNsk0iPqB1iW0cnUgjWH/FE0UlUHxbBTILrYFSGcesffja/j+07OV
9PcHJGJjseGsIcJEGRt8O83+NGwwlmU3fU0+fpXoq9L6gR6Pt6rcbEPIkNxal/Cj
WU0qLClqO5y+8L5BX2axXjdYtxUU3cG5EQbHNtlygfPu6WjZshDGBBnVlI9v9dhp
69FliG+6GT+xX08zR9kH+z89eyjMxHcMI+xzY6VFG+vZI5gH+FhMa67VhH2FKjie
75kBARWbjKM7FWgBnyHQiqQvRRR4yaeX25lx/HDAbaVyxQxl8Pshb3DzdNKLjaE1
MmolGr5UMFi93b8KiszSnV0rpSpqJxT3ozBds1ogoSmcAIL7/JhLIjQi1XoF8N4j
YXi/JW6IfJkw/oY5el/uKsd6QOZNmkFTIQiJAM/ldFbr6B4UXNE5A7KRr4tfF6gf
yF7rTCWYHK9iqSGVaRKXdpdQstQuLddcm3lCqHdmdmDM+d7QV5GMfHIjHTcJ8Ef0
5wMeNsvmAyJIGLokcrQBVCOYVkp8cwD47glNuDugy4wSE2NoDJKLb6uJthhsWDrw
kCjdY26sj+7jBwgweQxCTw7wjbhqWxiqlHVjD70Hna2iul5fl55jSJLm1qvP7o3X
xQt1Fyye9OYbo7y/nXZ+bjc+MW7RDRvpZWP1e0iU5mnWeVlLsrajxn0KjjrqkMVu
gUhnstNpa0ICS/RYspveK7wwcJo/7kKZuLcWWB+K5lO9SL1c0G6FH4K9dFfM5UY1
sepSefHDAu089/3e1NQQ5JRzjMhgCOB+/zCIFwvSZ46buSfmqiKhOFRweeil0Qyn
+YEg6/dOSO4SeuHapddrp+VFrhwB7nL54UHFbNrD1KTJ5pULqbEZRvXmGsytJ/3D
pedjNMJBhPpNYJbi0CnlVUdJ9D8loiFyeF8pSKN+F41yO0o7+kMosdiaVaGvzHrs
+JEQs2hs6QRvkhF/U2SEb3fhRUy5xTMIX9fx1a5WD4SRxXxzKPbEDxc9jYlXGsiS
EUy6RH3zzciCSNuCnN6OlWtEKYlbYEw4t7IoYBduAV+wOtMYAPRr/m7vR836ytnS
XEOxgyDrCzegXOZVco3bwA5avL/8GM2IFxOEJSHvpzFBXssmbhbvDcDXeU7tVcO2
aSJyH6jAzPAUiAjPoFLBBas+3K7/s8TIydnJlRzAAyAhf9XHoFtIrtE1SqaOXt6X
vCQ/gCa3O5RiqZtcTYjToGgPt4JbDnYndYa1h5GckiLE0MFf90uFpach9Pcinwcw
ypqU2Ul/PctZUvjrzal+q11hcTvq0YupTKBvH2+nVi7pQg6ew4z1+bGwhtbP5r/H
vPCeoSPGmg0kvg9DmS4i18TzoUYPXafvKSSIMGY4ljga7mqFlqHH7GD82VYXjngj
1GizVwhAsnvJwnQaZpt1jCKK1hDTv/MR7UGMuhOaET2V/1whEB26qp7ezBCbgeb0
/k5IAxTXSqvDAtdGCzOaXQHJlwl5Z0Jwz2StSm0051W4Sk5IGq1oMbQq/P4th/91
ezgRvXvexQjlsOoxZUIh1GqGyVsQWKHcjODUETMBrAeULREp8kRWopmyElVIx4g3
bT5xjRg3Fx0sezuSCnUvHl/OGaCjkPxS+VklYaCvFWYU2WyQ6z+TXnMIv3AHWYNZ
JQGyP9dT2SAT7LCDC7D2lm83W6ZNJqVhbT/j55zjpQoZJqSsx62wxCfhXEAhrIpm
W83hRUDPd9Bsdx8eGYntLqpIyXkOnrsx1yc95jUHn52udlZ/z1ccwsBgKk9cG2hu
WJI7CaD3AAIiigecngK3dN/BQSp4aSmOnOaqGAUTXdtaeOiqAc8wr9sjIDBwKWlm
ldj4lvYhsjdKX0QaIa1mXVF5cpT4pv0arONRycuCl1tyRUPP6d64NrYvYCtx3Sju
Mjrj36vDklmqltdOsIT1vRkiI6QzfzWVtIFqwyIkyabs6zcT35ksAMCaQF1+ZoEK
OXcC9EQc/j4ZbsGp2d1QIVkM7cH6gon+gNEZLeBhNQLGgGScZ48/EhSL9fmq2/co
ehfnbpoopmV3NmqzFctIDVEAYTa76o0/g9oBUkBDkTT34D/kNdQ+ZJ8YCNZ3VAPW
nURpzC99I0z0EtKXZ0i5svY2lVzLA6/lrtECsQ0VrFGAVaxLGXW0VHFcMoGXAWsk
Viw2zLYNcA9/flPdHTm0nB2zsTT6Ug9iN3rOSnc62RQm4baBfuEkgzqQRSjMkOdz
v4TbbjoynQBIjjEgLBCREDFBtxIIbzBjEoAi35xLxon3QbE1VODVIcOVzhQ2EJ6u
OkKvoS5mFBops4e2KeFEO2W4rV7I75A2koCY23YoU+qTlPWVxZB+v4RaZwo6V5Br
M5s10BzOFaKh9ZDoSnU9E2V8BgAOXndjW5JWNU5nFoJInLTWG1ROftsz7zZl3SHR
/wHiKFL1n19JceebhgzuCRuLwSpOqFVjrCBhkIIcVlXCcCUtRWjYHdsREvDXbiv+
SR4AmJ3FHFKWQ4ahtNG/+iVl/MLkLfJj6Nuz0liHSf8d32RUB53pnptwL5OqK8C7
hA/xfAC0EWLRKCTT+4zZ3RcslOyKXjGqiVf8pOHfb7Pk8Kuw6Vyq55sHXIvAuoQc
/BjD1t/NsAzXhnrE9rFj5ygljc16sThi3yZ3gt0Tg3utZidKLXMcQgERG1h16I2q
fZ2tqWv0qTTeEyzDqFRNDkz+gmX4WSzxqaEyg3LUHJ2oSu7Dvke+u/+cRqKgAKar
LL23gYckHU7q6eNVEk0XOBEcDEUAoihV1JxdGvGnLnYmvNGIFD5bOzJDbVPtdeXT
bK0g7Ved7C+yN85Em6eL/42UON8FyOcmb30w2v8PXicOr8l4cPMspoz76mwlyn/l
qXXxv+gkilhSxPO9J7hfBDsSMPQSpZj9Hejx2pbZVsJCiUzlzzrbNJQJfn3+BsWH
+FHsyM75wT7rn9lR2MK8P4nYeI4ruGQaxDrxMxsgGXzpiOKFc7x2Ty+56WTkD33B
JAH0rF81tvp8cirW8XadKItpOFbFo+dKII+qN9Y8GEJLwW4LDS8bBip5PscVo9P8
bhYdXHC6/zvvE/mx4Mr84QK5PqZ4XFk1MEzGD07aOspHQ7FXa81tHpnR27NDbels
F/+hsnrJdvlyNGvJreUUaE3vMDYDpERjDZ5TvIxL+/C1JlgjfiB54dg5CJVTuRjR
koNfwYb6+34TeIIXJu8tzqean006XvB4ge6WydH3YMuN0ipwabmoihn/eqWHnWdA
b9KkG0FuThVg/8g0kMzV143edrbxF8pQwrnEmZtJTPYFNRgZkcVM+/8KKP+v8m+E
wZrsEfajJp93zxb53/66L3CFHK7oYk/b86QAegVIDZnLQY5NqrXE1/Orn0+Hq3QK
OA2xUvYs3FDYXxX8oSpeq3wNdg6wrnVpsvZMKLJcnezyavRz1ZZi8ju2R8Jl3uI8
09/HWyjXUxSO+QDBucx0pM9Leczt3YkHq6XZCpq8a1K6CoiqqKSRjVpCYhgz9Hg1
R5jKEGCX321L5p/Hf+P6/dSugINjdKpCgxgMhMy8+FX9OrI5s4PEPA8om6cu24oU
iV8s9D7Z868wwFRXVN23bZu0uVPatze+gVweg993fe5XDcj74q7t1O9VNL/ekKDQ
ItWS4AKxqaSbaMFnEIOLOk641rjq63eKL54py6Oup0lpRi3XSjwRu5NZi3mYlXpI
IgZY1H3s0+Cq7K/mY6Tqa5GgHvVb8MBVMMGVSqsj16hXypYg48CHxt+RGRugIs0g
lvTdKp7iVEPvcQaw9BiYAoz9IEiVV8+atbjsDEYR1BnNUb42vNmDNqcTdtjA+sUr
AzEZZbWo0h5lsfz+XKICeLKibF96gVJCxqt0i/IaahRYyGO3YN7XRUd+VOIMYe5n
2g6KC/mIfdqSn9n/xOu7pvNkARSwdofoHOAmB90F6tvgIiz2TE0adcVgLBnDpMxU
RhsClnbMj/Mh/OGfZAU5+h/PBinvhChiKObx1fvsLOjLRhVUgFGj0lF9CltuC1f8
Gmg9I5dF2pOknSauHkNY44Qi7PNExjLnelQYc/GxasZmNUiJA23iIFKA6fFETyJ8
Hc/425Eck9HdzJor12dmTm3lNWsbXxxArNfGRlAHwdV/4Bfz+qiOtAVuwoWHmlx1
fS+Pz1cGO5ClzCfplyveaS1CYfDAyLOCd75Le+kxe4skR2ziw+T77oGpUbN5YpiN
w5fgK6oOZsQSeiRGpKD78mqkr9Bc7LuQboQeg/Vo+tkGEaB8TVR9kW8a4mMCCIPQ
31Jj1LrjzJ5fdjS3BbOXYCTjh2Vlp3rMjKQM6Awq3dbC3WFdqYJyWNGmrT0TWvxs
0aOZwgI0Dy1JQ2Vjsxm0oADlxkBVlBVvxtXkWwjT5JfmxY/rMVbqT07cRqZ/g1Dx
sSEZA37o6r5sEUeF6WgB23DOopV8WPXkideGlKp9NbpmMWle0SZXw3ncUXHLymk6
PuiQFJ1Xm8ZEpF4myjrrRZ/CJQjiDYEm6+QDCc47McqQWr4pM3xzo3dxi4uUVwJq
IBA0Tm7WOUnHOLO268hNSVBWzljIrInh8UglyM+GnSaADjFpdkWGZWjDBqQTuEoH
HW+EbeLN+iKWF9gYevlOsjq6aahlGdsjjPrFhiRFOygue1FpidPsR+rV5i51fqfy
f+S7q4WDPZ7xNOC2R23ZwkmfVVbW8Ri4EgF6bub4T0reX0i2GlFd0rv9FTtiFWOx
vf6lteOCdtfWe6ae/t1ZmJmW7TLVbYIqKgI5QwFq6WBNDsGqrozQmtxq+zQyNm/9
c6Z5gDKzm+anCShRL6jrBfmqYe2LMxdmk/8oAlHgIpnNv1B0QtEp3hJhJZt1jBPK
U6rahXXEeNgD7PMPcWGs/3xbVXbqc7fa42YC/v3r12JvIoKpGxNmiSM8Bk8gOvmU
9WUEpgv+DeX+RqYpOMCA45Xp/eMAuTDpUYZtE785Ej5aeRFSwSWME3FvEmMdo/md
RsvRTGywJ5+hIeWN24P1ofhLarmjbNi/FlGzIjgmUCxFIipa19pEMGh3y1KZXTqf
S3fix9mCHmwAdBsdqrWROEYuTIBJa2qD6GR6JvLlvgl80HAjSb96r/WSXRM4lLx0
XwI5n8pH0mgP4S8fi8z3gtaBzg0FkCLjsRY/aG8EOAUaM14VKUTRgW/Kxip4hnUH
nXYyN4+G4uNIB5ZZJOPotGPCdCLoHCLGhTvBnQWhQn4AbHBBi68g9zhLv2CGq56h
hV1gcRdHyD4qKJqUnagE6enBHCtIquWDoqIBN1Kgwr6lU97uC3H/DV+IgIS6txHu
V9wKsv911aCSkF/i8mk6Yjh7zynm/GzE0La6QT5tSmQY2JecoNNkmtEzfDZKwj4w
EEZ4AX2rQx2y6/9v4IE29UzbKHF5WsfubNqOOFxBgiYbKnKr0BvrXQGZhbmCO2nt
xroHCjYapGOEYzP85F4O0u2M0gg9nZ3VM48j+hvh20tMuG3knf2HfupI7uCGcFAI
rwkbFvbPDoViYatiO1w77EWETvs3iRPwYlskC1ryUcHFalmJjlmXeQpVt1yLJFLD
g6XOWoifQpVrkUcFNT3TSVb54t2HhbLfX61LgiOVeqka1QM1is4BjN+lV/uMupwy
hxfdgXq5SVEGfGkJJf4bET2mXIuauKfNeO1XA3yKucTsLe1LaEa0sKxpMLs5gnoj
9mlKfFcEbszPjuo+t25u/FvTRVElSyIlKPKWnqdEJ8ZZvVjZ6UkgWnNYR9m5jvms
8aIho3fcyzQvuB0gflnpfxsPERAeLJDdoYDo6wImiLv8UenhmvavoR4MggkwZTzt
kMydCP48UABaTWZoomsHJi1EZmZRqlhdK2gaFBkbN5pIFA9GJrPjqgT1F+fXvPsV
53uvphJ/8307zL2f/oI02/l74xNVdoXmyOZN2cPe5pSOG7E3z9TJtMJwjhmlHz3X
O4EcbscPeBd4d9ztFgP6V3lWGq85HH4hgtxIB/seUeEc/FDBveN3kmbSEnyeoL+e
EW0kQDMcjrupCmj/jRFUla4r48fSZTI3q4536URrxFBxiuo4W1UZZV1iIZHaX+Zn
/+hn3cn5OpJRST/lCy1G+uGBvcNaOk8W7s8iu54Y9C0tDmTMrdicr7OkR8OfqHVO
aoY0r1I8mcqhnOl37VvZxAfFD3VmvkZTdLQw8Cqm2F28DyOxR9meY07ZzW2WW86Y
iVOngsnId49UwPIPswi88QRh2o4iwDVnhf4nOlV7Zw0g44V4V/ncRTkZrxdW4ddV
71BLvyZR5t6/tbpoiasvWux2HE3RQXYTbB5LHiyrW6cuXZYAdrG7+jv5NKabFfqt
D91TB61xG53eNSWTI2Zeihcc8wq9m4/wQGNiKKIzsEFvPyaNgnwXgyrCVftCx4Xw
SPKIQ3pOn0K/HB5fik3ufFH3giqeDgLtO7Bdiwjv94/jOtPHDAaxhd34Xw5IGVWH
2a9s9u72q466adToSCReXaSQOTil7qXKQbWC75r5V+5vQW2nClzxN+x0aWs4C7C7
YmPVJ7dI6brXrtbYTm9NJz/eW5TuNkCoBJz6F19uSi6LBvWk/xTg/llS2Mmxam0M
CLL56brZp+JHeFEEJqTeJRqNHHX6xhjZqU1zAnDOwp0xjJpC4Ia+wBlOPUC18dXO
y25ogvsHW5jnVjrfHAmvKKwIUhCq+FGWcI/6+dFNlvgrB1bDDeISo1Nrg+QDadSa
SKGVtx1Mo/aBBF8s62CGaPcVvi6HspgTRQHh49nfAJL5EEa17fOHBTA5LWKtNW43
udCuktdiUcxG8zQ4ZleLLxYGHgXKKougDfy66m9hcKcVnzs3TPOaptvkkiWEFbIh
0Na/SQK07UeKmd2eFZtHb0oB+qgzsZtVYCqo8/Xqf4CQvBBdvuhfJ4w+QA3P7XP8
mp31z4qcBvgVomYLi3SgCx4yrPEZyqtzQjHLg0fiXTseUtPnPpSDsajABp0liFcW
qTtZtJXDed+Mrz4cd/Yg57C+BbuqLw1HTVnbKveqbMn66Y+CnkhLQIc/4dvnepY2
7I40uF2C9gE8m2oEoj6geUjmB/ECyqgC3SGn4hZIhtusBYRnaiQ+1xvpRLJFaF3H
ItWDbOI0l8iwUSaiS9b7h6g9wg4f4DjbtMJ9CgKweR+t815zJHNv6chS0Uu6hxZF
/bywciIfx6scnrhbDLGHYQRwdqeV9e3i/euh2Z1sTI+HKc6IOQeT8fgmovYmjlKX
V8Om8atAnWU7yR7UGO8HoEXRBhPCsYTm9RJDWVzbSFU6t0Rr6eQC9F1gJ7vTUamV
DN0z0BakSr2uViE+lBpshH5qXgl3TqzQJvyFXb3k4sSd7KNPJE9XuJdYmHyZ7xMK
GH1HoZtzn6ST3zEZjWNToYx4bqyK5Wf53F92fw6wZCI7XyjZapyGsCEEa814FPo/
Ui1HhN6G/NLuyX2iwiVQ+H/xM6baBzxi41tG+UMBw5tb6HxsQmUMtHjWEyWF4XaB
DqzaXsfIMg6quDMN8Ud6fX6ZhRRma8wTk9ag836xYa/icliw0JPNbf1P8jDOG06k
TibEjKmmxwnOFh3ubxvV3h7GkFSP+mik9DdBhN2Ah9R7GSyV+DajMbCaHxwZ+pVZ
HItdGPOIx8x/JblwqvWg9ayRsrIR71uvMkG2OA37L12Em6HGFChiVg4PMI/az7SV
HUF3JGCRfS8FsglCv/FHdgxAOgXxzRizQJEfHEbgD5fbuIsC6CJ+MDuv50fPf2Di
YV3Olht00h0YC7BF6qzpoJsJfv8FSTnMDVBL9senUKToFnCXVBMMi+9FRUeimTY7
Gup5mwCNbvON7EPRmEf+pAqTWq6ixCidckBfod0kBaa2TeAK+6bbqldvXNnC1u/K
C0QsCYL0A8TCLGjFltOfCPJBCkLNrg7csQTXpfoqAQLNIHAc/H7O1ykP4hsK5oaI
W1EgiP30f+Bl/OLQjJ+NS4BT3ERA1CYlL85MvBnmtrCMBj/FiPqNFNX2l9WHMHPi
djIOZgjkTg1Hg2KK4Ww2U+EOeX0OPs21iT3PW817oQSc2Q4CWLELc7DRLG3qBkaN
uucXfirUT2XM5GB4QMddc0iDsIY5eGWy9c65cSqwYD0u/PKrBfjiirACFVtCrWWK
vkL7KUG751aes9g9B2X3uxFDGgJ9VpCFcHXcksPTG6DyODVhatz/vnoAxXYWj5JR
ZJAXmSZoGpyS8k6Nd0BnrJXGTcKdfXQji05DUJ+EczD0hIGW2SXZ0OcqiOLq5Pli
lFYsg4T6l6bL/2jx3p1B6kNx+Yea6a+XGcWXZMLO+o9/BPRX9PYZYVbWNYeMP2Fw
GE2ygrPIVyChLnmg5FLx5/WvLO/6gSm8n+jwmYb8bgrXhydUnkkrptgnW4WYgtvq
N+5jrOuJ3kzQN8fHrWjxAbwAK4jVcpmrTjC80NW/FKeu4t2+HYPOW+HN1hy2W6Gb
NUCBqarWDs9JOhgWk8HL776tK0Dd0q3g7oWvHUrHRk/wL9BrEeeR06caTG7KCoZI
7qHNO6QeILAdVAyu2hMcmPj6PVgunk5xIJmx5w31P4r41h8Tb0uiRQYetph3W9pf
uyZnSdO1YW6vfiM0jzhOivDeFQ7q/mbH3eczQHM4ConVLjKrQqiQy6ymzCA00dGz
XgP/rK6HbqdozUjBYYCDhgHutna71DvKghJPTsgfJBlyNun5gKfTYwQ+g0+7Vctd
HI3WBnedDoxcapySqxzV+u7qwSB378LW2FhSJtN7RA74w0Eo5ucYeQwbCZijW/zN
Xms4tUG1cQ4E2uQKdfJsNwSakqfea/dyaF6lzPbYJuHg8j5A/MhQGZz6vLp9/gxw
00UFSlCN23PP+5gXl3f6Hx7fjL1g+O3dLGM5QzcOHODgvBEvrV8USQVHPCncfauR
AB1aD4InURAy9OPzuENleKAwxBwWLtupabrqRmLfEcfdJyjX0I9pF0cSUuaWnwSz
hxVglVDcaJlEhBWAWwe3Ep/1d/GdKm/CEXbFCSZKoUAj3wJl/oqNbnrO4t3D2jY/
dIcgcRP43LGf/vlCcK5L28Nzs/X4q+RKL8vaWSI7PVHRFhKZdxQN0Omz8s7Xu3cu
DpsYjxj+gCv394CHTbY7LS/EzFNl5yLV6Socp/UAAOACgkMqWMhkedjwE0a0Xub0
CdV8uRmFxUzrMAlbIeelRm7VHmhr+K49eMWmeB4o9jJwvzMfr6Hi8Sq9K1xNBtAq
we9+0tfoES69EMq80u2ZhQ0fGV6XNGxfti231dLeRjO8yXulUqYX/pW1ZG/XBniK
wsotBYX6cRGPLS7pRq8dsRnhWTnVta6BX2rDmvJ0tzWXU3hZ4f+11mECGlpl5Wma
OPBQa6O/8KK8NsM4O1FgfPfj+Qoyrq1IqlPyUGntLdk5wZdgsBta/1TGkK8/c4m6
SMq81ioArYIlNSsw8mZcTvFth//VOt0Ni00k+vlfA4TgnX3GcpK+7OaxG6ipCopQ
MZJIv4iSp81URhfn6XjaoYor/oQS2PFf4NGGQBWgBzNy/qRwn/vRMo91PCN8XADN
42CTwKQRixy/Q1pTovxarm5J6zDQMhoSRbroJcDgAa5XU++4EMEqVnGEvI+wxa8d
pIv/CiAXBj2X41xSP1zezx4ukytN9tWBG4QArvBrcGkPrO72xlSDATES1njdVR84
ha7+hGLoKQCiqb4mTGaJAXM4/aQpuJT1vB6UIO69HxFzZmp+IsVZuQFUIcBV+Cgd
YpZcpI3SP7/1BRkxVaVDA0MhrncNahNFNOibUc7N6reYqIFMfMB6CS6wE/uDfuuX
rHIy8ootUnXL4f6aYfjSCODtFMH81iuxkpVgTlss3n2ei/6OPti3Em3z/fjF0Khm
qDO5DOV10RDx4Xsex4gjlz6skWTD4AYVeBTv9wrcFNuQWL37b/MtAwsYurpK04H4
Ix5cK8OvR80cjxGsmqDvdal0/CoCwbUDsT/xc+5XiR/yuZkTcGpJbpZfrrC9OwDq
A7uesEDpXklT4IABBnc6bQ4tw6YpI9JXwzHYu60aDPo8fCl0PuftivXVNwL67DHK
lVzFrF+kcs2s09keWMTNXdz2O9eD99B0jbh/Y8fSAQWWaosQSojiC+Ii7pnJ177o
fKxuar88JhRYSOyWPCFjbgRbWM9+XwY19NsbcxKqUxLt8eSpIhTNzrcdsZooY/OR
wwYPXH+AI8geSB1YzShNAdfflPMJ3MK5b2uFByuqnO+RxvwZ0k78W1E+OWujCkHP
9Bkl355+aIvfDW11vkSgMlNSBuxfgBo0bXN42RjZ6WSjQafh0dAK/Z5rejngKums
TXbn4kW6/PoCO5RQMZFWyA6JXUqDX2rzg5i6IMjaA43pkwVkWTbrfSqgsGNob+Xv
+97Tx7dd/kHnnsmH0mwYHWF5nIVY4wxGcaXylof42d/uU7hAYe5BmFVQO3dQ4U4A
h0xxsii/BDXwTcnNokQem1TyjB3WSszQAuI2ngXyRKm0cn79TFI+sccErvByYhM0
vHD7Jkk7Ero0hYZkBYk1MrbLzsPpB7s9YmVYIq93G5MIleVlw7uWQXuqKNJp53B7
aoooFN/qiF+eS1fTj2x1PRb5+fFVwpWz0SefybTv4JS2sbepQzYawzePQgysg51/
khE1eyPtdqlUyJBppsUvjLu6wC+PWLDrFwkMySYzn32yJjVlaGNm6w4croYA55Bl
99v4HH2sgMbcr+TR228AsYv0w7Xe4v5HjzCajClRTLgNiAcTgUiSV39hMRXPXxxP
YNwUk9ThzFp8A7UfzOM9pLAIjrKNeeQDGlHAuSB6yZNdwLE4FC6HTGcUy5PnXc3Y
V58s3pqC+jBxurNu6Z8jJ4OgL2uOfBpDhbAk2bdiDdl+s6ghRM+MRc1dUGpy8ksa
Trhd9XRVo/CzEn/vsRPHNJVDspoZJ7/L8UfGUqVkDsKqh9aPXDd7NZr/ulB+XkKG
8rO7KXToCcq+EJdVPqw9WCuhSNtNFEsaWuBsMEL3rtkW/gOtyW0fhJJffZnUvEha
orSkL7xHKItW2jSEObwSMNWI1Y6FW6JN7tmbxacUnP7OYNYwhyATI9s5uoi+3f7Y
yqK5epTdtuqohVCTKwFAP1X8GTZhkAaoUYpMAJ2pbwIyaR8OJpawQKcSfMN1yPlu
iVA4Gm0q5vcg1yB29cKA5Ts97F+CamZYiadvK8Y9/1X17xCYaH8Q3/xD1zXwjK0N
x32hBuc04M/8EH8ZwlynTJMd/VkDI3cqgWq+FjD87ebdlnLHqy3HpBeb+lIbvm2v
ozBDPYBSc8pmK+GhM3eBh2Sho1Y2CvMcInrQTfufBE/kZNaad4SJgxbsXabJ8rPG
ePH6Jcof+zBSDFNQWbfmHZkZDXTaadpzcIRlLO/JBPCj8QDTGBNuXyqBukYaXbk7
XkxlXwqEzC4jnwFWbDHAxoe3rECbfeTULMDTTbL0VGd4tOqIYf+8xyKzXg6yyH0q
WpSSwatbl3ZS6SJ9MHcoxl6UJyaz7kB0n0vD+IaSm2qLTlUfTVEO1RVYYp8QE7xN
SwXkECEK1Bfsr5LpEnIBRJdy9rPe1giSn98dd4Sm/InwYTbQXxv/4UHgAEpKwfhy
IeB57PlEOUfA3JLyNKBmxftRnJ0ekRy90VMVUbyW+fzjIoyHlK7ymvykonnfSOMX
CiTbjesUiOttamUMzszCcui4xDbFInDF5whpJfGhHCfRIZi6mmdZ/dEPJ6QyUjjM
vpOhHZt2jbtwnx2c8PjRE3N68hkHCem8BD+ZGMCID2++uMzyNKb0yhUSAFu88OxW
CSz2aANze/N6jvY3IxFwpz3lRvxlbRDkGt1SgLjD+Lo94DhUXTomI6i3D/sw0rbS
Vw9BlGzwqV49pq/pwvjn/0bxL3X24kYxLcaOXgG/igZi+t/P4CSPZnk0Ui4yN10V
I1TdrDTrky3H7BSar/0os+YauA8Ol/sTfqfm+NzDBhqfufwLreWHX7DeAYLZAX8A
//U4pEglkLV6/KD59oSOXjm3qEJqTYL+9CqqJUmZe3GW0P1BDmjKMqAhIUIGseM0
MFHgJlKadl4aIKdna5N5Kxew+c0VOvObsevFs65vULGxqETb39zSWPX/FwpEmrVM
WfUnFg6NHvFmeRprM99Xk+y1f/l3+gzAaUMcveKYFP/hRrnmMei6b7ZnK4cOmhva
bYre+er/324ceJQBqwQs2ANdd+90IzJIc7LaoSKWuZNIvhGgIgrzor46Q6ATAESt
BuXbSNAyQdAeKFLUqzbeFRkoyzc0TeiZ9zLX6xie1idFDtQ0laG6PHZ2ZmEktbvg
bny2wa6N7r/I5nPTpCV4BnDlyMmEZnN32by25l+Su2N7d8El7kwqqSq7FCCqo5f7
hCCiSlBuPsn1/6C6b1Q0+8IN0uTZsC08K0FeUgBwcrTghRlKRQUKO961/TuL58+3
q6I2wLE5kwZSYMitUxmD1irMkSei1mVWujFrSCEPqwntEUwcOlv4vE83PKCF7PbH
iqIl3kbB/6DfkEXVThKr6XB7VUjmDPYxB5vUP4jOYplWYpO5OepEfIBt7jh7f63v
QjpA93kZayHwRImU41EnMhN6zfBCOWk19+Pra0cpSTIHJ6XxvDj1n3JUAW8m+HxR
BJTH+hTOqsEw22BukSeXJOX8YIgwuan0XtVm9feEBylP02nysKp8DIaIskqC0vPa
/H7mumw22IUN/pUpHRv/5OELpsTppiukzy/dr02Zv4ulsKpd84NL1+COiKYygKn9
94EeTTWweAWGz0eH1mlztnHrhXj1GBiViYhK8ga89v0M5cL0Fx/iqkZ79vcxPlbD
Acl+R6Gb9CoKfvfSGgmbmeSvPv/8JuEzIqlwBMLczimtfXc2TVhLfHPXg+o9OBPe
ZC7VeLbi3HxB3FyZyg51JiV7AaM8Yr5pzL7jao8yYp2LUob505yLnSSQhZcpqorj
viLOmiC9DuUZeIy71F6FVAZGPXNVUZnOYJQzipEinvYSQaiATOpEiZRdvqM/aVXm
Ye4sUGZVU3mqS3xrMlHm4MFZDWi860BYv1XYLGEroZr61I+HNhfBala+yVPoHUBg
qDm0lhllDxWzOE5cxfGZ/MWT+wbLhxts4jwoUUx3Te+huDfwPj5EG3yB7jKTHgR+
hn3NtlZGZevDBOPn6DZEE5lKJDJUFmtqXECypQAB1oQiMfNNP0yh6lRLJSE1XiYf
Ge4DFuKBR5GPA05T8gqvK/1NbuvMFchu0LRSrrHNyBTE3PeHgQzcdFOXqHeYcwzM
OpzUZ6G+caxDarKxuHLfC7EGwcZwFQCD1g/XnkuPiOqwOL5pfo/wRTZrnPckbhub
+jsnSSVVKEamdSR/cbN01JzRYmV0cfPwe2L0s0y79AG7EIUG7hFhtOCc5oEX7zcx
`protect end_protected