`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 8624 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/9huKRhRMtvnNqb3Z+UU7TahEoHV+T8U3P3ufru7l1O
3DlgtZzb9QxCbOjthp9+wDkjygH0eUfDrEl1ovhZG626rM6LzNyrxEUSurFkHnfv
UtiEaYTIrN6y5AxkSq/bhD9Vw1UVll8r4/dV0vn15/kz02bjBfM5/QQbGWOv4KM0
MGpb+UeM4MzNwJcndrrSyS6ycpLfYMzH8ETDowrmIAmTeXumW6LDbNGZ8t44YWsP
SOdJ4jaBgXeR+jkkvorc2V/aR15ktChb/JgwNmlGec3poMWfed+F5HwsZMj6fzOK
8PcWbK6WpqQPUyVUlLyRLMOepRuHilm9Z69JWG61Hzeg0YLDNj1nyAIS0Lo7jCKS
92HgXeDWKF4H/YyH6YmWxYYsD48ITyf2Zez+8z5PTATjtPYlgWiEOXLzfVJYdyB0
NmLOEI0VNzwn3tVG2C2C+7ybTFnES5s9CRW+Ji+OAvNYFPThaH+tmEDJmSGqTzZB
k6Ptj2SMh7wYW+dmc6sw9gyXMn2X0JrHi06S2+g3dkJsiWmHzMFF8qQpwgNnoqmR
nyHCBQ+pPov7OBeJtOZv8FO0b3v1YgqiSM5NuspiSKpMCxof/3G9gpdKvnWazeJS
u6eMsAuedEnGSc52kC/J+l3FEtA9pgTxil2w00cEroyN5tGrULe3HLtmaIkjIoos
K7GCPWjEvXOJxW+OnPvPZrXf4SCYKo5XCsHbfksjGM6qcy7PI5R09yMcLAk+CTR4
eNtQmUDeO9l1nJB6Ms/NaXFq8LqNs06uB4ZQP5WfPMsrLdVP59HSrKwmgJwYt4u9
dhBu+9+aU0ky2c5CDFOfP9t/aITUaBpkRea7DXCIGsQeWYuLhgTPFAAfo4QIwyK2
TUSdw0lpCIJZ9LV9TzvFiGIoEKaEiA1jANt8R2A6RjvzjtQ/oiSxJ+hr2PzNzrQ2
O4xkMDJAHILocqfeqoIJytbottSAAWZW6tT1R/ppFcN3SqoKsBzcqGRtssHb6uV/
KCKH33ZKdtdbVuARhwQcBPEJTQjpnIWqwF0gKyQi0guFuqJSkNycs3wcgpOIEjM8
IuF7VYTtnMybt4Wvwo9zcaTfw2bUyQZgSf6+UcMZ4vmfplo+NH6qP01OUkmlt1ya
h1XoXabYjnKHuh6e/m3jjCapIQbF79Fop9ujBjrmmbD5W25apXtULHLXzHv82qUT
9UxSJp+WznaitV9IXcfxhi1MZs14I/liSW9MC48gUiZmmQU87s1OhUMgL6Gy8KvQ
UlqEnqa3QRVUwWNArl6t/k5pBRof7+ll+XsmswEIIGZNAZBh+0xu8jxSoBwVJbgS
8MrCH/LUwKYarLzUdpxuMIWBcwtlOkOgkHv4YrhvaT5AiltaVBRKE0XcBIiOcPF0
69Nq1AUakNw5+E/8fD6+9h5asbBCVuNTPXUljInnerTh/gv4mFVbrFBq3EbMV6LO
H50Q3uBj6eVzP+SbaD5cyi2ofZHkX0C5eza0P8ygj6vOOwDGN/YS4JleaYDX0Ig7
PUed53mwqZ5DjxQFSBMB7/Q8/18Both7YZfUzNViHidv1HEJNuIFLxVHh7i2555g
ULzWVLQZSJbH1NqGUmVr07mgOfO2257eg+UQwLATJ+8ZwEjtb3AGoI+DkYR6l7vw
pwjc2W2HwO9Ryv4atLvlwstUQBJFuaXnzy3vYFqhAbQA7D5EtPwNMH4H3UeGjFFP
Sr3nlx0jlH3/YE3SruFCGWGavXmOGj2d3Bfwd4TfOFkclfwIP/96DzsnXoKcCQk2
/bx2ayFtjhBjrSGefjf0EBReEaLDz5P4To1LwFPP0s+Ttmq0HC3mCy/PRh6Lt4Mo
nNEqP/6TMrJgC1LmRj54KCPq2UZUp9054PwgPFx0jw42TzBB82phbcsrsZW3JZwX
NIYojGmTvl05YbGGcbOoImgFSihjfvFYLRpy8S4Vclrn2SngXbLDzAipVY5iW0x6
C1w6mJzrEzNjZY5ndegVupS+ULyTVqa9kmh45+m/e/zdpDEY7MDO1w1r9p5OQR6p
HczzEPcD/M+xS6Q8BkcxpD+YZCbUGFfWcKcbd2n5gjT3TI7FVImVmRMCU5PIfQzI
rUbWRuA71g6JWudulmY1BD7uikgauvAhwMyk8lqK3qXJCqKdW6R01sk4NBXZTAJs
VVhT33+0xJh9fJPPZFppjM0NFVTIUtc2NcMKB6NjvdvVoGiS3s1hVQAHhcHXXwUk
sU1aWsr7Pw5oZlJr6ItuLdXrI6KN3lVaobGZJtdQOe5Oso+q8nvuD91ff7FyEtly
xMvebZ7zP7tA6c/zlGEplPMQsZHc+wUA7yyohEJdsQC0VLl74LLo56H+WimdixiP
NFFckb06pfnjyqoS5DyniPtEkbNtbujW000FCfRCoZnFuzGIc3KnZXcYAW0QtTyC
aaR9dM0mps8dZ1yCyS1+7Tk9jMa//1NXzMD1dNI5Clw7nVC9opmQVsSJV2wDD8ra
rcxTHW5b42CHzgB9Tp/FKIUs0qwB4Bjmnnq1MtKHTZnMKzDZ4fDBNOfvAVdTuvgR
4UD2Q+crK/AP3u/GdckhvZUHM3K1DEeqwMLwEqxQwXc2Q9F72cA7y5yUgDByL8t+
qHcHwl0nh74Z05gP7a5QY9VAkMcAcztUrCpLYTjNC0Fb/R96YpsYvTzYoyAicXb8
V9UI8ROeFr0xGPN+lo37NwIXjqKEY7Hn58qnZvaeHgP9jFZGW0F1oN0ZvwvediZU
Q+GYQkpRu4kKgeLxU/iDCoYln+iMY6eCvW4SGrxoDOEcAMQ+qmxr5GOiTb+qd6UX
9pNOwWUooPSOHhNwmcPPUwtq4Zh3bkrTWNtXkfXICwdxqf2WqvIIJYt3vsMhTJMa
L3psMWEtnPCf8k9ZaTZEP0cDd71Z7q0z02ZmKD2W4LvuypTMZNlj9Rz85lYbuBRz
16LPfrPXWcGDdnr75EoAOBq836o81qL176/GXzos5SJ6dcfn9uJ3ms4W1BlNG58E
V3NgUWfNRGqHj8bnQ3TChwgkxziHN0RdP0H6DhdJGFdeHqlOA6cJS10i3rXNjYJk
Nx5YkeytTTccuQCUMmvJwXE5XNy+Qohy/SjQ1dsasnUCBUwtUwczLXMII7EF6XI0
sEaPsMMEqpWZk6ptzaMhdBqbs3KPYjQ37lP9lVacgB10GUp6Kq7qOdKqWL5J4QPW
KedjBE+4+MdkfCb/GtjdQRXvdZCUtjQva0jaKCqvEeU6/FqqClXs2REtKzJV77aM
lgGHUjHblj+ofVCkF3Zci3FSmNBzwXxJ9HOTKqSybL8YgfVtf5gp0KA4m0I291W6
cdSI07q5YdzBqTh5pYrMDnHaHenNc0lubYD9b9UJbYePlZPogcQf/Ux9QGv+7LT+
hjD8JhX6WT+Z52cLbzXxrmHekpCkJORMgmf6ysgdNulG1zwvmwb/m2JC9fOC2vot
c2J7jzyZ5w2UFuUhYFypWfYo2Dp+DstYDacDHXkKtPUuO3wD6z28fxgxgHSUygKR
NMYREp1FejIxuyqqKN8ewEmkSDOgiEdxvh1ZmrXRk2cpKyRZ2UBs3oYE1sEgUHLB
mBpQV7/vSOS6Grk4AR1RaaBOa45FRSl5vj990eshFIolwFhWuobWbvg6a3wYA4Hi
pXktLbu3W2LXWWtRSVncgCbqZpQXbOtn1YJIQaOGG2ML60KjlPVpNyDOR4eSQRAa
wI3ZyMOMC/WB/ZEAwgPjCzCrpAuSq35SJ8QQ68bxgAd8hw5z91AbnWaK+27WLYiD
4f73g89ZcONKtljkYwE951s0pIoUvx1zmuPsl0dYFuaoeXJ2VdKNtxjimqfAAZ4A
MfWsUyoi4sX12Imk4WHQc8y8E+CDltRmxmYON/q4LzzqEMGI2YObDwaX8auYb+sj
5des2hWiMuiFAo5F5u87RrZ/g6D4MibrPBU56YB7ryQo3j+bZvnrKGgBDCLWleW9
XeRRv/j/VKRSnqTS/xOUDU1XWPiXNjFD+WN2fU4mtMwsgILnmVu+pFMB+0GDQqdi
D+ZDH6copaU+YpoUe97/oXo96+3+K+EJN772HjHYeIehIgyvQ2z45gtvysWcuWM0
PtX9BInD4Kr+bXR2nhEM6+ikX8Pbth4QvhhGMObrgZnT3C0znAOyRYANBTIDAhn6
KXpTpBEP/zhTs/H/4n2AU11j/1OcjTojI9O/0K9RXfxkZVhzlKHwMobUza8bHfPm
a1EJcGydE5mlSbCWdpscc6AZKRpRbyiCoZaxRXkKKl4CX3Md+Vd2/5+VO5IfiIa6
4ZJEC418BoJvHcPwcZbhOJPd5r8XligfIHLgjShL1rvEGC4E83cGNuGyba1/pwmK
IAzbnXpr6UZtDkNTJRa6rW2YxQ6p7BBaHbUYW/lSKAArcgTcS5KNOWsqtX5CF4hO
vaF7guOlhEu1qWRspsSBmbFScGtjFpe0tbe0AwEwh1/oyl9YVpQN6P/ZzdZ4jG99
HIhKMnS+jlCh/aJmvJ65GNKMzxx6CSa3mLJIQw/l+/FUBk/X5kxM/lT/JlzJ3Fgr
AXhmNdUrATVAxxH+qSyPmVP5qM/qBZZ8cIym92XtLk56LMFPOC1MKIXNjZcr7+XV
7d+sXkRZTMEZa02kJ07Xmmp69TmPUmJHZOWmfuJ5QJC8FeqJcCfSn17XwpQmPWAB
2W107QR8WyuXgMfAwpLxoP5UTHPeb/5xZSMBnud5VXajoSHBA6Ri3v9xglxvp9fk
tObxkO/K/db3OBTQlbpf5OqwYF637s7jMtfgMX1yXcj5StbatnPb+hjHIBU13Gyj
nMfa5cbOJZ9w0F9KEQn0/r/pTQsvHtZ/RIfTM+3ja11tYLa2q2jCPTEBzHgq3FSF
5pQ62yzsrzSNZbzXrutvVtnNYQrqrr2/6t3jQKKMB1Miib04HnSr6pNRtTzoSMQe
QJLfNOHzVrINBnuyjpREaSfFihE+/+73VdJLlawWPgat2Zgs95TsV3Qp9JIDFmWJ
Scx5rvRtxMvvW901Z96zBCpCpJScJvbNrG2a/8uuy43omi4WOwuAoolvxrFUCwy8
YSFfUgsUWwkMONy7GJOPETSPvcnCtlMB3P3zW6TPyHoJGmVGcQRLsCsyPnPxp3Zv
gYFwkPzQ9BTfVRoK7yQVRzo2HfecOWKucbDC7oKmJ4WrTi19H8BWqPHhopf6vKaD
dYjCCggNCuA++/cQoVtXDZeb+SLnjKwCKs1HeCdNuKsju6n3YuID7MPKb7na7XbL
T9SN2Pf6nDLrgNl0sSlbXJd2Ofum2q2+sO93iwma+bds/timlSMi4FTZDujCGy6G
AtbIRBRhZ+7kDI03v7FasztQu/+iFXvHweYR2cO6DllTW1Lqu0gvOIrp77yGh4qz
LMfFVkxR16GR6LiCPs6wZQvYv4qwxweH2ehI7BTNHtHejVB68ykzbA5hNqCOg0cK
RF0W2fxt9RPz/SOvLZ/RqzFRcx4u/vOOJjBFp332N+CrfnjnC7QeObAemRs8VIae
9cDcjIp7oJPqc36PcFG2dTicowaY/JVCuCtLn6HYc6aXc6A8enWrscmoYfdKF/xx
smeCgt7Xd4asdZqoqZg2evpX2/cLea4gYDeKMuNdqONgS7MBVblqpcesd8cW3KX5
lN1eBzuvwnUz6Qd+fDtPKzBREXfDL7m5N+BXwQmEhskXG152xEfsuw4F7AoDPgQp
jJKLJEKoBUMXcfY5dPHyCHzgy2CqDrdVpbzXZRdOxyraV3nXHff3TWKjWIyasDkS
Brm2JbotDepIRgGdMvP1+BhAyF080TO7QoUMqUdQNE0BaF4xzSBWYzfXN7iDwFQz
bbEghCv5kOl8w5CPC93vfByNxqNCG1WsXZWbOPmHXe2SPzmDQp47FkZ1lsl0gyoT
fuP9wesNpDIsj7SBawNUmWJgWDm5J+6DgOuWVEK9tD/1g6jqm6uk6uPk6CHWzNLw
7aVQ/dhMpqzt6fQB/E3DOf6rpp+iZJGHaYMCNlL9mktljERBf0iipKJ5D9kerjLD
zsY1/mDqqkCQ/QTtf6KU2wK+Bq9QparGIXWwldk/k0jv5ioexefxG/Bz4ez6p80O
BG5qNCFflhHgsopYwkn3HX5Jf5xph/vqThR0UxFZyh4+ypzyQjG9nj7+GCfYKWV7
TUk2veNeIipCI/t6gyPozrLCI/R+Z0JI47vQjl3z4XS0t8u9Vms40WIQMue7h42Z
cl9DiRzv7F1Lm9MpOeo3lQQ6S6EqHjyABSgiXDM5mA/EdzkxhPzBuh3SbOiPBL1b
dTFRjSLorM3Gayp2YAekZGBlzKCbxKTMOCj1aAtCJuYodfEk8lo3TEU+ShRtOH/T
1l6XanlwTQonogC0y8zh2zZsiPVOQueUvsB5iM3tujx7cWkf44Qobl2eD4VBIUue
SjyYQSTyVUWllWWKvQdEOMQ+4zUDTG6T860CBMD3lHv9crI5fSVKDSzee/GJ/GQF
S14HgRCa4x/069Tdyw/fPPjd8QbBwksU29LRo0eg6bM2nIYoLexDYcNGLUtiFAKT
IqBZ81DXtJaEBtkXa8tAgysMqcwjPbITu1uy0zaAf1EBvjPNaIFfY3Irr6/K2VvF
DCAIWWiCYv8X/8C5+Jcrga/uchyae8IQyJv97B2zHc91RS2Dzy5YFO2UGbOSW6wu
OgyWlOOEFatrmYyvD0mcO2bkGtnSz4dJ4IMHzP4yqG7poees+rpuF7XXOO2QPK6M
HMRFlo4fp7Xns0eEwleP43w0Wj4Up4Sec3iwz5i8KPmvI7QV/bIkLF1pri+Dl7DR
1seTbbUDHTurv93zOFgSO3w7znejWWJJVEklQhZJR27SHatTsJHqXi8ibzuXLH+R
DeJdnvFDvSHN/M+J0VPXOqJiIOzcfyFEOjyoLiuHFx0prNSOLSww2tpZIuC5fBPR
ep24rFNx8rdierbgXOkvIPQ3Tm+hlw1bxUDknRum14p4EauQvY4lKcBOvCAlbxzh
u+3tCMipU+GYx497AeVr/gkBrWNRgOiAZpNVKj19bHEGM3hUn1vz4lmOKEr0qS7U
R/TylEB6kBQe5NMp11qjvwQMsuJYvw2BK1LlWmxCBvoboo8R3d0QAeDt/2qcdZPv
L4IqYRXnbLBiQTa7kxHkKsEmFFMIXF6v8y6ZlR4SdnBNDR5FIvqh//knoctVFvqu
C1pdMaXtFA+aQJgpBTDF0XPr8FtHKTHzKW8o9WTEN2ziqdec7hOk+9Zb7iq2dtnw
EiaLDWhaSB+IxGuMHuJxc1ch+pxkb52xqzM//XXkZAJk9osMxDPLoQD/w1pkN079
CpxEvxDE9KFPfk1pZhnX1YgjI2d9EqfBzFehGT2yPMEjGAr7NQUqtUa4JuCLDkw0
FJKYqjYYdBPXhRIGrWpdjWmjtcSHZqaJh4QvcLLqTqoonP4rpmuR5qv+9fTGGuCB
K1mMuV4kNN91M9wABRgR8II6sgV3pSbNwEGnS1oSDivq0l+9WCV9h29IpoDQEme9
c/mO/6za7bx4Pid2V80+8Z8n8vwD8fyxuXYPLfgadyBmaLX9yZjbgzhLY/w+IK16
0qFVeCNGdOKqRHCVanoBW7R3vzEWpj4BKGjlGX1AVwL/1RqX7yW9vzduAIBH3Be1
Natg/Vfjrb0a/xf24OraJkt7PxtBfJIuKh03UeVJrG2iq0p4x6ZtNPHvKXvRbBFD
+VtnMKnrw43D97DKnrP++zW1Z0FYzKGmYjACsvdv9zTew5bA3+DvjtRdV/F5Byf8
hCYMtcxcBkdkhrm4E+A4dY6cuSFqukx2eZH0lTf2kyldlT5A6oTXzmw7kt/LNqoI
C4Gtr44ahrz6RB5eGzwY5wrwKRyndl73vWhlFuIRH4NCOO6HwC2NcrNzyjRfHVwb
KmgpEqpdwW0W110t6ozOSkxm7B48nhh6mbBf2d3fSCmdzSCW3SZJXdY+l2Gr22oV
g07FTzmZrreykyW67k0yyHaWbNxmooEkN6wjjT+77IUA8kE0U3vtplVEekC0ra0p
bPjkBqtVw9JWvCmlCneILfTwQBguzItLz590cXx8WcJ9xDm7pseg29WaZ+y0/ZYO
GIV+alE/spwNtToGkcsy8qAvYNOoT/Q8lUPz5pqJPWhzhiJ6+CAScq9DbNISq2dJ
XrNsaX2uPwJymQHh3HTtXvtJAykqOvHnV4QXgBy6c5f9qpy1N0KKM/4INKydwBiU
gV/N/u2r6IwJig7hS26h3215koxn2+5YvG4uUVoG1+IxCM5dVMhbzN4tDllQLFke
Edu5OP9xnu3uCwS0jYeObRTF4HMPwfE+WHX7hdT7n9bJARR/idzohCOx479G/OGV
4actP6OH/Kjlf8KyLl/9R76TqR8HZBfbvCo7WhW8JforS2ZIOcvN9ewDKFei4NWo
kMoSB7anV1wkcnM0Tz9sv6+uZKwTpOHgzL7zVnf/3eR63Ljpzcjfb2SZhPfi8rLq
abECStYyYI3eoTMW2kzVXfo05npMXNjHSrop+y282AvxWZAeMjoc4OZ5bViwWisQ
+9p5qJknBWsVtg+//uKqFAR3QTyfpaPG9amRBaaTV1xlDkbLLGMmuvGemeZ3fwQN
6dt1pFLBSEOS3DgnfNvIKhneSqAPuPjyBsiJ3ossljxeTf/70E9d3b/mvzNJRRM6
QrcOSqbNd1FM/Rq99NBIgdwBGcQ0o+8Y3O2pjgztMUwfjzPBn1MMXHdxsXadG2Zx
05hrIir94Z2D9bsgfuT0XuKxKufp5nKw4TRvYhoJjztD4jVpzndBHEAJKVlntcNf
/aXLZBAJizWPjfs2sLenMKrJRTgqT+AFrNceMmkGZqC5s63Zuy7zheBE+4b6SysP
nAFB9jPFL3Oor+vRBzU9qtUvD+S6p4457N7TLWLrIUo7PdDjbcDjxXJMXJ1pSSPC
n8iQ0Nb5wRQZlKj9IdkNArWop7Remg/B5kkjKiCwOWhF5uDpTjS+cE8GMqLC+Ier
tvZlMvGhrRZwBMiq/4MVTNT345aH77jQRsPsGIZap3tTvDnUDXyRBGdE53kz7VAv
xvcU3efqPY73i6b9OQSu1G1MWDsdBiRed77Mf1H/V9ru71yQBm+iPxNKm6RYywZb
ggQlH2do0+ZDVLJfcLJvfNhIoBurbMbOoY8BpMtfWB0tQgF8vA3Jje3l2x2G+eme
H9JBBP1qdug9yXmHHFfzoRXpl/MfrmJdgAQ8KEo57CML+cE5FMcaNlpYIBt7VaD9
QVaQ6GGBk2En9gj+ps34VIWc3njM8W9NZc5VYzhasT/QbFRTs8jkA7Qzfm20xTZ3
2Z61rw7M6N4laH1fvxUtRPmniy21FnVE+tPt8ew0MGBIT8HOZ7JXhQTmaBHOQ5cn
apyKGPm6erCXgbpB+/iSBAdxdUrvEMFiW0Yf0q/TMxEXNNiOjBZKDLZOBxqOk5c/
HlRSWhr2P43AybRVDKRCKqwjJ/4iPcBixCvtkoDfCFGBjRhZ1hHIrJl7LsAjeq9a
tanVdPSicK8iOhHOgJd36wpM612Ab3dDRwe80CQcCEuiWsOjS3/Uq5Mi/aR/4c3v
ZKf8fZiuP5CIipp7WZmbBY5HFXs9QYSZMbNs5iPaleMjFHUbXlkvUthzzRSkZSdF
ogB3vOnLbvp2X5aOfDlWMe7fWHBAYqvumL1GynO3ogT/OITOvQK3fRinskytiOdy
V/w2yxUYzwGfC5OjG3O3yINDr1KPyX2c11BWkzZv6TVzOSAdTVrIjJ8hIFjiRku4
+s+oOHWK6e5UrwegshYgplJuV7sDXSd6ceDW+GyCGvU3nYn9FU+YSIto8cy5ihJO
2omQGc1rAwDi47xk74rBK82/gH47rPEpT9QR/W/oseaF9854msy168O0svh4Wuqh
eSCSsVT8FRJJqaYrCqQk6rn5ry/mTxDQ7CeGAibthcjl6TXcfpGkDhI7Os/gl4Hw
m1IeHDs7qfSnTISAGcEt2sM477OkNiQW5WNB+DCNGwbtYAFM6fzVFnCImvRAqk6n
Mdk5YDoqMnWQ0svnJOpG2Y70gmJ4Rnnr/SXTUoddWE5nru4hbLJNyPXu8IxK5c/H
QAKPKSOeydeAbG4U7lwQYO2ESEjMM9oDop2jUV9STPkACpwQxSrPu10kguTqOvI2
IE1cOrZLMQxF+QfmdYxQLaQRRpNzvmDuR9MSl4crVxEbZWo1weiKBswsPOJAufwA
Onyh88uyKDhCYfAd1c0lY97aeqgMneB6siIVgmTVgiBnAK8AosH5baFPcwKuNrEX
Z1dEXxtSsyqput6krOnJ55CHki3NUDBcl7VaqdsBxSK3v5hapvLyDvVA9uJAT4dR
RcLVB9eL4iSPzmQAtGnjlJOz27MPhF3hpFKhP2i0VtFLn5v8Wp6lGfjt7SayvDwM
0v29etHcDWfjD9Trs73/Wnp5DoG4LMYLWr17elisC7ywx/9ymttYEIAzqlp7ghYl
n8AJ33Vcp8XTqcFI44ivgwCLNAfah9+j7pCy1qRvqcfdFeQKURk4xcUyHlFZfbJy
F+PaB6NS3F2BgYpYgwWLczxJ1RNgR4QldTdwmsottGUd4KO/6ZZRB7ejG7Qf/EFf
BMfidnNQ8oSlJ8MQbmRWWFTdYL6rqEMCjFTXdjSiHc9/HUL5KOJ/CSnDGi1wcnu2
6/iUfw6F8iWqTWY3IJiY9oCNsemUNAKO/bMb0du+8eu/j6DcVu6SfmMNnkI3aB+m
TpduPcIZglvrbBmfOPAU0M+xaj+v7qDDkN+62Mz2YyDlapvKIWRZhjL+IZbnyz6t
vVo6GFqP80h0I3415mrX+xCMg4RWkyHfuL8BxjTaatEwtWW/33tAXs84qJQD0YWA
D0aaS+T6K37B+sipD4oeKKxf3nRGOxubMaxHWefZ1Yn9uswKb7504ISTVuy8MDD5
1JQ1gQJ9BugTNAsEQAoUe4KmEyG1ZwvYG7vRbMc8FpPQLGsggB3BnTpakj5PmiBR
FNKqCqlOWMLwjqYpz0PCXLcOJUNxxuP+hiUDeKKzamJy8UaJglnIzASNeh0l8Pe4
L0wQwCilO1jJUUpxnKl4IVsiwSsqNVH+c3fKwq2ygGyjYrc4R6zq33Ob8HXCxc87
piQJWixAtZzRgxr9e1c5Db+zvNDiROHVbCwj07qfgCZKYPAksYMTwoGwfvw10gCk
kn1hGstiMsn6qvL56AAh+sIFnJ+rQDzccn52Y1STZ5GBQ2dtis7UoBHU969aNAjJ
UcaKi395dfGLlLIG3tl0huDCEV4QKh+/Ps+wjT3p4FaLKPv3ClItAObsu51sRoui
1bqfCrC+Wu5a0JwHWonFpPr5JJ/0TeSEZOmdIyx36yjm0huEg0js9IcRdBVbR6qJ
8nmodlbDPbiz77NnczneqM49Aq/2Olqaijq6i/1xwNTohe8N1wuQZLtMPja6sT/N
1c0scHSCQCzf4hyEnvKuMxUOBrmSXXfhN80fKL2sjhBStaKb39LqqUVVo70s+YcH
DUDHDlGuG/C4w7pL+EMaZAA3EKrMATl6zz7v2Dspk10=
`protect end_protected