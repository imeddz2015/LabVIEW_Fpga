`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 2720 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/9huKRhRMtvnNqb3Z+UU7TahEoHV+T8U3P3ufru7l1O
3DlgtZzb9QxCbOjthp9+wDkjygH0eUfDrEl1ovhZG62av93pcepPPCqWC/8qqkfa
BfZckDVSCQgHCoKai4JL3NL0eJESqwMNOBHTks0j7xloFBpTNj9dozjUYqSsrOa1
ugo9f7TmP48EmYJDOKqtwEW+0bpE4r6uYe6vqOqeYeSbryry7tyGFGJ/ix8tE7E0
RV1VO7bKt0f0iNaNDTu8ZAfFiIRwQc0SVPcEv1iLsa3PNafSADQLDYqTCYhNC+F7
JsiBA4K6jUnCIMF0etOdPDuVz1hWVBr9rnZkeIQPU/dSn9ZadHiux0aweVBEAScE
gawGnDCL8dj+mojY6HV1ceDrpwAfQDgSqwPQS3Ac2PpFP7KaKk82TSp6kwq/YFdb
mvrF+rk+4tBIBzGI05gCu2Fh/F0UwUuEF9BBUw3KKNPEHPM0EFDyjCr2BdkxpO6U
mOqqCEQAW0wBH8oiO8R+uTxvCrNV8K9NN4nJ/hwUhLKqVe/lNiXx93ERlnH/L57G
cHnQjh86B8bvulgIx6/6PQVuqLfnPyaTcH4UWNpxP1/ssgIcnOts9Cltmoyh6aqw
iDSaLZEAwD+oB9WU/RG3lLd9Hc0GPkLakdrJ0C+/LlcaObU4Iehx2npNlWrggFTN
9uERwlGzPjWwFEJ3TDxiT4ttOZUuOGF06wK711Um8qUdlk6YaG+xFaGmmNNUptDm
qmO8OTsXfu6+Mrb697MhxKJDlvrvFWcWEMhZ1XP4ubFWrMN7GH3xNAaCpABWCycx
+76WNnKdP2Y1UJL0JHinQlwnuo7Ji4/RENZst1vLvKzo9kD8sHgJj9QJPWO3GCNi
fOKagtoN+umT/N+0APQdN1kqzN0yNdD9Y2YK4ET3d2liZ20FdpLKumKGa4750bkw
z+FKm6YNizUofqQFqZk/Mfu3AsDRaWAa8PgelRSRUGR2/sNUOZUw5y/2cnWrnoh8
LUPQbJJgNwXYOI65MaB7j2PkEFrmrhwi/gu4kvAeaj9g3e/CX4ZWfctCQBVG+9ID
l/PESIUAyV2OsAkJyigEGzAIIIo0RAj2aGcCwnQBjvHcveP/45XDGq2aJIeCB8HZ
TGiNhh4VFv8tkgcx45VcGuZo8H1sN1V37CqJEujwv+wa6ddvevfP9pZljxAzmkG3
cO4ZyePMdV9UZEZ4O7NdHLNQCIE2q5ZnabyhZrOUPnN2Wcy1pnSTM0czcVCqmjiz
GWTieqR2zBFnNUZ/M+xyvNPH8iMeVOWo//5QvemqN7qYDe3YjOHM6ShNrD8DWJuQ
Zu9TVLxNbp3tbiD1RnMzer3rPRignSuHjFpB3lA+e6GY70KJe7q8VXYLzuFi2ZzQ
DyCbQ3yTf4T/TUuwcqc3Nw1Jotfn51eAmtN5Y/vCQ8xatbEbcns9/CReW9xhcLtm
D06QF6xDK5f/oQujC8jNihxV+lq92B7MfQ32g8+l95HlKMgVhFoDQuwrsjoBWw56
BiT4AbhO0v5R7Bh3wXLYFLsWV14cWL2vOdqATVq+n22T0c6w/LQs9a2An1sPNRo5
tHYvuAc5Upvq9Op2LiJLx1m+tgwvzJCCgCRpnlqUJRc081zlIHHs6yh7Vv5e73sW
15PQ3pHyFXcxz5lzO04IdWMotQ96Gg9OWM93GU/bjnx/RRi1WgIoK3GYr8rdCJCY
qP1wSv509HBnwNHdxsS36xahhpdsXxbhqNcm+qTMeDhSH/7ToN0v53QwWVFHUiQp
3GdWHRObHWcutCcb/+xrEez22jtMa4/16zi2m/pKtiswTx/6rYVlzZ5ky3Jh7HnX
X32kVme4qeH1mtRomDCRO8/9i131Quj/KOsohDVU12KQPrWGX/Ym2gCg9+u3BWVX
bdgDo2WVmftZ2c5Qlebb6r1lRS2xF2kqAUkMtezMzv+YiFFxJJovYHz6MZEpECms
wJNpUKhhOFS1mI+xA/vkYQL31Qx+Itj63Plu/ZwImVwioL6cEcB5JomZ0SdmlB60
iPhC+ssbKaBw/bBoIpjVXsWEOq5oPum9Z79j+EMIyfA0b5Ps6S5zrC6eG7Jm167Q
l+sbAxsQY022SYObVxwcPD8FXrFVOalo4ejxMtor6MutyeF4wXKpQanwq084Yk0A
2CfycD+UgGbH8crVeFLqcWyp3dKQJAN3sz67KtuUgAHZoChWmy+PHSObiQ3iDQqu
TxeOyVfOMsEvhndx8IKtLFnPeWtTVD/UAkrGtGirb6/zrllSF5NWMupIMC/6qZyo
bPrGqWvWWb8bXw3Y8EDqa1D7f5b91NVBti57RQOMlB+a/X8FsLwoosMDskV5KeN9
gfxv9Ho6zEB29R+5f4NcuJbOvNw39erOoX0KLaYc4ylh7QilHRj+nnNo2C5SLn0t
2sxFdg0r2x4P2BpsY1GY4CDw8Zp7tQtic3SjNYy1/3EDuCMuEsx8z1tIg00y2vXC
8+EI84MC53x7A6x7nx4YN3JIgXiH+QsrJuDyE1pzMAKYwBxQd2IvjJSrnfMn0eYZ
6GAU2Dv13MaXPHsnGvFg+HR9jlgQMcHWWyh4MMkI4KRnuD97YuXny5FRX7QJ8TY5
yla1k3axW1Z5QXJVq5UUpLRUeptjuxOHbsI74iWkwEZX6RnW6DdyFgIRelqcD/ap
7efFpeGfWvdkNWBaYrOo1Ylsfy/LqwRxFFTMr3P+94ttdiOtANEAP7VS9uBFPUJV
DjeDyXoX25ibhNMWcE1qef6oG3X4heTj0KJHuU7/6KX6hDTVmrVP8ezQ5ou8s6tu
kNnOXCXv0yvToyqRs1q/9CQx0eoRP/L15VcRKra+2cIdKkSHVvuqmNRY9myotbjw
zRyrrYNKGyxr2gz4p0DExLZyw3L8MhfoLZy1lRtwMNPuTyaxNdIXbBMDd9aMUx/z
vxTIqhKxPfhVSeyWQPpp54Oa3ApvWD84EhA6hDIfXw6dQe1wQSE82y+7ELgKeWyo
r7lOk56g75ZNe4EGvgBf4SM1nxR58sODsYNFdAfCs43oXXwB9rhhD/zYrm8YhhIs
38xRxSaiog2C2hM5z0YOsJ3AQ63pbHtxxNRgD84c30yL6lvRQceZ4tfIbjcGtq4k
/MjwXj8qhYK7siQ0+StfgVbpWU7HM11ch6HyuHOyA36Im7+PUXAOqPskLPa+AAs3
oJr/0R/1XwvN2ahx7KDxWrXdCRxsFhK2xU2iRDmsMOoWt9Xm51I+Ty/hwZMgcudD
Gem5+UZ00pviGJvqcgzs/gNw4jg3rLYJy+GRD8odnEZ5Gi9E6YRXUGfgSclTwttL
S/zd+7n3qfIay1w02YV/jzQ9Wu2VfI7lb1qJoCzY0ExQQtrK8tO+VLeiuYYWyMEh
t5SIYDnCnL8PDoVhmRdW8yKZU1TUeqDGQFTT5O6/jqh4EtgNrk9bQVPmxTOv+Kbn
EFf85eq92BKkOh5nLzRSCODVeZIH8rbH4oX49c8vKJaQgi9D6AoqMKmYN4wVIN8m
FJe+L2n0VdQOax7LB0MiwYxuZUIXB+kZ9jTyUQfqsUyJrNwvrRAoMnAIF9oDq7Wb
Z8ZH3MT1S/I6HVtB4/2fm/fOlgnY0yzB6osHCP2GGhs=
`protect end_protected