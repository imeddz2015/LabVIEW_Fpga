`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 2960 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/9huKRhRMtvnNqb3Z+UU7TahEoHV+T8U3P3ufru7l1O
3DlgtZzb9QxCbOjthp9+wDkjygH0eUfDrEl1ovhZG60CPbBRqQFr1Ma9nzGwOTqJ
4wLl/cNm2XmLE/y/1MZHMHN7HagEGZPdhIOEL2kgtPBOuvvir70j+o2MlDhamAGv
L3OQBGe/NcwYR81OX/oNH5ydrpBvx59anE88EeyTSS7ijPBbsgteFpA7L0GFLUHn
JHClcWEQSNoD9cseX/6E0REuTKUVT3W29tQnC+UkW2fG9iw3+OTlrhzlKLE5dncb
j6ooyIBWpbXD5LAychl1E9kncIC4aPuuyWKMrHcxKU/VNW3aCnocUDxv4Zn15HBL
/WnWGZB5ZihrS7IxOyA6smkVWb4xT5bJucTlN2rtD1vbv07Ljy0qGLbGlTsplosW
QvGTe2uSaxIWI2ID2Qd414Ot6ZwRXbtfu6Z5fjUcr2sfoKqMwIXVqEZYYysh5TQa
IfaEOL+xQ/PpfEtTv5gSXXfRAQuxV0TaAYf2a1hvBLZ5Iw5dITqstzjssmPIwPn6
8GOPSZhkd7jxDLTQQ6gUIsRildfXAKAFtBcTNySbMz7Ibwee8sIhf9wAq5TkkKWk
NUzPqM0ktwUUC+NVGyBG6UDeTgljnYl3TBLwXM5nlMG7VW/EVFGA7/gWjcSxst7F
ieowLARrD9ucZPTDpLczDxIAmYQj3RrYX3XBuZhoi7Brh+e3OX0CX1d+j9RzZNmd
XVm9hn5fFKUG3M9HclyP9xCyh4L2ycSzcHHLYJffY1E9auOh2tVTv8pC4w+UvTcz
x9IgeMPrExBftbqThHc+nnQOU69zcwkfMszKSgZuSdDvzSMtCA3f85I98tVpr8J4
4YZuP6M4NbWb1SbDnyypvcn55GhAzozhmbNUTa5XfHxiSNdguucIEr4hcf5T/ngw
NWfmAOv1r4WuB13AogR+U5fUJ9aU6Ji2NgWK8mxAKpZnY1lU8L2RS+ekxb+AUQqt
hFGrFfrcIRv1/CV40BFJFL5PAknGn+Htxer3pIpR8BuhwLlMN4Fnvvc5EV69CQPp
OkgjxL6OQx5xi1wIdcvlDfYXKhZYGyeRwniq1mVptuD9hIDWN6hhW6nWzz0J0+Yu
YqG063SM+NfSirlPyPjMu3TAsyPZmH0TdC0a+tJF+KuLGKQQPUt7gR1rycgXXj3U
b1VqGFyP/8VoR14IFgO9L1xDHTr8NLB/fjE9hAFawD4DrcUl48MgAmpopjUBPlwS
UWMnYxTiY7tmyO8kIh+dDE6h1YGEwpxwuoPQwDD7RmsdARmuBfCDaXd5Ziob/YzU
Z1/1tm+vjmlYEvU/yjvDyz9K/bS0gE9Zk8OpyqaOBhrcJ8F7mGDZ1s5cgptbyWKf
vtqF9qwlZ21ICQrUQI+QBGjaMX5cyc70FSXMJxuiwSjUCENHBET3XgHz89VdoT8k
too2KDnEx4noeiN9ektiI8gXT7IdjLLS3X7OdSkY4Cr7+D0ZRbwpv7mSIt+jQvPM
FEngszNucxj2dCn6tpf0kQ3D54POgN/AUHFAL5XZV5LKckrgiFgYQVl+dXy2z5q8
2lQrO+n2XIKUmRtuBhwJLAyn32lQLrf58ESu55aDdSTxXksqwAMn18OjvrVeR0W+
0jkreKI0iF4oxKLSzDaYI95H+GyfW7j2mA8tXM4bpCVRKsQXH+/eIXDAHEbI40Aj
vGNRKTUba4Mqeym88/8CDGDssxEZKc3sPawIxjTDK8JG+Wo1tdMgKgA1d0xl+ctb
hwfoQIGOmsQR/Lqikum4wMxP8e3iDuVdWZAaYLnxDBwSEG6bXcWI7gawUA0JJMj9
2RtoWwvrGUSFScOcFz+2P69hWcDAAKiIeBiSgeWXF/Us+xRFeQjwbcL84nOCoESC
9eA+UrefMaV975Wj5lBbL6IGHr4cNUdj1aw4WGTgJJ8iD3dadh73gkjqjxdx1tYu
A6JF/kwX5aD7KrFtG1Zt382zBbNUiBYzKVVasjO8XJUdkSj3Kv1I7WQgMpthyJvG
3KCx5VsyudbNCc7GAg0JYarWx19IT70gkcN2RQLI71RVolXgTN2WGNEriV2KWggs
LsmIGNsWPjoa/0Jo76gvhcQightd8Zqjs8xO65mTuZ2N1bT2doURBCqeQCP80IL8
uiMzes2nkemxU5DogIPIvIyCC+EMS6HKmECSfYFfU1OVl5c386ztq1VgWkFsIUD2
7DFA7/hDQp+/RFqklbNaKkKuCor/0Dm5uXaQVk1lKuG8JOW/T6aL5nHKssOKPt2e
kC0rXSlMD9E9EHbP+IrK94fBj+b5oEw4tfMxVz45An8yQ126FR/mEXy7yF6mbVFU
84PtB7JKJpu1/qjxg1dA63Gn7dAtEW953HdAoxjS7VDd14FLAqIjHr9+JahSVBkp
+lPHx9a+/0/sZO4asRneBLkovle06B2ne3J50jYUrjGys1i1mQKhafA13UyD6oq+
GEanGcW47gK1bTcMMYHVCe1l6DRqeMQtjONyDaUeEKPMYvzNDPAdW7X30p9iSoqB
nIjXlpxL2n4nE+jCJfY4JxobDj6Miksu0+Wwr+WmOWdkDcuMjF5PnUERwPyEFmfg
SytvojLpZrFbLiyMVb2OwGvaFb0sy3tAiJT5tc51LSgeolTWkfT9suwGQsPsH1zl
nliIpRY8K6XPEUj4Iy2HJyIAA6tmp88CCfvl5CYXpZbsAGNUEfxNNRuvwrev6LV4
ll9gjtyTknpkSCljK4suucOJims7ASh0YHOGuLbfCuK9Q+uWWPl/psardCgjxIl+
0GyoHyR15HOA1Yio71WpdQBLgmpy1xob891PyLvM09NO7pR3bwGb8fu6W7IdK/CS
I51GSPsSbtsERIFeosNsw/hZnIacLIaohlGnKuFZfFDDlQTG6ES+Spx6X+6gaqbA
Jz3rGvExogFY2Yl2afeXVp2eUTpXn6Mb/p2SCH/7/nae6UxrcUwtvvQd/T8tphwJ
/ZavhrhRQVJQ9ubKVv0Yr28feGDgeVllFEHv0eONQ0cK/o41fopZq0raakFppIWg
oCGrFyOMVz6RWonUwOfj2/IBJsDwMvoHWOpUmDSpmN45v38OmecPRfD0mH1rqXjV
us9L3eqYN0IRp7k4R0cW7kBoAa7bPCRHeLMpKUqGXhk7+oQPlez7izZGHjiyZj7e
JRep/Js7EvYO/IR0AvoUG5F4lzQIlVaAMXwW9Zkr8XOFfwpjusQsQY60VkUHPPyH
EMKUomwHzM9hm0JHBPFDUDdRHav/CkcoCLWFDHy1vhDSKoqd3rxlat+tZhucCOVu
gKuftAUiNmj0k1S1CDdC4nyYFlPCoBcM0fT29p3N4TnvNfm8S35FAiRR8RZ64Oge
G+7MBe62xhd2tsucHIbzfvNZIFBkuf0xLrqwU9EyVwJxODHAWgLUtFR4xR5MMDp5
KJ/6ZnmNh3pgB0DZ9B6NkBGPrha3cStQ31LeM3EqUqtOW1X6+UzOU701ENGhMD+g
b6jWqOa4hc2TMamYYA5P9g+iWAleqX9bpvnrESNbx5QbgUeb5305+8raIe28Oo9r
gbjQ06ac1qXERcsOYtV/uxnAR/LEmFhkblI9ayBN1mLt4RyTB4+HtcYjJluEBPat
A77KWsYLlZJPeWSpiEjWiWTLF8l7Amih0RP9P4WjEM0XQQYpg/LEDiFPSd1YTyen
mTz4TrNsH1SBlJG0vmbBVr20zqfoesA8D/DAsiSoSR25G0NqDKD/C2iuXPiBaD8Z
1JNWX+o5RieHzIcac4a6ga0/nF7YcjhrVOKvvB+DwlqM2J9mOwDIhTyhXTuYq1In
U0WecILeAgQiqllgqYdlS8X5w8SFX9lPIct0mqllciEgCIN+NqDVqF7N0brWLcl7
YeANVNqD2e9c3/drpcWZxnLD/P2SUm20Cylytlf/a4k=
`protect end_protected