`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 27424 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/9huKRhRMtvnNqb3Z+UU7TahEoHV+T8U3P3ufru7l1O
3DlgtZzb9QxCbOjthp9+wDkjygH0eUfDrEl1ovhZG611U/QUXHp6s2dmr14S3F1S
VHKDzgpasngQyiRzy5nB777EWNII/n4j3FWdDZlReoVPoDUjCWJ9OpbJLTo3rCIz
vFSjS8352BEJ8c+eQaIrsIzqWlv4jJmoZKZC2y0sMC7L/YW5/4l6vR4VkaQdYK04
aUgOBI8xyEgTjSIS7s7afO40t9bxSmCC21K7rIhbNznimfJrNQ6ycRMZwwP5ojz5
o1mYdmPz2pRPJFbhzmzsSr+RKdfLnOJFxly+qBTcOuoAzoLEKBSod/zzUVBio3kp
LVryk4mkZc5U+0QlLwHQzMGsUqpwUgI3IFSzI/2Lg7dZ/wOBx5PuxIY2adlB5FyT
IsF5iW2t4rV30WXRyP9SD9tToBa3o+3CqsbhLFSVxWa5XDKbHyKXbQmrtJY8sZZY
6FiQ02m2OlJli/rAdJccq7FuY6KASEnAmTZ/pdBbcYtOGdgT/pejMA2JoUZgw2+K
DzVPyTWRhAApTQB9ocSClvauVz6HeGV9epJr/deHNhx5L7dIKH8P4nexq2aTir/Z
rRl12Mbbw2vH1prQbcokxks6D8LLFhG3aBKfSHbjYSfVdQs3rVbkybXqGChC72u6
du52W2NAIrnLOeAs8HhQZiZsv7XkdhrGSx0E+ZWvn0KdC3Ewp+u5IZMj1+bx32oB
SoPxpWmtHmNh4nSQZUONRxY3hRVGpZJaNyi82RwrGWLQFxLLI8p05dbZgCSvBSVJ
WfDPJZPzp0fzHmxS3lCbaHw5YFGIz4aSOyVAjWvygLzEJuLE6nFllcnJkXkxiN8C
wQBjHqLCz05My56iI4PVTCnqU+nfD97IQHAD/7uRPWor3h/AWmR8kfcMvQrTtfo2
uAfcN5Rr7amd93fhnRNLljribgkJJKzuXHRPcNnaeBvmqIfz9j8bptsqxdXuJSKg
tm0jYgh2WDq/jy5sqhbPHaiRrIadJqbz3PhDUx4mALZuLAE284hejsqWNqrXMJTT
8q2B/aMwKxk7ZpZhJ+Lczb9s7OKA97SWWrL/vAN6A5iWieFZRVvOYF7/58N95wka
wOJkx2Y7Qas6nRgwQIUu0RDs2uIVUo8bjaxbqh1Dl3P59xvyrdOzutezCyXzHJhm
oP4lHDJ8tXRRo1dNIA6nMSHBVZYUosXD9GxHQUuC7iTWJPho/G/KBhbglXe0/9Jv
8dQ1hbkZwxvbAb9jZ3cT3HM/N+zf4EjMz84zmORB6mNnWAaI9gQ6BojyJBDyhPgl
7A4PfCHjAkblTMqsOAa43YYc4yj44T+o+MmqSTEjjV4bVY5uiS+eB3jmn7lvbAGj
vwwVV4ENii3jxNBo9n1+NNeU0oLb9x2gVQlfZyNAZ3jKjbCt1CBR0vL0umO5CO8D
o/3BIJ3LZ33TJ9brE5tweWSHSz5Aynf7q2Fyaz63OqNGAymOpAPJnumFmwZcxIvu
OjMxzGaEHheIGqRBUSOTZ0mtwoEyD2aOQTGbfmW1DLcuyHoD4DHx3jHo+SYgmCnU
v18l7I8L6/X6RJvdEMYl8EdWqORyvvbgAc951TzOeqZQqPnRjwX0HOrsywZHN9Pu
dSlnQlsy6sqNqkdud0pp0bsPRJf20Ul5nx13zaseyJnymfbuYDs68Q9a2u4SRMDz
sCFj+BpIcJpJSIqOevHsW+AyDz1QqHZjvzerHKkxsIi70Qp1cOLwtSW2Stf7dpaV
bF1lwYr0goTdsT427zFPDT3FN89yMQL7NzV9pQ/uxq6aUWeXKWuNjDIsCF5Is5VW
KK5cb/2lHldfoo2z8C/7TSUeRWnnwbJ8jMdLPShUqbYbx2j0epWTuAwET/BHAB8x
xyqYckJe9LthAMzuM9c4eUhd2Q6holGiOxUQwA55AGpkZARIw8NRtdzp49DSBJEV
6RKzqgg/Ov/fPkY0+W558Qc+xQ1oBhCLxibchmnLV5FRum4tlb2+wUK1EtcBTOPg
fLR3SGjtDUIRE6HB+h/W6tXVOSZi2a6LSj8tiGJ5jjxlU02tg7DLZ1UQOgDsIuIK
0grkx5F0I7miZcMQPURFHnJzq/hx2bc0VgKFTAu49JAvGFVgiOoxiQwml61MOET2
L1Fu7mZWNan4By1tJ3J23RAbOtVJaKmWGVhkCpcss0p1pxarKasGTRxi2IReiVlp
kKTaxfKTTXArOw43acVevAzMtHreP17QfQV8naD1qCrdt5Q7q4HEaMprK/UkTqei
ih7KnQ4EzFk1sJ+Fn4KIAFBNvU9i63Gba5CLrhiXtAxbC9rj/27Lvt0QSo4CAKJT
TpgvPv1RV6AtIts4IvhEkMuF5BwlZca5B8fFYejUYmCDJKk9sa6IdnhmxWCKPY+g
ybrB+Ro0yF4/X5ZK6Hg+NlmnEjkhRCGTz7N8HPJKvGBgKdQQW8VFYqCAdYE0QCA1
M/kGE758ZPGw6aGfPRQILpm+hSXNearPGyNbftKVpINwSCXd4huS/253OF2Imi4P
/KPdkuwQRKDWJ/WZ3TwkOhmGtwfDwSnOimQBiUAtOrdtDgJO8S+D5Givu+KuOCDt
eWndfphif3zK83xJ0198ynMmIgED+MdLrdgYjF7zZkA7UDSe5G3cTAMlpOxsGn7a
7cHi84uXy7ywlFAwSnHA9/OPrjM4v6B9/Yusesaeq97NZYox8MmKGLbfqlaEGoHs
gZG/eLz3ACz3ezAKe8r3kOX96v5iQT9S5ZntgIVE+Ys3OASzZy2WE1wsBvwK03aL
XR7RfS1p3chhFRolo5WPOGXBU2l7cr/cGkoZkueKqyVEHnXwFceBbVAvN2KYFn6o
KopMKDEASddej/t8aWVQn0Q094nAXopEITaRCgBij1jHw3r6J3coh+UXKRN17DzS
VHrgBe6XTqU0BecAAZ40SMKkGC4kd8vyIgaCYgtfFb2UwdDbREhHqnkKrMEH8yEm
bZ5FmIPsUBjuCuNwbngerWp+6GXQbaUb16myd1CO7x0tmPRXTsC395ayUow5NYpZ
lrEZeRgEaRPrjmoZlxYUUPzeqDxcvJLLt/u75nhsCIh/Z+/yJRCoJu20gFNEAQN7
ByJ/a9uQDNf24fWoVIVcbBrBuHGq7DujGxM9HlP4kQtQGGhoHmUYYVopLXs//ptv
qLdY7EY3piKM/WahYLEFrZ9Izji7beeUQ7mys1CZ/b2yUZTcVg+woHXxl6cAb6aG
k5gqe5JBB6UKCzlVYuElH1tL+mrYVoKWM2/hFqEhx2m7LVFcm3jiclbr/abbFrru
UwmaQp/Qa0aVYY8eR/bN4Gn+OBbL1S3a5PDsu91dOY5AkEpv5a2vxQoocmxK2KO/
UDy/Tq3W9mR819Py5FeTf4HqTRqvZzJKT3saBjCEeAqU3K55X2GorvJtPR6wxoK6
b8eSRv32nCN4HkyYAR2IIJ8gW5ns72RafdDyvQnXNmFlo4eruM23YrcQkUQtRLoO
4zNpJFZG5BeTjmSaiAwFTmBzkYpJkLET8myvqm10M4YwrWo8ycJPYuFKqF2cwf7B
CN0/Xg+iyqTm4W/wgNMMdHH7dYJWRb05b6ro/+sFflBSlI32L+TwLx5Wj+1PNEhT
w+3Rde/+t9c0Xqtdq/fGWSHfOpmVZtCtnlbu2J0PaGHOkHe4ml1tkpLwxrJ6jUIQ
N7xf356Herr2iDD0rEZnABO9W2EyBelz/uBxFwQzEzTsC7nKz7yw6XBUOEyfqNTF
LXA2xbDTFXOLOqkcUH0k2CunWe/LJB2JLdUDs7h4nF04kE96cBx+imxEEnrEwOt6
cfEu/r7GsYJT+DydNH4TgXyyDlmrWpl2W2qENs+X4TMYCP24MfoIpZPPyj8625c2
RO2wKPkVoZuwWRnmgP31uBMDOJbbSA5duOmZKbBxoYVXKUs1Ut9kysL0eu43A6aM
0Xs6zGypd0JoRnpX08Sk3cfUCV4j25TGSeSfyjA0tieG5z3N5SQGKrgZcP0IQKni
dF0lIzwGlFKLWHOZLV4GjUmjhjoRxii6/y4DZczJG0uykv3EeI+4VwXXhgPr2cSN
zr6mOXSSS3QZlszjRovzMK6sQ7mPj/C0cI5cH6s/C3jdOsdM1a//42t9DnlV7/9H
y7vmVe7f77qXeP8/XzTF9ZosGAYSUqLQBKHzsYjOXYWy0TJvge7QyjNvlJmhpNTQ
hV8oE/sNw3XiyouFCeorCy6KY+RapmujJsuEIK9cFSoxgSbB07y8HSkw5Cc3ENsZ
SGg0/01X7pDcvuhNUvaRN/J5WMw4+gDEWmJj8Mp9s6UVU/wa0OZdND196wHVhNVZ
sZXpeZqksukfXdwFvfo2GFRUXpCTd6d9Y+L7dXQmPnJbGRhFCdAx0CjHs7OSvE7L
oLf7lqgv7PMabM7WU2yjAOsU5fji2CrksT9Yd12voZTorQhTZFwjgq3ujXY/I9pG
4UO3CF0snDyNCJSHo674rMdIQt9fmmweRb38H7HG0tQ9A8mjzCe8PsQ5ohXqA4XO
wumrpwNQF54lQcBkflrMoQIGEbau3k7nT94gzkII79uNf/kMAQF2cQwyQ9Qtdz7W
3NCTvAEEGb0YpaNpNbQsjMmPiGAVCqqs8KaOVA6o2gwXqJcfvC8D36L0fakGQM1N
JXT6EInGR+yWAd4HFWLFwa+ln9o/TIqoxt48kJkRhNttuW15BZQ6QllFeiSyGv9t
sciftZLPsSk19F3+O2HmOj3KW8DHSA7uPFUX3WnDIZU02tk4a2a1uQIc+DUdlBeO
X9sM87HKsjCXtnx3dXUlpqESKOvNhgUeXO/JYnJc2C5PmZAfMdRqbCpahklNXG1k
Jk73fPx4IESsLlR16uSSzaCz3hMD0gLGMkAWx6R9mikX0BhsByfYnKXiHnBfNkQO
ULcvBsdDf5bLRp182zxdDdCr/lvtNqfRLWWzgB3oRWk/Y+QnpoNIxhyp4JDOSI9K
oN+0rKI2ajCbOzpT5BQSlXLOD9oZwWfUODn70nMDOdx7Ah4veKK00IolgDoZ/V1i
v4Jik1Tm0Pd7t/wgKNFT2VFyGwd+HlGJSYzGdlVn825JwBOFv8bFeVkLT/1xCojo
RH0mNy+jXFF8i2QC/w3nGiHwSetjJ4nlCgoycfIqobOVp32RaRDMqC2FAi6rFtfF
JJ3jZk9KygL3RPCcVJbp9V4WwDQgInzbLq7/maNxgnR51xpGxicpm3/5SByiEyDY
WxMnqlrDG466HdVDnIfdkU+wOBWGTOBeo+gIPUVPHDd6e5iGqzkDW5PMe0JrKMoZ
EMQnnxxDsk4oOnbhEj+KT8in5Hgf911IiUg+NenDUyrKxO50v5ZO6x9bbfVChZYt
JIz6g0iX3AIKqq5NoAtc640tBwb9/VO8ObCL+jjuh+RTSnkYjf5VfkF+MnlhpWdn
bCPkdtOosFccQlps2+wROGUMPvfStyH8NCmYWC9IQCplzEpsIjpa32RnsQY3tQNZ
/bbfV4kJ9Eittu68s/FnwPt1L0076On3Xbpw/dqG+fgXdXc7luXRLjKs+4aRG7Uj
+6roXswIDF6u5+pj44AFWoX9kf8pF4D+gIbR3K1cc8gXn38K3yWubrJXJ8tnBIn8
iCxmNCIRLF/MPBP7byGefqhrJQ5p5cDVD497SSlgeHRo0dG6T5zJ3VtKGb/tDXT/
MFBP9p/R5NWBS2m7GrDqqH47ZJ4QayYVYono/I4n+Qfx3pU/s18aQHFXXvwr1nxa
3/nzGK7tQ1qjiB78BSOv1pUkWuxjAeJWqPMqS9rHW3/d4zR0X/xUcFmPoWhC6bWx
dyaJY70tFTnautxKBUQzuQxTAzsxfuMoc6+n1tHCs5ZnZRdpger163ZxipdfHzWE
SVUMZksoK8nFS2aRggfV263yeQ/yGDgpFG24bnYXqObEA9Sy09Q1PcFHxJVPlPqj
Bh1pU1NuRYexbMvs7LZMwMQ6Pg95qKV+yO5wbw6hL1xKom3q8uwaT6EU6cODWnCm
ZrgxfO+DwmRf5icCr9asZe7t6sSr7JZPaazafinzVRZLIHobJJ8y2uO9nqd+SN9q
6O7nEsv9FZom45P3n316rHtjiOTUoZ73tPi84xA0gC8FL7PA/3bUapcbCTITxnIu
y2CON/FijvMaVBZO6QlHU0JC1ss2PBHXubQFkprcrcY9ySW+o1JNtj+DCrlSDdZq
1EjKck75hYszUVShhInNZc8RDkRI8bem2dNpb8wW9eUcTFi2MS1R94cxlVp8lAWs
cu0DhZuznAAwSu+A98qo8SVtE5ya+vXc4Ftuvbe3R8f9DuejgpDrHJYgYITLmOQL
ThBihJY5iBJ+TJZFhYFCml2rT5LsFmAIWlMB5mhwJxVxjv/1bgD+/Ar08AWO04NS
sOgfFSV0ZRu8kNLWwWLUlOuxASRm9wu3D7gnyreOo1/TSnb8T7/IsdJOZ16ITy87
JIcufLYkK1jchclfAWFz018AKdYXr0B4qP2TgY58BFO+7Ik+Cs/HsoJz14bTnYkC
o2FBMtfxK1TcBvXYKXGXCwInwkpxRZh8Aepo5qPODifErmcj+z+C52cAguaxnN0v
LwQExIoXNJKJEtjp5BZNa9lQYq10AYw+NSbxaUKpFE0Vg9eaZojJ+lKfaZdPyoV4
AstSwd4jg+UFVH+TTSohT289JHM6hQv2Lc6LstlMDC91TwOFXiD2rCC3YZSI6KLe
sbafgPELY3RBSTQEEWWNNBGV1q3TpF+N0bQm8YVKmJMX5OLElHH70vno64t4TCYF
16JGJJvjOnu18RgkHDgbXAypvgG/A7SHaRhbTc6Vf0u9aWIlcCoRnW71FBUihZuv
QQAVJ/Mq58I+pCdWZWjQw8hAC1M577fMsX0z+nl2DrcjkYXTrFC1OCZge5dT3I2O
EX7vHnlFP4ETjMYw4RqctFjSK3DXkWqUPhRe2j92OEdErlphw/A1TS6iwQzyJHNa
JqsNe26Kvvg66L07omour9ZDF66Hf8WdKqEHBK8WREOj2ZtXhDTB/6fDy+NE3TAC
ACs9FzEwdTxS6MUKWOoeZsboZeriFGVVfbSTaRp0KGBBXZunsZ1iJR1kZwlXMl3T
gAIqj8TKrfjLakU4GIazEfPC6qJjplz88lH1jS6VGfl3HqMipDtN5M4LaQUrkplW
7a6ePRZTlobnqpsmfwgPS7L95aDd1dTrN7onQpJhtzTaVW0Re5M7vb8LS/Y3BF/L
eP3n78NaUok8oOVFVFdbm3fc2vmP1KINIlS4gYhBZtr8wrzliyXWtnDnzp6RT2nZ
kI/AC9xVu0vzlnIemMy8CzMQ1Mfu0kJ30C3CXtqz5JtUogF0PDubWBZ9CYGFaJSg
QwWfgQEUAyJEsuC4IChYiXZvhKoSNeM0PzTfVWZjXe2426udnbDxxgbXD6+ahz1f
mpSWqEZOxFcDjERbvCDLt5fxtt1OZ1hHY945rhWHV3Dj/ubXVnO78HiHJIajME7s
Xm+Tbfkp6VPmK45loWdGzDW0ZhIcd7lrdFsBJ1Jz/sojGZiEft0idyGWMND3Ietu
TvWhYdrSg7zQqigl1ln6DF40RdatpnhbfN++WyFUMjBqi2BDA1fDSO4ET7vNTcr6
ZCqXGmBWQOKbwqW+LB7qZDFMgBi5k3Q8iGh235MMDs2HyINN8jgey1Bfq7y/2WO1
/JFJd13AOZgEdaRQXHRYv7e4RZ6OJ/l3FJT42hnW8ohVn97SAnCh8usLDm+N6cip
I+b8PfNH8cAenCzbTpVv7K6FE5hQ0Z/ysAtO51e0CD4qJ87RhRAXZtdXPrAe0u/w
s4085WxYrrAwb27Qw+2aZYMM9n0eEZlpIBiOmT3BdHYqrcPTlRsFCz+CvZadhDuI
imvBlkulD2EXlMYt5WTOf0e1jT82q+VILAFh61/aS5y+RZt2fLFcVXC5evlb8vcJ
cHit19BrUfbtaXwooev3QFrcPU1f27wu0ul/UZZlELYV3tykYhq4FT2dtlBwPTAC
LkNq5mlbgMJc576Np7DyAElGLUQVrg0WtSXUok6S+Ea5kN8OzzPfiT9TyjvpUqha
8nomp8MAtcbAUn10mtSlU967NNYONyTGoRGFdt1V3RsL0d1Pn7z0KiP8noBihnA1
eKvR8g2loJaHk2J7nMZDSOHWWkdDUNteUS3A3ZqwZStRty8rDUg4eFQKRYqg2C+x
tT6W36h/wRYeHxSQYseTJ2/dWYzC1DbycU3YGKfZhBhvtOovpDoZA/Ia+cTCWHCv
gwfrxG8PG9aKdkQK/N53gC2SP1XMxKoUmzddhGnlf2kj3nFGt1+kGaVWPRUx3F7i
M4q5a5mEuOiQZ5T5A9J55AF8wQZ4cAB1WZObQorJfAVSHjCldruJZoH7JXGruO/f
dTyxuRAlO2RV9RGVREk/J2E/oe9YzC3HB1XjKW9nOfu2DubZ1t1raqRalaOAegXJ
Fv3JEneVcRtIx7q74xAjSrgF2kTIIEgTSb6YyKe5+vjXK+av5EbGByu/nAaMlBGo
tu5XLTZmjYTFwes3zbV3VhRsXnY0qTgiNf0+E7p8Xpl0o8nyudXrgQROunVTSF1k
LM9wCVzf9BqsgD0eYdu/9KkydnJ3xEPmcsJBF4cyvcLa0UVV3ptv4AQxUByN7n5j
JAI5G2ttT+pVu45M7OWAavPeQ/ojYhvrTPgzeX5Cdjnm/crwu1+3I3MstGd3nhLf
gjnLSU5sO3quEh/TR4r8faKPOiA+2gLk2Xu8ecsqqplpl6VfPn6LDiL5/bF3rFQV
oDNff/oxDqKthhBe9CAWYHBJ/IMz/WyODqXfvEDuFG4yWudMgse5vT8txTlo078N
7HZrGVZO5y/DM+X3tLWEF5FBWLgjvLoSm7cRcGo52I4w0q6n5z61912feZn2bIeu
p19bRlbtMSUdmZSkTP02pmbwqo0Q+sXngf9DtqtvpoAWPlc6/h8QXoYAE1ZPHroU
otMlgIZH4Vm3Z64qJBws708/51V5RapdsGmQMgX4A9uNbp+meHildfxKwVMUj45Z
gRNuVtmj3qXzeGDQ9hiCKZV8CtpDRbz2KUD2zJXYQu9wi51ZCx8wpaPjLrR9JoY0
45hoCS2LTsvOcY7u8UPMQbMuBRoDe5QAHH4JnI58XVKQ8VEWGmazW9FvcJJOSDkq
XbUH9rbEYN9XqbK6++4F/VNdOEqfj1yZ9EaDzLJUqpQuf5qqYqbb3JB0gn/PXHxR
kAUBVsaB135xciTqD8KKIcUGoCdlyBtLJe6E6kXEQ6O7hAGYA2DSHiUzHSsuNF1b
OkfAS0hsK3a0/fKQCbDvcfQ1+heyB0I5L7VKyh2Dy3+bYzUreQR4YKmIjdYGfGW+
NfdU/BW7uQw3bHqrHuqp0ebkwGsztLsIws14+hXzOkTjkomGl+XEddSHrqq7Fp9X
/vG/SDvoGVSVdzeHUJW5qW2lh6VVVArw8RFt0knCnPT6X7L3KbhxTILQk2TI+WG9
RIOlVlp2LBvVaoIAToHgayrFEIAiNFC84/mjCwa3yqsu9c6+sXbCYAQgXub4ghXs
RvL5Vwp8BI/QYBUBUnghoWW1z0bjo3AkfqBPaSKmKdNP3Fd1jCmyGD/7OLc9r9OL
1GWk1sVkEsGRsj1+o071OmUNX/69osrMCeV++WQQiMCbD1Is2QmwYnjJrBnIUD6p
GHHywHLLBRFY/gzCOajtasmwKQzWesuqNtYbFVvMykecsajqgS5o3hePAiuBEM/5
GixELAkWQG6cZt6z/sRC/x7AqXJZh0YluC7IFujUKYMXHumR9i6gxf4Wl4djRWjq
ezU42fuXriun+UThC4srBPqun+hZLCWz1657MGCn6epRMA1BoiajBKfl+9imijjk
gG4dVyZ5LogfEzVj7W4kQ9NmD/ZWCYAGxwWHboTzWiYH5WTXf0DYRN39p3ULNrV7
nyNV7iT6Foe6ro89+ctjBnI/HaeB1h2w5Xc8Z7fwpZlUNUXGLNa7vTv6UDoAUsuw
fO4ayS8M5YWoCYVAuJST8NMCDSGzerkK5uIpuNi3CrrwbYzTD5+kiqUEZA6UzkR3
bKKOQbuAIVNptL51zHnZJOr6Hawf0lggyf9YLX5WyU0W7uWmDSC9m1N3NpLYveGr
uRGKpEOEfCC3rjooPQIRIjU5XVx3wMz670ZR1hRU090wV6i/c+/uSk0zfYWNf4qM
CIvE+xOdvKCG++HrTvTpIuG+CsYSAWB7GGoShJCheuzCz3HAtcoU6m7qZymPV4Ws
P7Fj7FjYOMiWDVKFgN/zZQNEPxKSN28QyaYnFrlgQNuWWZOe4ROK+tEvKL5Y96Q8
KcptgN7P/bYwKkMTqFkCSLCQg3WJU1d7uzIz6rILbZBVJdZZ0DBQSxFv+OyEWnos
ai+twYdmSK6+J4LdmYcxQJFpeC8rBerJP9rW/WGlc0q41Bj6p8aiaNFl7YExaRRU
EvPncRIbJL7RH2KD6MKt6YjEs5j2nIf894uo6S/2fWAam4kCdDSJALVbzhQDslrG
4N1jkL7JIynIBZghlSHJyL7T4z3k2TeY/3gV95WyqIm7xWAxf+7Ds+daGQBDk8vD
+Pc6HdvPdFqH0c9dGsca/NYaYNMPJlUKBMKCM4bPWnNvCgxZ2TpDhwT7UnoRj0Nv
UX2J6pbj/LWT+TmelAWT0A6EoZAUEHNi4Eunsd4z/C3Ami3nJC8ilVj4QwTqDKaK
nSpjGIyHr3PAFsXc1ggiNhCj79ECHDcVtjdfGk0KSDHGtEzIrewalFxQVCg1IBci
vDNjrR0UrFIZbDvDBh1jUMTcmm+XZwTBPRxVXEpC8ypUi2kEv9jtZhl4jWSzcohE
8d+wJ2+Dyxw61mRnRg8dZh1WXtGkAPmcJQV9v+wdNQaYo6bMfFO168mw6I+Jkdh2
5X6xnylVb96Pw8xA3fh2WrQ/0tZb2QTAMroVLk1cbHOZz/PcWiT+iCdWksWvpyK4
ZNNKgwemfOIGTnHaGiG7bV+QnS7I7tbydQvhDX/GVR/y4pIuUhu+yHlcNzh7mBp8
WJTJdwKztA9OsgbrsuurWmPzuS2m8zXb/4lv280frhIMvFpGqgeUHCp42ujH+dW3
/IR2nJKrSLAmsKYq2IfMB+H+Wjgh/+QyppnhEzpQffoGUThHomJVu6UL9FNPduXq
Mh9knkQooGPOzEfPUicJDywSnpHDMuIE0CqB5oWvqvBLL77pvC7tUk/q2TXRDgAf
JG+9NcSMHUEYzApyWZpCwbdf0JmCfoxS/G0nTPH6+YNtFt9o5KwSsxH2ICfqJAhk
1xwoS1/a9fIVX54WzKccKzndSrPCjW/yiTkTv1erSFakxHP/NqJwldd48fC1pBRz
SHVK42MJ40Vw3+wMty2T/m820hC4u+6wg8iyS5nSP5rnpLYhBZnvxhrR30LMGH9j
LaDdp6V4KO8H4oPwFjT6a/JmuvHvptGGt8SlYwYu6VW64FIGk2cfs5kH3RwROb+P
L9Uc+GNuGGgkS/XIP3uTQoo0ptD88OiOBRgeTxnx2gz3KAw5rxQK4PswD3+BIJzh
2DqrO7YViJv6iw1Wtgh9dVUjjQfAbba7eyXOodo/Vk6S+PAF7NYqZkgJzF47dzmS
kakwmkU7HJdLMt/V150gacuxc3JlsEt/pMNFEX/dVJy44flhBvbz7oyWbLyX/gmx
092Y8DQpBT5W16nyBrkWKpvo27PT02+Jhf1E30sg4E4OCW8X/VjSHOsAtVdnGypU
UYdfglyYUMMF1rY4Q2nnRke4rxIMBsPXRG/hayDvRv/bSCyAC+nDv5LY3xS7Y1rI
tyzzsG8DlubKGCQF22kROPucG4sF7Ix24eP+T5FURteBfd1oyC/HsgMHA7r1aKWA
Qux58TCR1jMs5Rr2gAr6kVAnVnyzUF5sBhMNxseAwExDsN+fG9FQvIp3gM7O5X0O
eJ36wlls/f++f0Azyb3oQtIHKVbwZCE2YctN9qk5nCZ9DS0QY6SoaSxrwmrW32V9
4RxqdGd+0P2hLFYenhFiXBDUJv30wcTPU7xPgN5AP0UEHz3fuKuLocijXZohtW2q
Hj9r0O6tX8FkbFwNcNsiKcOA0HXoCIGTIyBpNUO3jJyUzlC8ceJPayZyZQAbVMoK
S3KmaRDTS6Fza2E2En6SWZexLKA3fKkkMZFNwIA2QLmVuayb5lYJhcA2VNvM8VKz
pTVRCX1SDHRYJv/Fk+TLK1tH9XtNwOnb+RfOHSdYzfZd5XCfUtY51IPvSIdMmceJ
sIZFug02V2s/6or77dPIjoyEsoIAr+MxrnyuGV8StoKHzTLBMdFwWD28RuiiJmMG
8k65e9nxSOMqL7GgymQyg2c22p5c/xKxRgnsNeUi6NDL5dG8sSdSO4KZmYV/Nlo6
+4mNT1cWy2VuJPMmIz68YEd4mo5/MoSxekUozTIKJBTzdghArQetGtj0jb2x8bFo
pcTgIBKuvHNect3szOO85qcXhL7nEopu4ScrBdpUa8Y3i/dCSccbWlz/LOae2pKa
UW2yAons7O+TAIyodW/Cn8aw4VHvv1JLqZkpTHIcgYnYeEyiJyHhbhgyhkIytqv2
OEuJ7pYypj/GNbttQylUCyL2OscPnamx9VZ42BIgUPGubIVSAPKkwV8Gh4WitP4S
dLG+voTBHZd84we8BIcwuBMG6Bf+XlrIYqIZoJEeDjuhuVOKjGbkBVlSWtF3tlLs
lofDeZeLVQWZfWVQpV9WzR7nMKESDjDKd0JcyWRg8SKbVQxFHH3pvy2SK+hgw1C3
/ELxOOALl+QGAIFsn1nmSjgp7mrtTqmdSHgVILCdfRbzDgqku+e3ZlEhCTyxVuag
mu4hgNpMYB197Ox9k182VfsIqe8TCL0uFj+r4cv5Zp4Oy/Rx6N7evIu9pDvDco45
PePBo1xhas9kqPSpdYv0KLu2U2A0WeeuG6vLPYSJ0ndB76l3L7zzjqLshrXC9pzw
Qxy8tNO7xWdnuVZk85KHsFG55R6KM977Koes/hGPAlBsIqq0rxSfUQ1OZeBLymHf
kZk8UnO+9VtVAASjEeMzJH80RlYSLmH4o4ejACLvyH1dNUkG0tfURyrcbstWsS2n
Bjfa0COFgz+aSsrXMfUeu9tfYGyEeQrdohXU0GQ0sbklQvdm6OrGCZGlXPT/Eq6P
M0IwlXuKQ/6eaUPzA1den5pjyGmZja3dGoE+ggdQZm1+Jx4xZXSbw2Eh2pA22SpG
XBy+4U70sRdjqdjTroJn9pL4/vJZZdxCCbtIUVf/iVOy4UaH6FdKNAhfFw/NHErE
oFeEfobyO3OTl3tb65O7Ix329IBNhgvWc7xzr69yB+oEOzly1rsmlM8lvJDpNu0a
OTq0pyOD/4IrUKrtSQY9wym/6RkZJ+HY2PgVjlZhlEXgRb+Hac7o75QheZwVWcef
WkuTourYTSKcxGXsUxRmOEVDT9ahi0WDpbxNBEHxf2+xmI0q5V0DpMzcFTnFMXEV
VsiGiVjnumrdb/FF4IhMYC46T3fJvDQShuTW1CFpj+LAbvFgSyRcUijI6wsIheRX
VIb3jiIzQTVhNXDrl7tc1M8zeAnJqjH/A5B3SIITXlzv6gA3BQ0DwtjcLX9iS/2f
aRHU+AP+TnxWbma71OAPXWPLItraYPnxU7djy8/IjZs0pefhN1pIjYmfr6n2tYjo
U/cl6mXuY2AntayHYAE14XPzmOkqvcUDBI4DBcnnVmYwCba8tj767SCaqsdn3vJS
q/EwO7hmi01mBAobpfXijojmhs266WnttCuSlYWcdas7Fj7GNxdZwPO8i3waNdZg
mle4c5/2jUxFFUyGe2E7EKAgjNSC83rP+M2utOTpZyHpZVf1ZJVOu+AVMgh3Jhu9
wHTgHGvzSSdVaiaPtRQnHwm6LWW5vVJArrjSQlFPlGC/VEtymxPuYqe8n8Fykbp8
RVfmdxwh00+lrJy1SChnGbpjKX4dFXO2hPf97bd15fDbao4WoSdM1Gljigh2MH6L
gF5z7DPQmlvZVi8G5dsscjL5UdKi2QHJ9aLGTBzYMroflKl9SkPwet2ad1Y+C3Qv
kg8Oi1QecWfHgxOpV97/aRZbwofvz66JMgsEOenAfQdzncKRiDkh1tyAgFB1x1/N
MfC2GSMH8WYAsLP48GlPlqpV5OMeLt+LRQ+5bU4tP1MKvxn52L8YaV7i2jmhpM6j
7PBk8OJWNI+b7MFgSw6qK49MeAbyw/1wS7lClIjPyjWvpFd2o8E0J52FrTJT4idC
CTng8wRVzSw1IKiIIAeU/YbLchFMYn+Jx33639U0jBeOjwDY3X+6apmtPrNXIKjU
sgWqLLamCQQ7/x0eoaI0zmFUwXi/NszzolwDPOXOUXYW6i8kximmoVYqrfWghqZD
QtVi8SC3xQoxXulHEt2vEUaxFzKEFcpMGvz9Kc37uO2f6CLc11pKamNHfjNt3suF
IRYzsW4EO7e2pYHsAXRBJjH78nTVLh7O15p7d0GFjiA2WiYaOAK5wrs0b5NeD62s
w59Eiv+xL5pQlSVK7gVDU2qh1WyvRHzWQb1NzjNFilL4RnXMWIkTigvLdzY4M+Gg
EgI57KwWyvuW9DGOVqMmt/nWgCBV7BKboFoOMfb0UJOzr0SYJO8ghqf2CqKTiaLT
Fs6H46+UJKlH7NfZzMZHtpovOFamOXlDDjIT2S+R0d7dILi6n9kmyY8mY0G5oiH/
6pRev+Qa5AaWl3dyKgzMa6VWMhom8UAf+uclVgt7gFRv4jaUQbZCg+988zX8MdFi
kNO9Zz9e8KS6BMNaA/yyRjumeWhXBDfCMRzekdus1e73lyGTEruakbjP8yLLwYtW
+3d5TGprvux6iSn4nctF7NdIggXB/bor++UkOpTCu1Wh6X6hcJMGZABhTTLi7n2V
dG0OvZ770nYLIdMxm5eoQDsoOkkbLwblKK08jZtVBASbro246IerGJX7z/3Lm9Iu
fUlNE77JR0L4RV8JJ12wsbhRKtq4LrmtOLhWS9maZKWzjwYx525VFLZIWc5/5YjA
uphMcCKzATBU8KFJkOAuKbiFzfCn6bv1aWhmLc5/p/Q0sMhIaeahQ+tQvSjCUpnw
3NuTyhSk6LFV/MwGfGKS/0vwLDvqAUvteFntmZTrtJxxpEWyNvwhUDb8+jGYrHGH
SZfA+c512OMyoN9z1xDuDQbwXDsJ2uHN8HVJvtZEZwuhKTWhq5rkMKd0RHkaBRCw
SO2oZzzLJIlZq3/yCTftNlrb3RDQ8yLWZSnNAq/YIlZGlCsik3N82JdlWFmkE4jR
u/XX93okrBnts0fir7H4nWKBE5N1rZDuZCQhaLHeLO0bHmWuc6vjBrowfjcKMKCT
L1Bw6cN+14qqyvJuhZtMNWiUp2HMdPc3zdGBac4EkxI08EwM4/fxDw42Jjbsimzi
J/5lqKA6fwJtv7Czaap+f5oaER6HSMcjBROKChuJnofDsL8YaD47rJaxq7gz/mUR
1M7Svv1R6pgOfCNHeWtIBhf59IrOlq4PB80kGoH9iav527m0mF8eWS3HNwg0qFR3
hZGw0955lTE2FPHPghE5/wNHOZT3pqyDHr0QD5g7FXBto3DfWPxDHiOxIKFlbB+m
HgRPQNcxxQHiNzqGryatr9wJS2r/7+bsF0fWvx6a3lWpxrQfvu47ZFZTxeQKgUW4
BhbulN2WRm5i6sOf9YSKQUMorIFMO+0dSAQBDr7FMDHA5LNOGJztSzqL2r8qv0WQ
d7XtHf7vw6XNVcV4W6yMKWzD1ULsaxmA33T4lcybLQWRzuWq1DqhCN8NSUtkdENb
crcH94pfj/uqgFA9nKuI7j3jz6EkYSkl/71iGS52UfCPM/vHBC8sC+DkTu8k6EaG
IV8ZX6BvNZyVr7MRHvLpgOJnZLnKwexMz9VS5R/nHL9PXMqYuaEFDT/fkpbQWBOZ
OnzVgxWLfwCIbTutKZUuBggksv9bTbNmdfhq3kyk7klc6qxHPREpgkJv8SDK0pi9
iLVkJFQSeNjLzD/2GSVbwNry4b+oHVdVI6saWTaFvbkP7uypS+yuGyG/Dda70kG7
YqS9C8ygow3AdYQ/bju6bEbkDuOLKCmOk1qd5kRK3gMHfF5OTN8Gep6uXEoavjPN
qZWAwf54R8Bc0Dq3159b5cIwcEfu3ayeDoAfdgNc85++gwK7V+OwUwJfJAdXzSJC
2dnpZQ/OzcX20eoD0zHEwvVN2IaBZUgvrgDHOMaLpLZ6fR4SEjtYu4/LHH0qQtSm
ondji6oAKSSLkK20MMNlQ8/P8FfUpkPJadUKPfWFLj6nxAzkxjUKJYKbYboKbVOM
gRK6aP1l7UzUfBpPHiyxZDsPegJ6tz4zWkHDGO2383WuZgwPg16tm+CqAEQZLaoq
fQ+oVWy4Qe25sNqkHnzHsNohcx7DZSXeARVlM0c9uAFgbhsc9f457gEXM33HcZbH
VA1rWM08i0n1ehV5la/iFWnTX8ZKmMa8XS8tYEMVORTJcEx6ryaKSMDGBs3btSE0
CsAiaD8cSbsMcAGGSjPx3RY4vG22hkydwJZN4ZHqkd+feo3S4vup+L8ejSkmAKI+
aaHcwlBQ+63p2WtqwuQLJbyL/xFPMLciaN5ZH5Jyxgn6C5zFirBJVpd7PYKn9Fia
VVEgh6LIiKXwgRYVfCO0G72r0oE+bagidMA1OjEBqWwE8jiGCoZ+xlz3wfA3OfRa
x5z9PCkqrAie+R1gAoPy2DEVbN278RxMfoWDRJwdBCxIj0oCoIKYyWesYwNzVHY/
zlWhbChCwYyXvdJOBINvZhf8CsLD5lwYKtCZ/g6TrJ4Nc6VmTgZObh8s3bhNVf/Z
aVS8xqtgi1j9ApSsDnLYU6P17fesFhmB8AsadWZBcogzlLZG10zVyDrSCG5rWahe
qkrMphzLD4j2X0LF5epsTLIpTZeEddc6uHM3sOTIPo/PJ2S4ABmN6pg0hPsS4oFM
MhIJOtXySsOm/i493MJoFgB6aQ2Ccl0XNwZ1RrpWI1S9rvEghyP+H0Q7sk4bteep
3SuMqUJJe40umi8/sk+tIKTMMUSPCLfRkCiKzLohXYKcG2E5NkkW/2FhGXsPqw7s
hvIu4bxIZ2sf3J41u6VwdF2kar2E2V/8YQlTNkVu+ECgcOB3uqlbo4LXPijEfluR
NEUFiIOW3U3s5Y8Yn43kj+p0PIli91w7kiFVq0GalLdYU8uihLP8N4hc105Yqd0F
b3mC5kIwnLn9R/Ex+jIaU6qg6XSTreIjjS5iDxYgQLfUWvj51jnmJFsQifj1INgv
nzukuNG8nokBDnpe/S+FYKFunmOs1PiSYcBpSR9n2FuMMkPOwaj6QhptHrp4qXkY
eA8teiG4ZGK+J6YI9evn0y4un831zq+KW3d+L1tBEpSsIhq4eiIkj3klbwJWCDGA
65+648KEFCDjZw2ulsDFktrPXyZPh35qvr2hqwHXObKjgsz6XBeaw6USWOVeuuXm
xVZcyzpx7iU8I6BaheJoVIcP0Zs8zq82e5ljv7dCvaqCmwEkNRyQdQvD33HYPHNz
0i6TfGp5G0RZQVMdwWavfIIvfKhifkcP3H/GHWn1Pms8REWWXl/TnMuECPIW6jZc
o0ywmYUmlqytheDbwlCE8cN6mBXTfnSrYVdHoZNQUpX7X7x7Z03v7xvtNWSeGVhB
y/PB21hBdI7QsQxGXifIdTMySZ/ZxZeZ6BT2bkhK8Hkab8ikJzMA0MSRCvkszqp0
h3KFYHSYPGsJcgp5iJeSU3Bn3cRrFqp6BKUqzhkMzjNIAePpprvoStZh1zlpfqcy
AYKLguubPHgMgw7DNOVC04T516NRUxvQJKN12tsXgVwt0OUW6etsGTmvmI2QtlZ4
ryJpXLX7pPCsS3TvXG3k5+ZXlNbyuxhyqhi6XnPG2Qf+VcFOQu/kUuyhqk9zARuN
pRIVk7n0J2afYFDV8mPMLA41cPULkuc3/ZZ5Af/ORheciwzxf8vZX2aMBITtJ0lZ
vSej75tpU7iNEOOMIho2MsVDE8FzD3u6Ew4zlIKOapUfhOIKZLNRXy6XbfiJiIiX
bW+rKVPIhYERR81brVJqgYTdMEmNARd3FkjxL2qytPU0OJsRovEctE2aAFzGZqsZ
E5CUpxYQtYdCdXnjhhK8zD9q5oiEaVLmcB+1iTxOb2dv+QgTYis51ON8kO7UMhh0
0JkYcw+OE41/ChMnkdKO31oW9k+/texqV1fMiaiSb+jIfgWNBxKzxjDgngdpVmTL
EKgPwRiEgHqmVfVRV0stuiv1E2R+9PNQ7IadyMygWvKRhPGmVoqeRBU5ifeEmLE2
kjTmbcyk8Ph5jnr9xbJejysq1hA9SDTuyAQoHLEiVndsuuVU45NRiy3kY5vlZIg/
ZndehvIG874odRjvlv8R96gPWMlW4u5QAbDJS+hiIx+7FdzNxeR50j/5t+dRdtRH
7de/kpiFDbE9kUKtU0MA/Q8y7SWH3p4PqkAej11QuSxm+XZUexl9ojYPiDACH0KL
2Fc1zb0/Qzco1v5zA+Nq0cEoo5ktJEqsIQj5G1v7RVTgNI4vACoPAOns+vol9hTk
os9cazNvUQY7iiyZc9s+U/e4LM/OZqTZVVyfGqujyWjWwS+cyNQQkxwWygFYXXaC
g6vCD1w8CAR1rH3H0VVjN5/qAhAwcPNLjui7sHQh8/C2W6q0EYs5L+eWoTncGOwc
bfscc55qrwpMM1UH1gqtHeM6N3lVFAzU+AsjY3kTfxrleO3QiCDthT4ulZEjtjeX
d+KjtyMkFn0TCM/Q3/YhG2CFcuf/WRdvCiDQRS3Vki6wHcdM/e9znnB/BmF0BU1r
KDZdz6ukZbErpAKb7jczHNz1FrMd1IkJjZGB8eSFGKqnMuTOh+BQcvvQbF66P/Kw
DUia2rbfdAqfwxpZIcdLkJ2T1EsS3g6iQAgotB8ZDNGAzqhfD2INdlFdCNtt0aFB
UXmAP5Xc2eyhLKVJtzoBfJkSP2Zr+LrmN5igkDRRlukA6zUvhq8Ph6a6S6fjnCPb
U9ZmohyrUYztz58G/onOjoGK1NrFarkk2y0f1KzL2Ap/bLNh41ej8d7rH/tHXsqn
0ZcaxfY0e9/QfBlD1nw/uABBsyBxnczU5KgTcJrKQ8mCYwFweOqiamt4SG1/pG7h
ZoWUJRKUeQbwtSw9M40lQTJsF+/BbH+QHfCPRqddROM7Lla3ag9ylJkjcgStUC2n
7fdmxrpd6Qhlgkh4arpgxFq2MP+gZzPokmGduVQ0Sw9TnDUaC3v+iQYQZVqqUVDL
QX7EzB5Pm3KAME4GVorvJk1QEQRGLhJMi9dhxAlMb79sr3JtUJYWQeOLGfnBAjk8
O56fOkshbqBpBPkQbFUv+G1Ix2yUQ3rxYQOGQIbhGqN+UJ/X58UiAlzqmsGSutQ5
He6XoiSaG/MlW1nBVf080d9KhG3rupCzNEsLFcTyPm8fjmGw2iisGFyfnKXfcujS
rj4svS301ggp6BINv/lxFhJ08aoAGs0+epY45k+zz+nTYL6wXv9rcVGcKGXBpYCQ
GNOWPBsivHqmO8yeQC4oF+8k3bUeHkZYlncMzXfCOFmzoxR5q5dz8JWTwe3xmgBs
SjwJegc9m8fh3xP7WYz3/TXPv8bl51zY4Ms6vCbBe14ZfcnitIqfHYWkR74NBqxy
yYNZO1JR0Yu9FDGUNfIBTRrffdCnvx0Yjopkjm12NRSHmG4GCs1BwpLY2vQrUXiq
DOTw1Nu/P+3NXOLelSQM+QbxBJm2BaPhrk9FvuVhOj2ztad92TeieHZf9nSr12Bi
2B6TkpmhrzDkf8DTfPEkm9p+vM3b3jnA1oDwutbk/DT1PXOpmYNOZ1tdYk9fIppo
4JfhYcYY87Ia3a6FSJ+ifA9e9Aaca+1E5sj5DkA3jzjSxNLuY4LcAF5cioN2RFwQ
/cEUzgkwGV4OjwNuMeVBRr9aaDUKcZiuQDHEZFmOZYAdWCXKaKfSs4uNk5eW7lHS
vVLjvHEIjV299xIo/04KygGv01nvyn4vZBx5/UtlFNtFWe4j6Id/BoiI2sK5gTNl
R2Pkmj3AJ/I2ERpij4L+lqK/C0UutPJ99BUNNQDGKA811iT+NDMdvAWy1yEqc+5B
Yfpd6wgIizheqPO83gjtXcKQPDtwzgQ0Hw4WkxpWRIbtc6ahgmB75B5WqsTE6l1r
AUO58oek5MkWwHXyF5pbsZnYFUX+GGpxtnNnd+C1SrQMua+OZXDgCXw4aqWGBQF9
cPuZXR4e+XoYJtWXegLw5HuIXdIHikeRtVIrywJxpKkte5grjG7Ix31Z1QiVVsLw
BM+QYHUX3Fy0Sf6+lix2fBT9Tv7Phu6MeSu0cqgQeWoLPUxEUlUjZI1m3FiBCQCi
9USs8MXbFtYgtUA8rudSpVOjy4P9D4QxxE/31NYNKdEunT1thTpu4Prw+ZizfVl2
oY86QucCV04dhlDiE4bkLA+VwMuREyY78SmdppzeKG3mXZTrYCOMgE46F6Q9is6q
KSdMnmKaby14izAYhBsw5P0NPcHbrFz3Z7nPeWNUhQMaGJnSyujQ3NhJlq+ATpUY
LedrGnnfYXV4LU+pVZDRi9xlAFL+QsI6W7VXcsJ5l5TGHAlGboXGwpT4v6h3Cb6H
Wy3VK/WRCIFZJNfxWkiobEa+jJHTma2wGJz2JPd+OY3lKTfPezoLnU/NFfbmKHZs
RFPg3n9HNXBSeFjLqMm5m9ia3UmL2iT27/7v6RKSKX9EfLmav5oz0K+aslbbgz5B
VF+hNNNRjf3vaDVMRGcM/BFvACFInPgFxVL1xEDK4aYbCCIc64njue6U+xkMYl2+
xnpdu49GL1JPaSzehmQPXqfraTTVOAkq5LIHMXDNehvRf4YdKo3Rems5fFKZzEZt
iokxELWjt63yvzLAidkYd8jzN6/DP0l1nizVNGt9Bxx8aOWfeXCgDKRNPsXwyE/G
p+hwwIvIN0ZI7TOgtvJJ6id6l1vyUXnRjd2wu5LBsLuGB2OfWZzekDXNydjjdc+T
v+nJTyYHiHd9EjbunmRDm0fIGOrwF+uEi2UiAZs45W4RC9uR4bKp6J4DcTmCuYm8
7H9/gumzZfBS2WZWbdFQsb03K71U2ma8vz3wvvfCpD4u8EsDb+5sALYJV+4hBCTa
3mNCEBylpiNIk3T9hZn3lxzLyjGkR4wsKVorNZUKDEPtTLy/rRgVwcMv8dB7t8XA
mxMOI2WBh/YEzXTpjshvUehuTWIdoNWJiDCF+dT/3QPxD8d4UpxMV2XvO8OafW52
ESU4fONLB6bRX4cgTXFNEnJC2jF5bA4Le35464GgOTMtrrrQnm0jLB2tJwbCUVvb
qSNm4Dj7pM5fVU/BIs9i3tOIl5vD+pLpC/gI8vIX+GRQHshvfEbno4qlrEPyQ5cn
LWECyTDsnOGQy1XBareDW28718iOVZfWfHAIFjmJHZLYukmHLI4gUnP93K5d6+jU
d3mMCWK0Ii0W6Tkiaxzz5dgjXGJWgNfeeiJYdsHoMnAyvRWcLfe9uoW/R2yZetVb
B9ytmUCF3x9PPWy7r+Q9HzNCmh9vhTymi8BLIi9llYokxmJg647NSjqQu+F0nruw
KX1AYUmPeN7qBqIF5wIFsIHiZwxIerK3NPvWIn+OSTMD+waCiiCwT2u7Rpd4q5ue
61/cDg3N8Z+DRsOPI/rRhWJy2FbdHuZ3alVcngRXkjZqkd0/WHlo3BLoHTgmR6Um
5AjG2/5ww1ia2s313mwYf70H3SvANrbyGKKV8173nq2K8ECkaxuovSTm+aA7x8+8
8YGVPb0CpBoufZzba+w1tQFf+3IQQZUW9cWgeIRH4J2jqEkI3WOQZPl5jcQGO0nw
BKeCSUkgX6pdRZoa7ARVL7OAdo+RGLw4aP1VMz9bnqbNeVPAessOV9jFzxO/4lT4
UNmuF9aLhX2VARPsAeE2iPFvYzGI/+6tstsSLtZYJcnbyo4xlw00koF7XEViwQwV
bPZtz0wCK6qv31x3NREN1zKtSOYX3DpTRZ6Wl/R3+1S/bbkAJ58+Rgn6p0zBARt8
8tQ2eZCeVyl2Ma1JNqzteAygj3EszxNjC7htsPTzrXQevH08V7pzQe+TCUx8WF/t
+5+XIrhAaOqj2TYWD6bLwwakOp1Ys8zIkzvhFPFoSyUxu1030bPTVSJG9Rm4yaKv
cKIF5b/j5yFMUacy4SQsnCcAMUeaL5KQrZzdEjQGnD6TbmyPszo6os8ktCX2sFSS
xgC1w+H7yiVxIjLFHoLAyuZseKSjIhAui1ZXBIzUElwzLM+749JO099qnj0Qb6Ot
fDmHoFN7pUkpqm+8TLJawRWx0TFX8Wi9881mYBGsx+xGaSiSVdkmsVemuZ3ojTSr
K8H3/AW731yVDY9b+1knsoP3VImDjVaFFBRaGqnC7an9+Vocmzf4LyOZbAWCTQ56
hXrfrcyoLV+rZ44bC7exRlnChFKyQduhnY0KJOzB60Ekema/dlwGfmnvetVSN1zS
nFVbIzdJqdZ3TNLloYrTEpjUvEpOtfvT6XfAqrtqqdmNTirVAKMw+j7qNIj4IWRS
wRKr/uQXzDZIPr9TzNlNTApIGJbidO7bx/+2f09jYJ3H4CDdFDahTQo7M4BP4z31
u+QAcRmBYG2Xcj4AacFW773vmPEBzPp+B0ng7/V/HkoojuCwCdQ+pBetvE7FjRhR
Psmdak6yKIeoYVx3eo+G1Usv77+ZKdEGorK46mBohq8hl6R5qQogocJDkBRS7QDJ
kvcBk+4JfxIceNfJel/6ekBsg0mizvSVRGqfFFmr2r2OIF/T/w5ebLjhSsSfgiCk
mHccbjgAfh2j/x1MQM5tgwBdMpUYUPvjoWhgdLxqREDuM9+eOZylX5MkRw4dYTic
WwOTU/NAiRkg2AV/2UcFIHaCoKZc1buDZv/EGNNCjuvZF9icCjQ9ewj1G1neNOWw
95DLLPRF18jUkEE0DP17AA19rHjCUdtl3SjgyaIRDpy3J50vfZJ4LyXPYtrwdFUT
EkpNwa3MMQvjVvaapGvM89udmAMyLlobxrIjadGd+oTgTyRCd2t12oQ7jgQfuZL4
XkSL/CWLanSrpWNI9PKdRRYV2FgD/mn+2YDzz4ZTHPobnx4fCmXhu8byVOMMM90+
QirHDMtElpmVMsr3s3mWqKNburRCyKvIYpqOlJi8vsfmhbvigWCas3tamT7MMg3W
Zld2G2tscs7KjlJFpPBtUPeWPIyDz9IIhwRKfJovqoeu7CteB6rg5BW1nPkfA4T7
dmkzhk6wtXzzD5tJEHMUbOWwMJkW3wmz2EUZR2h1wsEqUDAekUj3KrVUshhtnNTL
9nWUcshOJ/fQM8nf45yUKzZsLLbdxho6KYjGn0klLMrUPzX6n7hQZpNxNHFBH/l5
ByPuMonAJePq1l3kyV7UDaNx4lVa64bChH8vqQyCuyutdvv7THHporvPnzjWjRsg
H84CQneLFpk2m4Y0eceAWszMNoztLTGo0mCRky1CpUydbssm8F06Ok1ckmGJ6r+0
fDVCZ4nc3LdbCixSyg/9m2JtIKb7WErF4DYSw3xPV1UVO2cb6H0Q9iTboGP9Q/VX
0kkUtZ68EhaU/Wg+KiLUW44RJ4PAUPEyKQk+LJuwo64pqhsx1wVSR0N8thR6UpGe
GBa6Cey5SfjleWmaF57cyM8PcfEoJbpx/3PMcqRI2KjU5HW5UquluX5RHDIJUaxu
m1sRQvQqts3ozDPmRECqPlbVg1ikaG05+9v2wA03DBC5iP2LNpDW+KL5ZHjDQNg1
MTa3+Mmh4gybd89X6A+ePxM3y9iOKtG+JiUbvMmdB4mexJ6e67Aq0DZw9q0iCXS3
MdJ0B2t3LAMs+lo4I4c00McCRoFCqfzJNwMme2DS7XbW3K5kGvwci+WFXu2KSftS
KqmcE1n7k+Li9vMMK/26/z4BLxeBMSFM5RdXLY0y6F1EXY4XSBZJiovHBiZhNR4i
KcBVxasmTjNFE6CVvL+IIrU6VUY6Zcj20Sn3a0AkLEK6A5FDjKiknh4L+kyXk+wG
i4QM2mX6WKLEJzjN3JBH/9Bdsp3eR9b+MpHR+aeGzALYu+ZL6/uKpbS7zmBNxx/c
KsSZBBTrGRJ8FBtkN1nuJIvUfI129M6tb3KZux8D/udJ89AfykJyl/1JfaCGQpLk
UWuLyqBK4fBHBXEh6pvBtczl4eG6NCD/8eBgdl3EQtkNtgvLSyYHOF8VC1Kpown7
17QG+ohiNcn3WIyKXwSxkMi+COHXUYpQXVILbS1y27hmRjS1Oc573fiJOMezAk05
lQ72jja10pHROtc3ZKah17vMR7bYh1Oe9gGwQZLS4ZoheVRZE4Tf2nGQ7v1py7wu
IatX/1sw73Fo24fsocDayptWVNbxTJynYb0Lsa+09Sro+YObLNO7TX67X1GYZQ/H
dQAuStzXA1UDMuTCYrJVhFoEeD8DMY9Nss398CUzoH5NrpyujqvKcjwQQ7NGXD8J
v5g59cE3V2sL3Oc3mneVu32EewBztFMeyRpgxtIo743wBG6+MtYEWT5L9RGq170W
5NeLL+Wt3LJDAFkGQAgiioLf21sShBxB9el84/8udgTjthCoyKpz+64v3w2RiTyG
uDLzFxpD5DsJxSjj0sH+b0l7Ya1NiUGPtJ+dD9T05yax3zKJvAhlTtLmrWa0+SdA
DWl8Dg527UhON78VUPY8+Fyj50qI0IUfveoLgHFZkrxr4CwcNB1pmN7m7zvMtrSP
TNOrFHeG3f1cQhkYGPy+wrvKblzbYfx/sTMgwvmJwFq2s6gMUmE0E1lUhQsBjwRX
Yc/CRNpzFZEhGTVliFUW6QI204N3L8XFG82JyydESIu0o6VrfWFLVqEW1n2DcR0a
bPMqIHkubbm5vr2ux/0MlPvYmLKJY4xUAP6ZjePn1aV06ucxYVeMPX5cykwY3Odo
aqV6jX5tyRLwM/SzsnQmqRGMODadlSyz0rzZxrINNUM9K8/gXopAgzd8Lructwm5
Rk2alVowzXmCsfXNV2PQXp5DR4vhy/pJZbKNOqJcU/pp4TtfAcsyB1uHfH71V50f
I4yXc5DPai29Y0Zf7+dzY4M19u56/jGRH+tnK43Bd6KCFnmJV9eS84eh0yvisxDh
0czpdD/mNdLEzYMpccEf3BRYSFu0nOgcwyevf8REb2hBRz1/uMFxCLKlXLEZuHXy
VSHwNv4kn+POfJfKRMui72AmWyCcTl1z4/agL5cVQ0Pw214+RLYUWo8VcBynDjnW
s/W2Wzqk1z3NRI04Q1/9NnyAxvvcwIozQKk9ZOxsN0PyM0uJg362nsubh+5cLoS9
A51SFY1L+iizo00q50yh4/ImcztFmV60sWA+yLxCHVJdUb8nYNadLZXWm4SgXiUS
56axokfwUq79hfKgBSQUoz3xAPGP7/8XkIbvubYuEYvA2R4QbiT6Nnbm5uHEqlX9
O1EOlG/h2g0DzK1s789OhG277C9lTb626ZQNFhMElR8pMlqzM1qzUThfs7nNTqnB
DW4Gf3dT7nu4hv/jbAKNwJXkRIGOeyC8rNz7kD77AupB13ZzBzTp+EFaLMAhSCCo
rnExFO/EXJp+24DrXMkSplvyYxPCwh95t897gH22DBONsUAMXi/OFTXUm5DhZ51T
DppC9c0y+P3hInkVnGr4UpHInlpEsWnm5nymS12Ahyn4jlZzAlEPciBne3DlCX7M
/u9aFDAvuleQ6EIvNfXKT2gr8tYgZRVn3Ao/qSuODjD6zC7bfcA8RLlz8BgcvVyg
tP3x3PNagUFCHD8upaV8VmL27vWbnxT0Emy/nBZgdGcql1qipCHGt9dfJDgdntE2
TNVTZHRpU91pzBxFm73uWYJEqCqO/99w0UcszY29Ti78CLnQhu26fFKxDPFtAM8I
20QtCyueNr3rOdEwm7x0nLgIEsXg1/b7tNtSGnrRhqMdbRpciCK4tGXwLpSj2sQd
E9Hx/WtlmflgPHBW+2pMEnEpGfgnqGQxoVQidz/imJI7c/rjPM/xOwA+bAJu6RQ1
3kuzB3ZDTTguDeF1evAPVL+1UCLubsK3phw5Pr98UYZ4Lk6fY6P8XQYYBJ+iWwi2
kI/lrIwiS01K3l8FM4m65A5DJJyq+S26BEOebjbO/fMAVazYnDO20bb9UqnF/EXk
C2DHy/hjQ2vjuEUaNIgzRkbWWHp+L4T07kyKvdq2U8ifSakPjQiFPZdINg3+vh27
3ygvwSFLvWBHljpV5ciO0soj5sxepGVOAnlXa0OyK2zmCYfPSwhOjDLgrQTPHe1L
gf40Lj3C/OAguUATRHzPBByZAQsuINE9sHPDJ3GjzOZ4BR5IbWyb/GWiLzg57myR
7JFVZfZv6yrZvlbVOk74Z4J/skot+iEN2QO0Wmv43FfFrfKuz2ZBhtNS7sgkwlJM
1nzQeNFniAwjZgsDvzv9ZF0N6mvm6s1RB2D+OK7H61qy78OL2zOx95sNNBjqf5pg
0AHqsk0HwOUFlbpFwuZnIBg8ONTHIFSfRamI6DSRCJ2Zsnq8D6tHE/YsYH6z821M
Uls1qKfP6kBpfVoXG1bEhu3sk3Bg/RWYvei5Bss8xsJjBLzDqSvdlX+1gKuDuKs6
quDtG1Sflt2uBw6G5l/hl9Cm/uPrTqp1lokq91hqLh+jeJyZIXs4jIxKfv9ANdAd
P+DEUP8GBdYfbinwtjBc09XpY2hw1+YfhM1eVjnVqdInKgYVQkx2HjqyRVj+1Ju3
bAlw16ythGTCf+sZXWIP4uJgKb4lcge6httb6KDWpPHGEql03VEUsvHDvIdfbzCZ
RWy72G4my8zn+NCKsQewUjDLn+mTGxZybmh4+U7B2iX4xzctLCXNRXxIMFACWRhx
b2oL1OCBa/uoAl2eH60t+o/82gOF2wX9d6jBQ3cZhbzcFtHN1XkL2JFJhRsOpNvD
YYiGojjyMrpyjpDwlAfHBQqF7tFRkcyPoi4r0d9m8qnZKfK6VoSQjMn+zcFVD5j8
46fIE+Z9d3rp34uwrdZ7nj3BVIZcgxtV3UhkyzFhtzymiVPqnuEcsdTR+T6t0Mk0
q0dcKV392gZFdOPwoJQBzDK2cl4eGSYFzX0xlfrb5Pnc//Q27dxTWKXgnTe5X5B3
zcFVXMMHPcfM4OEholUQpHtg4ARKhro9io6WW4TohKUAUXJK0lwDiG9BW8MjkWuY
TSjSRKntS3a1E2DPnOPaaPsA+gA/wq8ClY0WB9UIMPrBVGwbGNUKMNaELm2vRTsC
3ShAiatSyjriipCsP31udeVZIXEdTL9Mlg2G2d7cRGL3eNF47+qhUU33jEDQJsUc
fj9lV2p8RsTcIqD8kHREljQlNNgjUnNoVIgUGHk1QNRTIeZ82wIyzBhuGaB3gCM3
v663EBbcWqRLLiMDmp0W08MK5Iwt25C6NAfYtNmeusur3J4zTFhKFcOHi57qyNUj
zrjClE7Db6czSMOdIw87XK8AbnJ5P5RrkMeWE2ITv6lY2M1l9jvIPwk1s1RRlHPW
htPpV9cXqiYNM5lHy0p6//uTjLiqCiOdcRMuz8ou1wmdW2l7fnxz3/rUGKwCi8Ju
PTADgvrqC/SvwcX29bAGmyKLH6B9qGcNGFbzX0mCdgpO7Z5wBUFRj8K/mzuS/AY2
eAB7SlpoYzwITfbI/va8Akk7cZuIi3RJXfJYOenxHwe+DGK0nKTZ930UHGGrhlIO
oGf+8g3VjTrSv9Smb2LHFx7WJnM9Nkock3RgsIrDIOj/64yvvUYTDs7mUlPXpdFo
EPkthJFcpL6EKdUzyWg+w+4cXrloHApgyyfDYRBS/Xx2zkQkEi+Jhx/i4Of8F3e5
4TsY5jWhG6vyIGQdybhJXIPRzNHw3YR/dWsM5A3WWY7pmgCZ+bWNcFJe4q9TgMUv
Ya1lfE8uv3BNWpKAwVtvgVfVkihOOXZaTCh5hD4U5jY3/pqToJixqJfiaVbxLTt+
LHCx5oxZqs/m1Lzh73LS3B2LMxoGt/0/Qf8q7pg5jORfOIonxIrW9hXfZBsPuYeX
0opdCAs1LJT5QNw1sep5GzXDGZSXhG6Q4ZVa2krbo8kA/bzxng+w3Z54dR2EUWQ7
cUsXun6/iwqrS2JYphmgZ6WcZZSuALn3wZQTU+PygIsqAbTOoBj8y1Txj5zRGv7y
3RvQQ2GInON9QWVv8bzc31jFjmEET3YKbBDzMz/epbeAVkWBnUKQeJMYqCj1huJN
z2a+shhrTxLkKwXA5mr9TbWC/N207/yRGIT7sKwC25a1du4muhXBU0EJL55FPPsb
IihWYdaOVHHFQ8ugY2E94Tsw8F5mF6/HTG9Y0OditOuCuO5ZZ1keI8GUWdXInXpG
WQTMjwhK3d/V8YmJoSVpZXZoeWd9zntxG2GcKONtmi6BM76wBDvNL000HSS4vxkC
BeaN++mfheZLFEpz6SWRazIlibpryJjwgzIbofpeTZPwxlgqVI5kW/FAhVrRp+qb
lnl/xHAnqZc+oB9PCFFrLVBg7wxKaPvPwZ0zCECvDL4gucsfJKmbf0CHaKMY1rmN
9aJM+WyaPKQP+xBmBut2dL33JD7vbTkCBTTDCBP6MQq1xIeyU08lLD2fT/6gsQAa
w+OaGCZuuXyEGq46LsSs8zI+54K95NL4lOe07rBLKi/aSJSS32FYgf4HhPLPlC9y
vbzD17avuo8ixwKXmC6Wb0lugESsj3rx+AmuPiOFkBEGsK/zOiaNQEn5ELshO3hK
RGHxXHiIdZ8tmnaiW2+AJRL3X6/IfBGzDCiPA9Q3EoGG4XAPuk/F8My6AMRmTyMs
scrokyq3iKrqDpQril6JdlxCafSo+8S9rq4+fNCOrYg1kpgQDhQ4G2wlbDOwHjAX
hw7zLqmuoxpjvWbrb+xKAKCDWTkFlIpARAuq49RxeEQhPHNexj8Y2bc3tUPP5yGB
B5nJk3iEK87JK/bVBFiQMDP1bABWR50XFIrL6haM1FbsaAy1G9mNRavqfrgDPJY7
1n2mGIdsKI3xZbPJ6/xr/YH761/GtfQOOcuDtUeeLznw4bNsOeDgAczb/DxZrHNY
rQue0NK1C54jO6GotDMFKciowyRhCxo7IA5lOJyx/dQfpY/OxGHuN+xFBb3x0quP
LAJmsjPXf2nigUlU/voecCcNHyBaoeC07S7JOD91jUnca0BFJcLw/zRP8kEHnyn0
Rd1YtselOKI+WcYKgQZFngxULdgaPwEKrOOUnV5KIMqZPHPk2slC20huNBttU4EB
aHD6nB7KNdQxG+4/12LIFGpXqPBtvvHcXyc5VYt8u3L+46f35XN8fxnClmfr2R1B
jw5EoGuLMglsbXjzVfHCVIxqrJvwr49rTyaTuYh+sJKf3BJO0jaiqASwNZO51E8x
X4sAXSIlbHiKJHiaTDMcCv+R3zU8OKpDPI/9vgiZLLO/y3li1dIIDe7b8Ss4Xc0n
4rAve0/s3yna+idHzIX30UDcUYvFqqx9NmIz7ENOEsvgZMCOK86/C4tK5j3NwWBK
8hJ3WsMPtxfswrI9f2YBshhbSzjSf1efNQZGoecG9sOoi2jiMXFXswbB0MHBBC9u
JvIg4RUe0s6pgUylCSgi3pKwJMMVEQpR1oJt8C9GvD6JjnPSjNoiDDFGs0x8g+pU
mg8eoO/fd3hKjjSt6QuofBXHx66nHccnFJMF6IsGeAP4wLv474SCboPYUuCYGfsA
7W5BXvzpoJzpN2l9Y91CSIJooxmoGqbHuVi43XUHkPg1GNWXZPg2I5G31jR85Jlv
zAww3ejNLTEVwkNdbNSNEduDDRjBTg2He1wW67JzLyseNzptspKRfSxCS7roI9Ox
eebQLe31PvIIbxjIMy05kvXSOb5DWQzZamdPZIV/hbSemtTEeO5onDFvRO7NXnpn
/wmYvSPFr47ktgne8AvIgi0ztEwfXvb+gOSzOA7QuXw7Kxm0nqXUOWXO1UWu2pDR
Q+ZrVew1c+rtN4+x3ekH351QGEB0+ff3TAakO2Ta1zE3J2Sw+TzCe6Oh5mkFbTh3
Q/EAfreUOwItJAO+mRINSmxeAK4nvLuRUfZFIbE6jTTA5hw0f1nZnA/zqldatLDI
YkWfObE02A4VLWS5FKU1ZhAFKlJHg1pkfGH57VvMBQLJp18K49N7ZdshB81TCBUN
5lLGHSG1gEtzEvtaTJsijnm3q9Xt6DVxZE9R6+yjvX5VUQsZLP/k8vMO6Oaygwmf
BoMoKx1GeNGRpvPaIBISHmgFrErKlXz6ljMiIDvkcMmfzYNC0uBouv8ylVEV/AX+
bwvTTcwfDK7N2dX1WIR1cUGKhFAqBJpCv6Rn2v0AH/WtBdPp3g/D3csVeVIiu95U
nXqO6EXJD5BPdK5mhZTKg/7DuwuxN6e96AxH2cYbXCVR89zS2MZeYQ8QGPC0Iu78
5PtEuyqBbbeMOIH7npTcDNjrclKJqe9G6t1RQ+rTNON5dbE0WM2Xoz5Ua5uGiYWf
B6+54DuqgR+IvmnPZh+1kQek+fpSGfIRx5AxLqJXW/Qa4JeFygx1ysIruiVzVcbn
pc1YzE69wjcIxVKOrY7PoG12QDzntR1GL2jkf3dENzgEldeCXhs8eIa/NLg467c/
o+B19PfIRuzCRGNNwU8awb6X8fl7/i9QjAXpa4Wqa3fv5BBIYKB47Afz/IIxXCq3
9j6BwciDfuQyen3EItKm12Ztzk0d6v9VkM9XmyrPTFx5ktH8MUVK6chJbOyqg8Pt
7n3Xf9Fk5TdB1s1vc8mZ6rqKaRJ8r5PLB1BlrmljMzscaFYoEbdMkn7y3ym5E2gX
vYFuwhfqO+L+gjnglTz0d/mTd913ppKHFp4xK5UhohPervXz8+CpAlz8ivxOQnQi
Dpawiys1KhAPnDfR/MSlWv69A9D5iyJjUbFPcBIrnjr8Yy+8szHcqmut3snkbcLT
24fU6dpX5HpcyDBKUKhfL0zAlAZammU/gi137q76Kk2hN457Z3bh+L3uMy7WjcFE
RYsiUDhXmUA4iWHxEbWsnvx6MNXI90fxel69Hygs4l70xzmMqsdsY0EUHuAP1JG3
EazD4iH2TSdpi3wnUucZ+niNBt2zs9vu57fzEccTWGgcYxqETzWso2kDKlep6IGY
3Sq+2pIvMcPF8Dalc8NyrQgsCuoxckFi9zvp4anYRlWKuyoSDecV+iirNog8Orte
xln/FG8oqHhPpCAvMEj8TkfWzXnTclYYpcVBH89O9o090vOdqOEkwpBoPHTrGfgO
U2zfYM5Wp+voF4wEYLtxiIU627Oqk/h83bDo/T9jXn0KNARdOXrgI4l60gtm0D3G
CYKUOQzxSUnKl5a+milRHIamqZdnRQ4M/PtFj5Erso8QaacO35KRcuvvH9AoDOyG
lRMtKQGzOCtEfCYhARhAlfebn48FNe3kttinnNyuXnrdJnEZ3wNwYuQWExffGvKT
+o0e6Ssf6oJoPw2+or13OIZ/9TsyE2J46XHut/f6bQgktTbxvQJOIr+bKdOmrX05
yYyoLtK3Z7l0xgPLpvkQQ1J3PmgH4Z64wyOEuYmyFn7wjhNNyak/UKv8nTMAtF8w
RhB0NfeazMdbsWEdnemjAVpbZAmT+34pF19hmTQKtFdmcyGHAqsZiXnuLaY4PLDM
73TxFV+1O01uqTuGqqv7zrHNv2E30vPLSpJ4Gl/3DAYSAtHQPevHkV4C74zer5XG
exXzZY/ZGhjaFnpEfrHTIEt3wM1FTLnuTGGB6pQnBWsAQgaPlzQ+j1r9SQTmxmsS
srQklxBX+zhx1GQXKtxuMAv5eqEBtrHrsR2bs0F7w/ztN2C3iIp5NDeQ9v+qwHxL
rCbvplpU0kJ+emJsbG20qvJCaqFSbDc3xVB7hZMvjqUzYfslYlTye2E5NO0UMisF
hk35ZRm14j9FyN/lUX2O9lhMRk350eDOWZR7Rb5/go2WkpA5mse99u5mEsPT4yK8
kcPRduZqmHkQoODqxv/WAZ9KkRH5p64WawJOIzA3207if/i2y0QDYPl6awJArvHe
WvLh2zuIKM9sFsUv++DmXe8mu+/GkIQCuNpx7r4q7VwOwIQTko8cdN14pg2XtDv0
yCEUBO9kg4JWQoOxuxSzh88C6Q1cnjnTqXgbPFknuJA1gahjFycc7n7GGSi8ui6Y
ZKXiInU+LEpYp/4FT8DMrK0RhagMsjaTeBKudE6MuklenTyDfX0nxWggZaR6iDMQ
ON5IMYOe2vzE0zN9c4DIQLl8z0FuVHDMN0VVL9yoPsxI9mVS9uH4wLiamyE5R02R
5KDEAn3wIf7Rctg66DX3UC65qvb1y4/cz9Zo4qsE4v0p3nz+RaS2xqQzsDu0wMic
kNn0ktrMtAHzyRid0q+F1F9OQrHC5daFuyeHkB/kw47YLaVbpadvlsegWxg9t3PN
MTxJNz3H/68GEgFYonW+xeQj3OLd0hfcCLmCLwK6GtwZnu3qPImhb9ALoCGtlPOh
9PfkEWjcV7PrpSHsVFbgj8CVyAnvlS6Pml+FpTIQG68y9q8VcfnCXgEnvxRWTBkD
Gcv/VcKyxXv/dAVs5xfYUtQ1+AuWUpDkm4SgmAeY4ROJ6VGoni1KBsT2fPPK5c6K
sZp/uSDz0m2mB8I2Oedrd2L62SxTiMtERhpEDmcAS/eE+53tuXCm9HgPcCOHNDKb
Xt3Fs7PQEpZ9ygthdt6KM7v3A8CPjRDx0ZfzmyCMOkC9bMggPo12mFV+JLjAWsg7
s/AqOFwD7WN8khIcQkh7aBaZnrZG2ei2/C+ZIWqCw2aQQ4gn68oKZ+AURcFt0JXi
V/tb9crL8YaBtqECh6P4444DN4qEknkYW4phPRemVcqjFdnHcUat7zqX16gGZDpX
ah1v9DmY1K8JOa6WJaiFpCr6BgOlwFpfNBNgIZ78ihhNL3U6PBAAgUW1o14Rcedg
w4S4+310OyFusrGLDT9sZBIcgIBEkx5vrrASklrdQkg8XWam9xwWbf+KaKCjW3g+
DT35XguuWAXdoMTNTDH2UTL6bpKOQc9heeiK6BMqjNV2IEKuaR5EeNAkOf6yuHpG
4Dx0NtDeoyc/j2iKrlaoatyCulnD7sZ+700HjfLd6VJQAhXT5iMm1FCLJJjDTBsY
mQUoB5nY960YgKk8XTN00q/By4Q5/UESJPgLMYu3jjC1RZBoQJ5GarS7wjYMJ7rb
SQWj3kl2NZKAuRCxL/NakUQAsXtUORca/hu3kgeEVta91LFAdlUytBfJoqJdrph1
T4AAkr4X95ZdzjzLrnVC2/WKxtthFN8cz8I0JrVykcodODl/yRl1MNCsysf5k2qA
tFJfBBoPN0JoqqtD5o5u6EhTmjYt9Z2+1SN+jr8gHkYuDdtIJbaMjvLIsJuAcCfT
RefbKafRQ/XnNCucYM2442BPHvVBAKx61UFE/1/M4mpXDqL/EBZZglU5DrlQY6VV
HnV9FTTruXWV9xQctQdmEV34qCTWE7c6WfKz5vg8emymZPsiaYCil1kcXZK+uwtd
gUURrP8WXC36iihsID7SJRLpu6U9k0wCIpgYdq0ZG/H3gcQ9h+Q3K2gHXNKLjC+l
4cu+RsI/9CDF+HUsk42X5DZ5t4MFTlIDaAs3gzMB4CFLRpKhBfNQ/GVwoJqnjviM
kyTjy1cLYcsX/jbOkNQfFQdHViKGvoc9ejKhkgWXSVRn3ZzyC4ZKfJkEYoDVL4MZ
byAWC8rzy8qRraPdbHtwcBTufaEwDKrncqjdmhdQqBIh380HvUntpWr9/T2bclLB
75/QPkL26xH+CNxg4r3Ozf8wXuP/AVL+88PMoP9TmklTjUS3+S9hvcN7P4gi53XW
gehzSi0kvhhFWySBErgRbtV95SizwzKulTOOZqfdu9oaL4lnl8J7jLnjJ2+MqV3A
nt392NRkaAG9b0QdtXUSrGK4gpMd8uTJpSbKg8Oiw9hWTS92vt/Hb3iVegCN7Pg+
n7Vc8QIgH3To2ZZuohhomUjakNKJAHySdp0HIGHpbSUQYplJnzajBkcFjjNSsD7i
d+sqypVnpoF2+Owbmp/JCOTt0YX5zPMEY0XSmbUyrbKv/skwlnFBtid/uSdEwSa/
blb6K3PFE0N2lsg+1TnsKqnOpW231TktwkFjemO5sxWZBA+ZGM3I9djJuYCyqOI9
utQyvoQVYWaH17HjYlqV5o0nkUVbDmHK7uRNCI/8AMrCiCfJR2YzHetMtDavo6P/
Gwal1NK/G0rbRL1Qsg2lexfDExie3BAyt+urB/jwuE4ibxQh3iVoSGo6Cp9xMmAN
HvRWiIOXpAewllD/hq4R9caN5ppOo3jmMIGQUPlhlrR3FufYF6TbblrZyE+idh7N
e7gbP6Xa5EHOgtu83FvU8YRUPucrhHr48D0Eev+DqgZIj5SWlQSLQdvKX85jHpi6
Gq/18VHoxLY8wqc3wiFdZHPnK0UHBI8HK0madJBJce1SoUmEDVYzLOAUxrX/59Og
jaGVqH6GmLanBeqHuWzApXwQP119aV4ISQkoQj5ZwmpMoXIa/Q6LV0Nu6q5S9O/e
46wYu/xj2FufipqOyYcP9ZqzZmDtFIq1m3xxa1hBrNzKcJtM6C6yvUimg1JPM2xe
aU9tBd7SvncAz0ve/JJ7HH0rvkyyeOhAukxV1O2ZFA6HfRP246M9j9mbvysQQPNp
kWNxcU9k+lu9TKni5aqzaB4ypP8HN0DNAJDWBy1vOfGj1re1YItVia8Fjn7CeEBp
TxZurnlM8Zo0vltTVwBzBsBY+zWu/g7NSRXJSXcrjAHML2K6lvfhbIWYimWkJo7W
a2xTB8iO2lvABQ7w3oDkj9rsch0ZjwKl5NIac0b5vX8p4kIizVKIsqDfiAihyiV/
dg8LNsFO6Ns9n/xJy52Z9NgGc21df1SeBQOSFzoBhsf/yvUVfdZU7UqZIzBjoVVj
jvAbXJiP/9IoyhT1beeFqMv07kezr5RFqbsZ80LVniFjjPnr5ZGkLS6yNsOe/8/0
bhAnw99IY+LEETEI9hhuuqDdDMCTjohMOrAMy43E1OU2Cr3jMRd1LJt8WMhMjFQr
xZI+1oR8JF34W5l1+QiP9nh6HMCm484Z58aPfmT6sSi9mynxLtfg2nNYdVCqm0LY
HsuvbWVHltDlzXGXYoxvubH+5/QvN7C4wJHxYXx/mOo3hL65wIfGc9360kIj/ady
eWGspa0DH/sTNvG5Uno2j/v8O5L88fsUg56w+OSaLxWqSK05bcrTpxgMdvxiL42+
t4su5nTB+bPhwrdx9bIKSBe7H/AkoBXNEk1Skv6mTY7+Sf+W3THVb8D2FMquV8BP
CSzkyr0RpZk/EbWJtbIm4Yls7fs95KljB4jdmueEk8qPSGvhQVPBUNc6Vhhv/qts
8iEDtzYNvvKQ2E2i5uOnEQly2QJPNIFY48BaUIISFxn78L6vPsn3ZIr4vglfMums
kxjmFP3EiPQqWMksNg7Cs0P6LooCojlCqErvqzbU0mItx91iWdmf1Ug9UtQpfAc4
m4getOx5FIC0i3AGRokrWAJeD69uCo8DX60AFyP5+u6QDeJmW6aMOL6ENJzYiqQn
0OKxvoz+o1w57F5DsPRu+D9cEANutr9C/4mGCsjphxpESv2NWpo+CZ6PnyCFC8q7
5BtWhgLLbDZyOuPkU3O19yvp/CB3gSk5fJE3LDFg2rOTzZcYMnz+Q60rNfJXzH4D
XMFtOe8/zFrRWij/PxkvkL3dF1v/rTr6+Km4s+1FQLFiXVHwpuOvSBU3pvU1FU09
ziFX6ifh39RFzGd968wnb5OcYZ06O4kZs0h8vGfmRXVsArhSwnslLCKwAXUciONx
VAaSb7d6FHD/U4Y/DW7YxXxTksCmvQoOaucDZ9nZHf4PKeuRYUW7ZbOj12mhqmy8
Q6aOVlticVvkYdy42GOnNLCV3slSMe4l0uqHs0MXnaLmVNFHfImCUyLRmYwuc2yt
C4opiWseZUisL/aklBrCI813JfcCBeI0fXouE7Xqtimsj9YtYeeqsp63MjKe143u
vuk8D5jU/GfDxsPNyCCW+LzBWf7r6hNvxkiiB1ufe+9KVPYYwjbEURT37KDJMQ+a
vOti/vqVpLu+yffpSAcg9jcC4Iq6rGVsN8jjLBYei8trxogcmv1gsP5qs0SpuLwA
yEXwF2rNhhw9ZQ89qINgwF/Uwfou9eY4jBJjKVPJmph+MxV6thQH3lFurYvQotIV
2PwXq386XAFTX2mpKiTJuyeKGVjjSpU1bzzu5YuooGyNAwssJePhdl2kc7lmEJGg
feJ4N0GhGn+xPYuItLt+3fak1CwUXrshtiX7VlB1TbfKAPz5d7NrTx2IIjO1bfRr
GDQQYtuaPahSvTc6BKTRMzKffe6rUjEwfzjLKXReI711Uj5VEJBsQ02ozTZvx81U
N8hNVvHbPRn4aiAc6PX2bO9wGrI7kI0cKF1hEBPcrC3IlgHurOqBEpCLkZjMTZvP
Kxp61VosMvH06LKL2uutc/QrsJIYtRLZ0gMw7VJbOhb2nbQppNLmj+5NlKSXcY91
FDC0MRvA65F8SLY6kWn9rGcZVao9Vszc1EZY1+k51AixnSPiKVG4J8WRN/HQl5Cx
gmUjcVzsRINy40E0ajS7Sn0iiKLCW3ZwV+1HcskQBAoq/BYEm3rIy3FGVB8o4YyQ
LpzNM+4Jwcm9dsq07GwLD+QcLojjeRIKExhQmOnpXy3YwOTIfqR8LWbY9IRzM8i8
lw/va9vv2SYRII90qhnthw==
`protect end_protected