`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 7632 )
`protect data_block
XAYzcToIY1VIPqVIYOouMwaXR6+iabrWSAEf0x/eFj8GuEaEd0S1cjNRhN4pe3ey
dScutQVB7r/7WEWDYSh8KlQIia3LXI2SBE8xjX/tk5LCgNzhno9H5DapHBuHJsgO
EulfYGnLpOIT24L07xg5PzKrc2ymrZ4gjUqPTfBF0Ss3PszGYcsO3f0HYOd0pQpJ
14QMNQMknx/+sYdZc0mXkvRITU3k6j1v+0IcI/TlDRCCo7x0WWFJEHVkDfkFmDWu
O91lwapitj/X+drib++nhEaXpHzcdZ0Znuq89oOjwBl43r5OlC1CMddPPS0SRuHo
pwhENX2PiywCpAKBoNFLEo9R+UZb+Yfn9Um4qxTNU3fLSYmbBIbe8XQGZ9FBu7NH
BzJNqEbckUgj3Z1QqfE/8KRlUndxs7sMOtNhSJz9QbxFy948cicmT+hOMZwg6c7Y
noekm2K4aE9ZFY1C/G3LhTc9MfWptTaFV9yFcSn/9cCINOz9La6G0YdYCbiCSDd9
5R+TS6yw8PHjetKdvxPlWoHDy91ZoxFRk4BeqIJCEVKGsuu71YlBSN3BtOdpOKVr
NVfTxztXokpWXKncf7wKp1fA/8iBs1heeIYYOSVzaSXXHlgNigBvQHNdet8tUlbD
89NCYu1MuPTuSNxGcppAPTl776/Bzu3SOIp0jhGqg7yT5/YHd6GXFy4hmYr07gz/
9Yj+ogx5H1PvXWTiYCJjZp+x2NSqS6Zp492g5S4e/SSdiyYmy97S2PhtxR/QItp5
Iv4cR7bh0wWgnHCzGGvrKlTwWTzEZq+Ocd5Zv+ssgEeY7bKB7X/o7i0Wx0KkJ5KK
NEoN7UuNGC5bTsCMMTC9B1i4ZjtI6XFrQKyZECf1RauyBQ06bV5dPC9IjehgmmeI
oyz4FDXB+1hEICBK/eZC25bopJvMMtyB3AP4V+umQ5ZBZdmKShiMqIuWPR+ojQbx
CFGZ4VCkKff3EHK7R8JkHy6ZC2gC8SBZjv5cwswPt54wc2nCv8qw44ml20QMZmCH
eflCveJAHlXeyEkhMaZBTIKyfjZOhO1YEzgv+rwccNoL8yGT3h4QHioy/DeqO29d
l+Y87OkAm+3GcMkVOv4UZnNopaOyBeGCXACSbm2O3d/cImfp0wHSCmHRQuxysmmj
PaWuZ+vvzLnTcAm7LV1CYu6CHj+zTks8apGfz5pvpbAcHHDluYOlifL5dnCuATSq
8gAMyL7tuSExtL2n1SieSw0m8kg3AtGXKszv4jUn7wxIopwIgR8qih2m81RYcWVZ
lpUj1am5v9yGlQLxaq5y5Ev3lvzYiEIPFGaa+vjVuCDMtlqdn6dUr8iPAiOwMAbw
A2ariOov9tkJCFxp96zMiBdE9Rv7bU6AipUC7LhU3/5ufR8d/5vFXpJF8fTnqrsc
HuHxdh0hVapj0fuKDM9GwDyUPUWiQqdWEiF9GOKabZWS7GOr+2OIIo/lkWCNg+cv
8NjLpEXpzu5SZBidla+yzlZ+zM0PdO7RHcX44mXdVcaSwCofNnAL2AaGalfbRJx3
UF9kECooFAXxxXJr03sWZijPQhxlqK0rGht3KAQtI1xWucZk/p9rXBFyoH7FRSXd
QFqLcJxXhI5zEPzaKgksWxZ22gIiKQk9QRy11Nt5KG+PnZ4CQ5wWlvqMYVGcENfk
WI/G+VFH+ATLc9t2XljhPzK2abU7UAHUwK+mivuKeQrmkqpr1Obnd5vfaEskhO4V
ruTHznTgEkNdzbAw8ghxWKjl2NhTGaQfs25te8/AjDdsxjKKYC2uIV+PTAi1INPT
gXQK5NADhQ0CwWOke7QsawCfGCq3NGpJH6VcC0H/tmq5umQAr1IAvGUB0njFIGc3
t6seGhF9h6rbfDRa/tm8XnR2P5cLedu0wEl4SMmzOga3M56zM7kiRGAM/GQQZy4w
t4QJQj9tGaRSKNgpo+liAutLwXXPsFVDODEf/8O9a67NEdTUAum7MpwFO+BrfgK+
4X/mVmy4PTy81/0Ht1f2R+D6XVbP8UgiByoi4BPcEIGiqdHXvs0tdfToFkx1FZV8
4iqIf4Z2FCPW/ZzN/cHIPi8U7+4UxfeesmeLprUgKPeWBV20lESp7JC+kGZ/G215
ODyEvrezkySnok79dwsegC4iv3HI2uSV9VpYRfmfwIiYMLZd4S82ZMWV6rMZZXIE
om+xwvZ7fF6TTWVHI3S8OPyr8jOz6aYt66vXwM+PeKNu3xf2pcgcrluqJicTmi+M
aQXYc8cA44XH013YHmaACFq9VCloC61C/qqMIWvU4oEARRMHwNEfPTI7hv2cfDmv
+gqCiqQMeLvui7ctRknTZiliLdh6sfWdzfHxRrFuw84K5wYOKYx/RXJRGU9V+fBf
9Se+0W9CYeEfSZKnBY3ku+41pfqmKCoyS1wIJ0HXFzteTGnXGLLu3GmTwEyENNk/
ZLt92wMcCtjrCEK2oy1n5XyGbubTBENYfGiMyK5rkR11inXtxlSiU3C0qrmRRdlI
Y+K/YvDAlfFT96g6Bsm3YvxCLbEgVDhRUijIIzQnJwdiVukRn1u4q2qgGnVVBR4D
TJ+aYzAj226aFxxepIti4B+alOZqw6b5IEpP5BNmIu1IJkhZg7GzEFQkYQObYdoh
eE99vPHtPizOOj1EYsWAd7hSU0p4hAyjJCCXmZXAyJTERIDXCRdJyZpVf8ikp0Z1
FSFpWKfSrxoVSNPW+vbLgsWaIhx5xEXwsmjk/Zrb2IytkrnF28aRzxZSQOLG7Txt
G9vntNyMFQC0ljcEOsLoskXGMYrFzL/G7QGDiU3vNT7v2vGRUfV0bsZFxq2S2c6l
IGdjjSl1EU4rvhadNdXW3Od7KqZTIvU0HaHv+3vIlHZWffLHKz88eiFqqwNlabWD
3CkRVg2haEBKT4gr6pheGPJBwscB4K0eh8dhKum+i0Typ2rettrhCDGN5WiOu47j
tLURzUAq3nejm5S3h+grLXDC3OuQTYdZyVXnvBx1E9005n5eRGS6y+D1C1sTovbe
C4d1s5+6DfmVnPRyI/aCcLtTYlOdE2/DnkerC/+jKfxczwoBcbX/x5rOoAyfftIN
XfY7bzXTCIhgZhMzzqKS4sjNUVKXeV/qGgSGK+dfnqg/tkicDmcGnLGH0beJN415
HlcmJsYEte0AdYMDWU8gREtWCoId/k8rZG1+HsD6+jOWDNRvfhKj+ByQuSJcbiHF
CTba3Z18FmtFPHo3dkm5+ZQXVEks5h0EqFEOvq02CCluc86mVbQs1aDxQ5ngfCtR
6x+Vrht6OrO/NY2obmssmLlpChZ7kSCDcMK1tbsX63Tzl/IXjdAN+AVhixywfJRE
yGPbR9L1siIu2fhkI49xtIOsov6uG4RndAuOVQ8qHWp8H3qIgkQJN4rmOr13tBr6
ASIwGWt5hKM0Owv245bTg8c227qFKaaDJj6WLLS5a9ZUeJePDvyNIeHkgMHNHm/y
Fdzkc3yAfIkklTMdp+lWzPEt1EiSWTOA6IPaMmYzOhRqnCukelQEUutctU0ngrob
QH7E6btGbwAQw8s9B7X4dg3GTj94AZaPtyhnnNn66kVjQK8Fzc0xTy1aHwdSoOVs
yA5dOY/cduPTc4T03x6r3mLS6vGdlAu4fkedkM2nWO4OWZP56DnEqY4UljLCp4Nw
8U2bgGVqdfcSG+nJeFZxvOYA9JbgN920nl05bDIUCRrhQ8u78+aTjVbk5C6YYG60
fyNlzn6NHf1MIXDN7U8fHaB8SFtOVX3g9ECA0F+0psya/ix9i1ciK42Ne5ST274B
D2UL2jX48rN7JZG9U2f8zIiapC8peyNkd18BV8l2PzOp4z1Vn2Jx3cUefrLrsHDW
hBczR/5u0HKZE7iC8Z82JuMJEkK9xMF0R7Ypq3HJvDp7F9KgwUL6JvfwYLV3rZWl
J2mhCnJZuR4NYMT4jAZf5JN+o4BVnM6LNHQJhefhySByul/4G2vcVfaeQonNO3lp
+lHupQ4cHvVLQQXF6VRJ0PIPux1UbBdUqa5u6oM3Cum77lJ8UMTFNWQpu17g8FS4
1TXnv2n4821Y+MZr28Eonx+siNmNdSkVZKkSI5SQd0Pa38TD48kOEJCi86V+Y/70
f4K6uuzZ9q2j5m2KxTw9XikOf+HGkVVx3LZe9Iir5UBb/Bgg3vo6pCr75O9D8f3W
89d5U4S4LpWWckC0m6Qa58i4YPCHuUSyiP2t6v5ore6dIlGhaewlpSApPBlzdcFB
O8VJ5/1fUbZe7xvoR7upo71BLAgGx9rIo4k+GZrb1LTSY8Jq6/1qtxhVLJO1ZXyq
z4eNfTRnEojgM15trUqtoXoGHrjcCxBd6/Z/VHW72yIKugc+qA8m6Cfa988H+G8x
eH+uGpDtce7ygUwakJiMEXT7IPwbRkr2OlXWSb9F/6d9sAoVRwcxVuV7KgFcOCCE
VTDjUnTsXRVY3zzClxYLtcf+fNPdNpAtIlSVvdSdchhRwFfQaHDUJfdOrT/KSuuD
lnxVy4yDXImwU6q/hSQYHKUqOsdifMC2/2cChPeezVUo2hmIotK/mgS1o/gkm269
/VyN5xqRlWXy0XuFsYDFoeGSZUvIhYGq8MnYTdCYw3MkRyZExwTfU7siwfw+2IX3
bJGSknz3G0+GQlfb8i7Qwhh4myezMMZ7C5WTVyLMbuBuerSBFYN2FDj3ZVwNHvUW
5x+zQKN7uNijO+MMqSaPsDbnJa1E3+NsaHXxIwHTY/NcirCIU3od7BmFdzYFPuUD
bYsgAMxo3wyiVSjvsFkUsvmJuqwX0+aSHqlqeMfq5gzXcC+nBAexVL8v9Mjuv6AT
Uvs0Ce83Dy7fvPRFWy58nuCbFldwQpcqLjsTV3tJWxi/cv3gWr+s/SkBmW1PqUfp
V+Rlu9JPS78W42U1ApFdI/21Bo/F9jzWpsP9uMXIePgoWaTEY4rp2vFn81e3K6GR
eKhda9/W4N21w0kiE2203deJXfCFqoMRzweS2fXZYs0TF9kU3EAJK+DMMqAuAjRE
OuITMiLCtVEpWSYPBej82eK7WxBQRj5bs2iitFFBV1VSke4jmYMtUns9N3SnsomM
xB6sYjCyIwOZGt0hb75nlMQ+tQyQMqXuSMHluaCVOj8fOqhmm47ydPGWYMiNhK+F
ybUOHMc+5XSIg5ZxaRecAFmlGu/orPRtEJsRgnEXVhxZvWOC94dhsV9fOr4olBA+
Gw4wNgY2CIpnul6DRh23u4d+DdVvDGOCqoT0DrRU6nqCqyOpVsaymqyLHlV0QEmS
eTLm3Rdd/4vaJ2L/NNRikKFYmgsWelYH7WBp/jInmplDj6rfw/oZOd9U08ktvZqk
vgPxE99OzcQUzoOCAf6O2HPHNjuhZxGfOLKPwzvAL3vYiWTn/OlN04Zy5zNRnRJZ
KX38pZ07KdZGMw1uOge26F6h9wMY9r1ugUd2nus3oQ8GM9FRx7SYe78i0BL0XVqW
xk6GtkjIdHSNKIPUDzRjZzLOLeqn1UtTPdQtBCu50Bkb/c1LBV4WafX1/2UWFVrw
utl1z2zSj/brE5Gtp3DfwOGBkFm4Wzs/omeCVMym2gH0TLjsraC6vfomfBD402xW
4pA+stOUiJcS4jLMYbD/ChXNY4JLnL4pmDCU9ylq6N5g70AHWS9eGCPzD5oMNkyE
jWjCxW8aStKLpPZKLYAOJFhf0Tjaxrc7C5fJlk0ePKpL9BzPnwAJUubJcySOpxJT
R7GckWYjSasFx81QiVihEFc0ZPGvNg1jc+JkzQXyawM0TTAAz19L/hKEudiVsz8s
YIzoFw/ChWqNdS0JwjkD30b1/r6vTpXOga244cSuY99IoXOTyilrEQubJUi7Emux
ndGXgInFqcOPvpFPLT43l88okKZ3IAuAhHnivia1+LYKbn/FtV0tuJBqfMWRGVLP
Zm37hyUabqKt+SLWVgfaH9YzDlFI2izSIUlBqF0MgZvqjpcHvH1duiAuxAZ5yOJl
6e/7jB0B+fm8m45CV3LbAnChX/TVkGmbGdAZ2sbk1M8kWMLiof/7ONhJgYFWl+N7
7edfst7RJpI4mW7FjoYrCFs3fyglcrcyShN8EAMTEdoXFIibXX4mP6aEVfhMPTPw
sI+m0wQb0+zzKGKmCYFkPhoi6UWt4JqzbiAT+6w5tkyKb7mz9JJL5kRrsRLJZf0W
YuKGcAdlSL6mkdbui70jBsBGjhhQ/QyZ33SPNARnmyESZu+bhdDs03A6A2k4imwS
U5otYRuSzrHlrP7ukrPCqmcWeCoPbHVCKIZwGHM2YM7mLn5cgSoHNWv6zSsIrtcu
cMk5G/fu0LVATQFXMb6wSsK9LuVZQrcVKRViZPSgHsXqZ83SBA3mgEJAimLN789h
7OUSzL+eSf46O2FZaEUw7z12ivBYdoyx6uAKCvAwo0xYC3RrAEQ/V0/q3Ne06QLG
bSJFiCIJb8ILsCh29wkznrYJ89D6iJwxinpKE9+QRisUfREjN+nJuGq9KZWAMlAb
fJm+ZUvP4DaK8mF3vAZOrbl2i54ONuHJl/fo7p/kJoL28XW/NHPB5YaMP9msPJVW
JABq1zYAEe/w7z+vLPC5hvfpMI40JBepuQKyaw98LRV+Jobt+Jfyt47B1MMXbo8/
rAGKdm7/zbWSLSOVlOlcsbk6d59jSZxxyl+Sh6vS8jYCQz9HKycqNVARl7toROMX
8NvRxBPpyxYidp8LFKZ9uk1D6A272VFLv9cGK/olAAjEk8C1cA3GJHHmvGSz0nfk
MeiZfQr66fPAE+scTEyE1iFI6lxGA+oKVpicX8hTmTfQ0OZOIaJjhsGkTWFHjfYu
q3wP4IAo1PAH1ixJoavxFUz373mlkLs4f4jLlSXAXsan1VaTbdMSzg9NKmHctsBx
jzyBQL3xPntFtjAv38ue1Lx3aGA5cpPHR04jTxhjHpmc+fnDu0eVdyeUw1IQfT1B
f7EoiesUydHAQStyfwM5NS6P6Wmc7lRiillgEMmfjOmtbeR/tVgXFctTP/z8qEKG
5OPVbfDm6fF+2QGs7Ie2eGrnQPjhsqMhvhek4SaE2ElrLO9gyptoCXIAAsdbZ+1O
t0Y34AhvJ9mEdf6uPqs+L9om3gWEtg44np+ESKef1EA5itjqI/LVEUBhVAbZ6Q0U
exDks4CO0mL740yg8wup01wxSfYMD+Cg2tlkr8Usiqh2k/ZPJW5OAT+CjRw/0TUY
eupTvEvX4gLfgruCUOAhoIUXYJihVN5qtSCDKqZAtIdLo2Jmm4gngjmpCwWypjXE
XvBZxfDDfSI/18DzULwN8QqkxE4nd2CkN7y3w8bxC3XHNs7hbubYme/09ISQMv+c
Q/rLGpfiBqY+AC5rWpdmmoVf02NUTC6XUupoFJ3v9BbCWmcOSOV7qR287XORCtnf
2DgcJKw0TmJK1N4PxjYFzs/nLgVqCFVH3jd4c9sfOFPMA5WBbZOCf1v0syp1Q7Ys
tw02vkVfsUIEQp/mG5mpFBEhjy+JZGbxXja9mbFSzGWywSMRjxHbp6f8w3iKRQZB
ocEn5cQdqO2iiyJI0VLrvXP8Z3RMz6Nb+xBnH2Phzk8a57x3UuX6MLzCzGPW2NUP
MQK7Kd8Uc69nERGuNdzGQTbmxCfyntkx6eJYo+ffxQKCJ6v5bQR24P3fHHPm1v3n
FADp/OnpBZhz59yQJgbHJTknSAFHBtJ6o680iRYGk9t+QEKVXkT4FLTTIi/tY0eF
es37bReAxAW++SK82wf+K5W/6Qs7wdXKmbKcx76AsLan/4Tv+9brxstPpUAc8qJm
8FClcQrTuYh6lSDtt3gmCZBmn81b0YOBIRdCW2hgnoOcEPsiy+xBLOEk5gTmVBM2
cBNk7+uTO5l1yy/MfJJ+I4mD2x+7Ke4/91Kry/oM9zdn7zQUMSXOVkUM2S+srjjO
r/0N8IaGxGuCLvBmTwgF7YHXs3PLBt6G/FyyMB4jSsgAETDyJMnESEbKHpepCpX7
7xlNp201yTdyUh/OiD3nK0hY2Pj5GkQrU83C/ahhq5rSkQf4TFi1jzW7ITYG/wLB
jziwKRx0jDWVKpXfMmcCC1QzynqdmVvmJ2nYp7JMAH1uT6SEIg0IzdKBDlhSY+yK
rdP31BFBwj/S9D5by9VBIObFTiTAWQSpfdlbyJz8RrWaiU7mipA2LdQ471mDz5MN
uLhr/5Xij+aeifB5Q0MGqtJOmwKC6Uzab8cTtHv4Ue642cKMbffjYeaLRN0b804U
QAvMBKPRCKwqqWQNSQW9S4agBEHKSeMZyit/+4YgqrpQZ80n8//rRwiVkCav7htF
zi0Xayt3PqZgkiqB/w42qH1oeOwj8ZTRYP1pTtXUWJkwicsWewsvhpgPIcnfH1D4
q9xl2tlpzAGD+yltn9mTVGYsha6UieI4YTyDtsimYTwmTz4Nt30YbUlb2kUMiUOp
I80WnVh4qIpJRS9iBCfpMx8UmZ14xfyJD3DMQOtakpG6Z/9iBgOdRXPNPdWBiANZ
5UCPTqT8dsyo6+48br/+/0AURpX0wuJd/J+WNrjpQIT9a0OLr4wJtAhznUiO7psT
6eMSUNinWSPLxrtfCUgqkNEcHLJc0xQZaO7FnayCeDTHuRXjQlkZcrCuezuV0+CB
16bRfj8ac30ZGmslU5HGmasNtU0SwK2qPdgOwCrIk/5URboBclwEWevyDV6K6SKM
2iFbc55l7P3BFvJ6P/TwBY3wrbC/UGFCX11bJ/790ucQml75FbeUdGuZyEqoRfcl
4QanxJRQetZB+8KnFBCvqP0zy6A92YuvZIBc9CTlc2dwaGTwJhJnR+5w6lhHM/vq
BxZ9EpTx31YugFGRt60Qau4EkoQfBn3ryRC+zBAQN+JjHrYPP6hRAMXU+ayBQ7mq
1ee4xWPGE6C4isabB6gczimthymjHhaWHGS4YqmHCOFTNTcjSDDOLTEz6mpCrM6b
4kfBlFOImwOZ1CUZQ1t/+tzc+wrE3XWoF1NT64RlXnYNrQmDBK1sFkH2b/Ierhpn
YqPSZj5VRH3OlSKi3Ke1+xVRcDFMrE+T1skCUjEXxIVa/2W5IUnBGmF5w0J8JW/C
pJv9QtRhqDaS5jwDyOajaU3f1Dw9rJFH4svDJImMR2qvkOuT8sRYi71psI3r50ol
gnQcOrcMkkU470+KyBcsmn1OUGsPyF2CtCwELZrq5bJizV+y4ehgirZzBC7h/EaI
HX4kYdoUvhHCPbadCY2BmfKt9vXY0wR6TcLt9S454DyoIdtZPiJGW/eAwqkTQuEP
lMn1p99sG9gkCjBCAB4j3VB82a6eNxeeBc07t69MWBd2Q1DLonhX7X78+j5mS1T9
RJw+ec0tCClhYQYfBf/GcUuYNxvLPspkFpfv0WWd4HdYnjQVVDMpDKFqAxBfpnWA
rbRYWVk6AgBR+GwNbGtV1tEh5HEU7RQkHitj0I9qZ1AZyquWEUCSvNsDqPCPyPbG
P8FvY9Y6xx+qTE5LxZdTD/HYP3lXoGqtuggWn0tcjldmhXl3uHEZx1hMthTjhmhT
YbABUo0uwoFohVZdanPhDHcCvAOlnWBWbo4HIctNAxt6f94d1UYzker29PhsePh8
ITZmkm3mAnCY9GjA4iPspU7bdFadfcw2qAMmkgSNwWtEw5ssrpaLwMqa/31yfgJO
yfkZvTMk25MUhuAhm2kN7CmVklE2me06UZ10iS6kd9IELFYLHz4/OSILFfkZKudb
+mpTMhp/r4zKjsttkBK0OWfPap1+ymBdB8FwHB4VPWpPD5JcAtTVkfGH5k48KnaE
Gm6n8VKtUNYnrWUeFgrFdeCJIEbA66IqYv0bL0ydQrCi7k65H+4sT9V7v4iVqj1N
HpMG1gVv4n1PDz9DK0YJkHoGoZ+QdZ0Kk7t4M3FMph8LPBHrrZcast6A1JEZsfwJ
TjUbuzfJrmSGLVdgIL/IAWIxbG4tapLP19+NEfEZPPWixbi9VjXa2z30Txr+AuPQ
FhX0Npm8V1iFs1dD46bil8PaYqqfEFq9nN9v+5u9whIMpPJf/pPety7/JQIX4igi
FLrv+in45k05LwC2iwjz8SY7ZN6nqG9kxqj9peOrwUl7D41hZbdbQa1wlzVSPPdN
qO30+nt0I54s/VeEfVJqNehccMF7S5I0++mtcgyp8mFsWh6kKJE7FaKD6xcaNWgY
jFPf6tFyvIbXd7KK/+Urtyn/ysDb0l/Nd0nbToKLvIw7dLgBgQjbGto8/maBbri5
`protect end_protected