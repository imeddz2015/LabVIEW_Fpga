`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 21408 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/9huKRhRMtvnNqb3Z+UU7TahEoHV+T8U3P3ufru7l1O
3DlgtZzb9QxCbOjthp9+wDkjygH0eUfDrEl1ovhZG61jZkkzENayPRivduqiGlqQ
3JusN4/7mY/80xGlabj81a0/CSDcKvTtGsl9TjozIRRINCVZeZQx6+5JlkCyvgh2
DjEhDqjPJj3DWgDrht//S9zfv1PLW9A6xo1+/8ZAoak3URRTXpp4azL64avbm/lb
jw7blY1WUhjxa2dQ3alJZFvXZXDfyRaC3fumeaM8Nh3bSORtd6Pmw1PTAZosy36X
TY+rOahuQ5mLDIByuPFlzkkZFEOJZQy4fgiTFwe4JI23TIZEWqQjQxkU8Qd02K85
5qyV1+xiOg7EgQS1rm+wVuwU1KTz16F51sVypuEPzfUBvwbCordbMUYD5qZtMJjG
jIXCEpEUfvwKE3p1LinPE9Q/dHf88s9G0Fadj0hKaDwz+ooI8Jz8JslgLn/ZO2OQ
atFJbHg7LnyZWnbsre0pnb3nUaAmtN5sQMVTfqPlxYgfxQHF5t9MeNjt3UM1W+mN
H03SpYQ08nTi0i/Wqny5/4fTGXZKkekVBXsD0Oh+Gk6BmwRWfCw2AkKuAzdmZOm0
51viHLqBLJ7t8sOHddhXmWv8f3mLWS9XZNa47uUkcazZeSamhcSnRrhKdFRWiA5D
F2bFK7rMLo8FT2jcV1/Ffq/aCUEjcXGlstj2aB8EtOrB7IVQg9aiAy3k734ggAnA
oE5BtyUCevgKiy0WSh1gcdbxIg+gq7c2srFz/VI3LJESCM7OAfjmckdCFNl4J9T2
1F1xio/ybpa60H15IV/R75617Rw3cQ7+LtFk3pKSRCAxO8AvC9j+lMrPiJI/V2iU
NttQ0sVIJV2TNS6yvc89KicxRG3pY1xdvD3csDcG2ql7W0+AlIul+5u04Mo3o8wM
s0jZDu6Nbyip/DLcZ3h/RHoD7MmJ0oyUEEevTXqvbmnMJXX5ktQTtHQjQi5KtrLw
tjL7qG5srNO3gJBoJHr/hHJGb6F1MjAH+cZdrF8Hcm4dum1Yc5AjqgKYDZBo+M63
/ymlBb+XhHgozMYDtxhGKQywnyoddJKciY0K67SquqULgWQjj0tiT2+WHVT/IK1S
pBABCFbwjvL6BlUfyP6eX8kTcUZjwstFbfaSz3sdgz20Il87TImR4tb3Gd53uNG7
HsoiGU1EmDUl9t4rn9ryszeeT2YoTSQDMX/CR6v98qtxxt8pRV356uX7nRCu4BH0
FkSXIpv3eJMgvAT2mcWUeeyrfUE0PxEW5WsJItcwMDIqwGPOleBgHKOxPKCdrC1X
XxQjY0saSB/zH0PAXu4Rwju0vIbiCKFYNYJIuhMNjAFXaNP4DsXgmyg3vXs0sKFX
pyd+brYggBmgEY03YorfQpWT5E9Rk+zmqrdRBRTqR1xWX1OaikkExLkXn8FFSPdd
iHJoNi29H4tMzozoM5xfECGru/UWQl8cbNdrNkD8XDjyrIbWT/DiNxw0zw0xSCGe
CiPz+/bt+O5R360nK0u8yGPEhFVy5TNIf4rvsamQ8l7Kqxpov91BWdKNCM+/pHJG
biAweeLRZwQ7Yx8GUJECQSJMEcXrfV4aQppmuRUr6QznNwT7v2YmGP/d1NTp5n8d
IYuZFxpp6VFw+3gltzA5krx2VkplE1ajvJqEHI7ygUjLjg4s6raPEjNN2KjkPgUD
KkCGvxPWvlJ62FeKJWC341SRZvkST/qsmN4aE9ZFt5R6uRv+r9J0Rn1RC3EYz8H5
Dv85Bqk4AmCvGl4tydWP2VbT/fYx+6Ph7j/OZWZ0gQZ9BuouctP/Ea3jdAXtr33i
dnwis7ciZ4Vi3tNJ8S1mXRxyg//ktD7/o3qDY2Ql14oTItrtQajaNhEa850CRW5M
NCP14BNvB0/z6q2YARsYUO4ExvDwEM9OtMTbWVvqE1h1g0krOtl9NGn+wF8Q1lK5
XC4rkYUp57ZHIrp4NbdDfPB5f3FDDeLg4WEuD8j8/5R6m4i5+AIvTMqKHlBAL0sM
cenh/CeQmGC/VR06B3ZirkELwMuqrOzbgjfrBpGpIvsgyxmYIdvf8YmidOVrl+89
awxxmdHJHEFLUtsZBIEjnGKWjHBPyMsjjMS1xl8d+IsRy7JRyQY4QMvq9tf8Wgzu
a4/XY7L2whEVtQt3XWQhrHu2rHQlbsoUT19HkdSBmOlDI/byrJBYCXwAStmZ64ww
xwJtUBu0LXPhqk/LNfd/cir25+yCWsWKFXOvmJThrztyhzZI1ckFGVGmEWI6noGO
REmExuweUH9inamdnicJOn/WzEjrSgFEQzc50cm0Gon7Ewr1zAhM6Sn8C6RazZzY
n39M7ZqQFx/6lekPntttjMDs/aYFBo+RlgBpl1iup3JWeKXLjGYLD6+iyg61ci5P
/yTKbO9riElL9mmzyDgfCTIjbombG+hzDFLtCCkD0acf/DvoNICMwDDsQA/HYFKq
wk8XICBImd9/qs02BlqaYTc112DDW0AX8e5FxJJRvm1ZRCvSMFcFN3qnq22U5lWz
DPbY6mHgRQbuNodcTkKAJaFfjo3IZYqEIcL/NavCT8jUuulF7mbtIS1tRZeitkwD
PrwK+uAexAXj4nphytBO3IUZOQbElEBDPrl+oWWWRrlTzXKLFY8JjetxejcwE9s/
mftU8egaolHfoWsKA5yTpV64nFyNce7gjGhWez53k1AzcQCOk+/tTA62nY0Dh5p5
RR1K/DbYZZWQFWLfykds35YsJhergwDDTyLSC1xmP24Lp5hb6X907NNl2gyl6Y+v
/ihdnGd8JCtxjcPRb+eyHjaWOixM8CL8jcLXZXjSFtT2/HDEXzDx5xqXlynjZUJ3
o6D39aIXaC5abkUdeiMrDNKcvcgPAMMHz/sIP0XxxIkS7A7fn3Cm6651SqvOkZpj
J5sqn25IJLkuACf/uwaKYOPITtURnSvio4MziNKGu6SEZLVH3GNQ6GlDh2unJZ8h
oFOT98h6jR7ugBbKn1pbeqf7QccYp4OyBO0sBM04Az670p0dXwAMCLHTywpJ/KPy
32NW4NOIUtClYi57yNg5HarKLjnkF3mJDER5TIL0Op/P/oVjPjv1zJ1S2dXgPwrA
D0PMsRKjFhe12lVZiEr8euzrYWzLpBO2URjPTBFyw/LsHu3/rPXhkTFLjb/D08oC
Cc3jlY6wYm8hS2cMEdJnV8PnLDwQaT4IjyJpN64+WBL3lE5WQQ06vgoRJMKgzyk/
+hwcrKREjDYgwhjRnvcSF/y1ZMqdHI5GDL5xJ7tjUjWRteWIXK5ydU3kIhwaiL5p
jp1kYp08VHRMG39pAoxmNAjv8BXGdlSE7caI/+884Q+ScBSD79Va6VRO/YsuoVx2
GcGDZVS+CipYo20qzVH7B0aFVZOQCjXQmSelgtgHZG2eOdycdDiztAK7VwrzubOs
nAiaJjiMAVmNiWirNmzKl00RjfuNAWwjgj9/ACmf953sIijJuZXqQ5iBXQ2A4iSj
U5TZN9gD62RCF28Xu9LrjDDnknAEufNOf0z5s2Avk3ZuBUEkoMeMxX/krkgp/JON
vHyD8wECEwDGDpoAziqBgIKzzBqZb3OvMARGgMeovosbxQ6LDvueQ7X2METq+1qZ
BFKqKr0nJ51AoJwT2IerDeQrSQcCA8auuePHtYcVkzpPpDG3VVIjOlXGAg6Iwx5w
7E8/27AwncgB3oSkmG7tmGbk2fEVH0jVg1fz7w5VXCygaIg2E2x4qH8uSUZGMDgn
Yr7h61RS/Xh3Zp8LTYRo8up22b0mCrnC4u3Pq1kcX77rx1bndl6j7kV8WOikKkQb
YaYtxtwk6PrlrSQ+XvzwGoqbkJQiWFBw92RWEu5eHhsmHiqX4085hyRgobUSQ3/l
TpmhiN5nJeXecCKVIi9ixqZclzejrjo2rijC0auR4BnDS3KsS/nQVSQwdj1bWl9j
5iaVdvniLvjgsOqX4C2p0v4mAl2oBRD9fnUR+i4y4u6q2JrcANqJqu03yl8zTw7F
5yLJcprWaj1rB18McofsLGUepDwvgRt0dShInGYMaKu/SZ2tceKXBuQvjR8hqQGH
3qzCxY4OymMcnSY3Y/KvorG42VMypXpsJBGyGB4XLtlJfjv7QILznm95rfvotGlm
xUbT2h7w1IrbgI5BTsipymkm1DazbUzZ7fsPwQNngTpiQxMSCtUCl4F6UV1f8fQ/
zwVhdWGWJC1rGedp3fmNtYnKp1hDvcA1Mz8U7nm2iK0d7jrrzczx1Wk7hkfFFTje
OVdlsjQgDhexkuOHzp9Nm+3KHHaSsy5offpnRja2vZyUKu/nNEoapAMK2HmiVZHH
PWjNmKV76vu3xvpaMCG0M4SCQ4phWgFY+Y3dZNKzrjq2tmYCQF96foPox+4LinSL
3p2fNwrHmlV7NvKZmxPzT6oFjnjDskoTPiNaWijiYV6qu0yatdgoyEoCszll8tfp
uaa3jb2f2SxqiQ8KlBSLhc/y389VXl3VweJ/GQ78VYywjeZ5nOg6AxN54nTfcc6M
jppYOFlHuzJ7/oyioxRbX1/CFRomdPrJ65oBjsCb8SzGOh1zHpWi0IO5KHgUbnXH
bHFWwyELWED9WyTnGKlqC0pstolC7I5LLNLJZ6WyvxPvdYJtZQX+YVjWLxFHTtE+
4CXIbCoDCat8gnV2eEWJOzgQ8pSsSX+Fc0AQ8mDIp1yNIdZr/Qg+kJ3eE8cdT1Xz
SxqnY4BCm48Az+hQW/6XeIKZMiO4gYYBaMHA1XmhmmOPE2opGPGdM53qKo6x6Gp9
Hc2tg/4SIEwpv3+mepRmvIodiy/k4sRQXDMul8guFjsxrJMFRHk/79t8Go2lbI/J
y7U1cbvtBDfwCbVhwrHm8lTZ80rbb9qJtwvR+IZRiwkXHNgpRHN0HM2sU1QKDLF2
9DTNNWdUOJ6MQoaeGjDpYf5g+LEc5zNslpy0o0lj/i0Fcb8yQn6Hi8A5uplE2bT3
zWQcDtd/kXjoYm4sTJ4WSixqjQp/ZNM9ibN6xrUfnCBQ0WQ9cb/2lkWAqaW57tL7
zlpRofoFaOfbMA7AwdB+TDZpggNO6REsVQgTXnslX7POBWLDN5yhZ8n+BPHvxPIL
yJW3CvDxfihXKtQn+D8zmTRuYB85z63cqsxLM9wzGX2xm+kz9rNrOLwy7IAV5VrJ
yMDClAY6vFON5mQ8/pjXHLp9sDWHcqxLzRDtnsvS9LGA0RevH67+oOGQ6+6RSrUy
9R5aT+Rf8X766CKorNVj/P+IeM4JFGDEnrwH9zdsd25ug0bAObO6BQZeZK2SwXW8
co9lE0Grpdp4VmfaurqMdJU/nm2caIBBt3aRW0ZcmBegDgAHiiPsjT2puSc4K8y8
poVVeyh5EpAanPnbwhHfNKp81jmmILH4bWoSCldQVoF4s+sB4GnTpIeha2B8TbSr
i2q3j9a9GjT4SuFDlMava/q+WBIO/Q4+Ddpg0VPzwqrUfcAQ2rLGJnuH7uigWwKY
xTCxF9zYBUilxtHnTQmNlIX9rLmSOWMlMT9trrbbZJM+yzaiKhWVD6x1UWUfBwrV
NX4rkay+wa8xjqdp615/NfACejfF0xwXqyj6xpjkHcCpAPRvvxrnATVSJFW0jakr
Q7hYTseSopMkHIWjJjsDxDLIc4bv/W+p/0CihXYeV56E5QfOSf63GeNrWjx08cEF
q5gMfih2WEHF/TckTtNB66kSbDM1VUUkR210eZqLxwVXbqLEa8FT9uvmuF43mv4Y
1da4CKrOvh3HnNfDpQa/9lgtFo5izVaoN2KsnPuw68XvyI0SYVrp/l0hyL7IFGeG
/w8KbjWPoDeiejfnmFYJvNDfbYcYXfpspsYChjlF30+fOT8OQWjrV+hXe3VqXYVE
4EmL7DAOtKiBkYJCbkPf1fJL2FbELnIPJ+ecDyGchbOTohHSkKD0k7ThZtAEL1rV
BOG3WWoBQv69zM4amBe6NrD0OqMGUhcjby3pNO81Mr0jd+mn8UTd6DK1ZUNNUCsx
3Q4mjDM1MZavaVeyYFijh7ljPElWIAJH5szD6/ZKYt4ZxwqgfJ2zaZLBv2Bqwle4
Zd/yFSiOIedHjX/cOE5JHpAxX/B1ShTZsLdcS/LULPZoaFBiGiYAg6ShP3Aml3n0
uVUXEgyBbmlT9dBYRuKfpJWa3Ekmz7Mljsy+BMv5odchT8p2oxeBzrlSnbbmbeH6
4Oq9KI/LBMomm/nEosj1AekGgpttOuz2HACOp9K9aVPkZ4M0NZ/bkVvsm4kwH9/c
MyWU6BdAuwx2I6HOwQAWbn1iHjVxI2iF32quFIuGutV8RFyRH3pkxwoDaEt5eNuv
SDhnQNV1bP5syBr1gdykfPCh2y88zoWI2bGtnjgs/XuzLcvKaCxPNp91UiHUREX/
yeHNhM1hLc2cPHOZcT79L3ptZGLMpQn3Cr+RyN99WCGuxul0Gyf1GT+1U/P6AJoT
cE0OIC5dkcgSwCnKODWR9txtpCfY/rv2YT0J28P4DM+0RK4zDlEWOK6HFSSrt+7G
xK60RvuxsKF08jXGrT2gqXR91MWdbictVYKbrENICUyDAoXBakVZE1wLRvlV4eSI
jDhFab1aMc2XeBSm9jFRrSfASoM4A1MioAm5cuM7jx87cL58MYpY/EzspyjVaNmQ
a+pYwEx/HgSSIiErsOonp2jI0gCPATMrXWJS+jHNdns3uF5bsLmq+G49Ma8upOss
y+ANtK8LJTpFoxiV0vGwDTdcdbTZNZ+BXj4lz+p8++3vq436EMkTSidfEwIH4728
jdM+RMfenaL9kkQXesIgFaMfMW+JPEUjcnsZD/NbB1xNoAjs9/txosErXyJjDkcd
qcZimvDY6sy6YlROffwVN+SErJGgG5cLaFsDg5FOGWTDpDw5gIbNBsQjADRHxgpX
F4jLDHKCB9ocQZCN+XFLGNz/T3XFe3F5Wknoe1AxG4D6oS6DfLmK7G/XpZwZdvw2
Lxp5MHIG8Miirzqr4fjOKsdc+AowLKV636W5NqW2sUy161cd/srLvP+g7bchKZAi
pFKU2y1YjKURUQEdD0+FAeKWi7oNmY8tT/+KnJPJehH93n4742rixbuJjp+dbK1c
UMd3Ct9CkwcihX9h+npm3lnx7ry9S7N1gRlisoq0tg6NvKx5tsDfGQ0l7KA2w4CK
A1D5r6want44+jfqe7tCjgL/VXqXiTLzpVUyfVjFMqI+Iw3emnK5Au+06CYYOOhJ
lVvfGB5bNBdPqPxVDaTI1dUwrOnCHyNNSLG1Oxkr8p3KemG5w27Lf94EhtwP/uRq
SzylPimCHPH67lb+bDuJRlzMdNN/ag4wZumQalGAgO/9WjeL+DdNeOJf8mM/UGJR
4R3rIawtui4RVpSTeZ1zMB7NXNJGOmkiOL9ocYUseoYPcx0UNkO3wIH6Dwv+4PYV
TQf4241dWqVf768OL3wyFREHKPABxDFA7BKzh/g5Zcm309yfCLJBtkdJaDrwOi/e
xY15Egx/tTc78KYTSzLX+wuzidzjJuLz2sjJMfy+VEYlwPi+5gmwJ84Tv/gbcvYx
Q6VtoCVmPcOhM+4V2dGCBdf1cSv0pgSNoAfVNKkWxTOE1MDWYBnBTCWJM2d044Jz
bTw/xt/dlQivc3Gc37ARiha4pvhzJJzLsl3xP4YQIDAug4nsL97YTms85ZS5UUds
QVXRSDIdFTTox0yHmOBqs3KFA+7ehgHbRIDPQYAT4a21MFMTGz6h+z7GyNLlPBfU
NlvLPLJTP9uScxgzl9IKikxpn0a8iJd06tOzNZeRP2DtaItFAGWKENKm8f8vvmPS
WzqehUCG9au1G/ZICzn0A1gzjmFiOkKeFEfaO0J3IIwYaG4R8LzV7b4HVBd2ny+B
LdDzaUbnJpc9O1MkvnM7yK6zaTp3rYpEgrrTq5EQbm9Ubf43UGZ7KMv8kjNsdY8v
AjfZuA4B3BckoNLFLfsLB7ZtMY89X/z8HztpU0I7v05Im3YSQugNWD8wvDIekJQH
rHD3Guwu9QBxZANBm79P+ByNkvItoBi7q2kcQR/GzQAmBLCpbEsErck5Gg1G8NB9
QIjkJEi6MFLA88gX/qxd/9e59Gqdq6Giu6Kx2mjfzkp/jL8nSfsSjuuNjOJE6Zx7
Wjx6q9mt2KzIfZDC2z/7CP68ea9vMhyAG2wnSUEXxdF2g5UuBRNRI5iTB08yWkb8
B+iGqUMmlAfmxWksHUF7c2w4LjuYG/4spgDU/tbVOLPx+x0KrB/bGoxFiFk5E3Mn
OgSREH5/awxPuANRAjHYE1PwdMc4JWvVtbRYSEX9tmSLPQZpj5bS9LdsS/YUS4wV
hsk5GKR8rVZ8KLzWpo1gtHJkR24xlBc7g6G+3JLfAICeJIJqEUNWyWgEz2EYFNhM
qJ/ZnTAYCVvUMXgPig5n2FT/df9kO8Iim84LxymawxlDBciQQ1IP/UQrzdwx3TtH
iwfVxyDhRwSuiBofpD1YxjrnV8BapW36v+ItYp4mI64NxqS9wejyFtpbt/uwYMY9
LTKwUkg3uCPAdbCAaHB6McZisTA/CP4NyXhlNo5BcI4ONh2PPB0ly/hjrMAuKpKC
AXUipsbRLXaZuJ90xkqqNr9rtwWT2P7LVXnh1MAvoBQREgDXtWrZAyEAD0ECl9G/
b7p+8fNZnbXMTfBZ/Yxr6ix4LmkCkQT/TqwTYz3W0z1hUWW7cSyarRkFifJNPXAV
0S7ZMCXppnSMDfsDntBpcWL3NBUUpuEN9V5q7PPRY99MaCafbIfdy0eVcwDJ7G+m
t3L+MxO5UplU+qPL94vYFwnCqUByU9S8OEJGmHZUPBFZ8Dw5SXGl3i91NVYTVU7w
AjdYVaohtFZG/MFq7CZg7ZW0ZxQcdwEK40Uabgw67YN6gvv+M6Aoh7q3Wr2S4Vth
FJSnCuadPROErfH9mGtgvW1iE8aDTprzNfOBngOzrJaUxjQOabp2vRA1muO3G2os
vjH7GPfIfE/djbOEgV47UhVhkqLA6+n3lU+jXN28BfSCDNz4qahnvs4DTJKYexfQ
cqwke75cwotr/zm2quOh1btgfOPbQA4r9Zl/T3UAtTB0ZE5lEckYRLZN7sSYdPrU
R18Ng73kjSpbkx/Dc9tGLT9kl5mEHy3elcW3HEVT6vwiNXJEBorv29Tmf9yCnl0O
2bkgKeuBfgtv2LrXOoPk4OfNeD5JsJVAv6eTG32uZ5QabIqew+X/kiw4LdExH11P
VBsnbWkS7UYBFuu5+0rGQHN1HdWdEvuPsT9lrphizC3EPSMiaekrhuHjOg6lhf3R
ZSP0DCx3GjJyzSH9jGd2pNxwFCJqRvJVyTNAyg0Mj9g42MSofBx61A9hX76Q41WQ
BlJ25C+1RBbmtOKuqLTS9/01kHp1uX/dWqtwBs5O8386hcuLz4rhmgIbgObDHcI2
P3wMTgrB6kHMktKHsatYRCQNI46lqaL3ht3NrCnF05bsaLVuPbMqMG4n3jDSBGPa
oL5OXoBrqr+3vg3V7b+bgbT9sxvmNLyrL0PiP16UN3Uft978SY1mywRAZ7J436VZ
RVIMVpPGW35sRpqnXEu97T36N28BsHUeJU+a/FEWBCCTZapCMZnlKaSDMBOL9cPe
I3hRMgX9wRanbWV09xLA8cCe579E1dBRrsIt0ZkuvDp8NcMj6hV1PHonci11+Qkf
bnogqsrFusvq/T+m9KaD7hzE7Rasl15bOf9scSz95wru1IZpDYPpblE0NcREl31G
1L2+TLiRqcMdbt9RJ+/KtR+aF82pyM1VvfrsanTWrJNpgSnNlx3U353edAiKPU0F
HVi2uFFdTcbRhDv1M8SrzgEiXLwTUfw5O/Tmw8+AIX4y+fHGZ7dwmjDpLoJpE56K
O2qoUTUuVVdSDz/GJ65yEZk0AdUUMinqFsCidBL3Ul90cM89HFsbywq19c7RZTFd
ic0DHnnh4DbhZWSF7nHv2J18fLteCm/UTHSUZAcCYy7EMOVMbyEuneW928cNrGGY
zjBAPm5PREmsmx3lSQBt54Hy70CsGWfbDE3AFIo6EfCiGmHrSFK3st23y9XNYOf8
r8KxCzZMzcF7h/PtZqYOsW8/8k/k6SXrjK9FzxozW82tRf9H4/b8MU3bLn3qC3U7
kig8WFQnoiG78ylKqJGj/2JUmtl38t+7t3995QVHRfbMO6QUV+emIIJ0TQHvbeiL
FjGzXBqCTRoqiZ4CG8SmWg+Ytck4Qurrp2bx39jorMtYSajVBCR053GELmg+oIRk
UOssQfKGPeC/x8iKNra1z97IOuOJv2BUD0Tq1DNtwKvevzFkFGPaksg5gk9xCN7N
2VyX/i2Gb3xwIZiSTIyt8gfIPAQScqb89RsL5hT/8DNDKXZ0sgdxuuoOAeKCh/Ws
JPRqDH/+QQS+UHgi/lM+vBtDCv7NN14m9P1swZ9lgkGzWL5GR4gDTdVv0PXbelEU
qc7iXi1sOjk78k+gaf2MQOKZuDk4JFT6Uc4hXAI0Am6EFhgpJaok+zmOcNgS4aNq
m2SnFucwCRvvv0vmotZb3kuVHi+vxbzvnFF7pjGrkcvTtcOsmjdgmlJ1v5PXf2Kx
xKaDXyhxN/GFUHiLG6HbwUBzEbo8DyHT7elVsFxaZdYHSshzhBw12NeSZcRlPi/j
4lu/QFnaqWgB4ZfPB/TLE0p92ou1LyrcY4ndGxoRhO7r+EielFt7uP4aeJLNjenv
SOmrOUQUWfpdM3q1haRLJmZnirmK1g3dSGVFpDcty7EtEdBz1QYGBv8Lk08esy5G
16oxzhg6JnwAGrXOfnZBtMdFOhgpqrfMUiVPkGvk0IW8v3mva6wMRmtHu8eKGzvt
azmX3ACsJaTPb6Gr+VFtl+Il949QYoVJyWWju2TuQT4DN2/1exFbJcyidkS+iLD0
/Z7FuNRVZ9L1jCTjrY0YZkrlkjwW2pfOMq7DmSd3bUJHe3hNpgATuT456+/aumYb
he7Z+9gs0t2UzysXL+q3GfvGfaXvMpeRe1nUXq0y/TsjjUzNDCFYOWYWjI34NIFY
Q+4LE/6ANtcnjb1gCRoWn55NRtUwWFkHT5lMGxzJWkgY++s8npQPyS6f5OI9sjhD
MbxfGEFHzI5Kl975RXa68qvJp59SYIsnQLhSCTKodsFeHxhNKDcdkdXmi+du6mtj
5mRVshAFlW7q5BDDcLVyuRBNElCzBw+X6LviVckWv3y5lNSXWFJFv9RbkTfq0S2X
i44PcfP8+l53rgKYSTotXoUKMltAW8KV1z6EW+gF7waZjPl8g86mTo7stug0flLg
5aQujCY3adkVseyVNmfY8XKt6BRNe6LR1gHj7ReEUPcMrdmMa8a3xOoQSAnxEVo4
kwBZ8VCZdftP5UI3LLof3LsRFXWZwfuqfdZtaZNg1z6vNrQCWj21uLE3ds3H2kz3
EN/DdAyEgOFoZ3Luq7RktdkGnYOQOEuE97VflccmsBjRlTULKADip/0mXgfaDROs
JJ5noo8JrlFaQyvrrBdbXYXNrp+7xhpleb41SAKEZpsKLu+FYd1Mvsz+GrlsKH1l
IEsX69qGCIbixW3fQ5p1LfXVgd7yp6zpBD6HoaBYjC+RkEDICyAvYsdOIWfVBZ/9
2ECKju99ONHoJoM72/7aduek2Hq4L26pKs93ZVfPYLrTBh466MYrBQ47gggvcxW3
xYh5aPjw8KL6pdw7jB4iFyhQYH8wRSWaMvVFTVwlE8pnfPC8yC14VwxF1oRg3fRv
Tt9bOSDB5nyiwjf2a7n4KmdmoJlnkYUzpVFU9/2PIQgS4k/ePfZKd7cF/1hFs5Hj
lWBNw1SJpPPLxolzlBZJruHN0d9S1n5xwee0o+fTmWtZDYzN6KpT2kS0B9kwW1iw
z7p8oT5Cxz6TkbtAvXxWRsdD8/4medKX1Uq0ZuLx88rHPvsK7IPExUj614YoCJIn
xMC9aBmMEQ/+E69vpluVN+qCsfqap1/pDOqNd7p5PGunU/f0oBQqFJ9YxgWQO+ek
Gdoz2CV138LucBHe8qCD00sDvAkIiIniKC3Ls2sK8n79slQGKNvUQ7Y6udMaAtCq
Sz8Y7GbJc1ZUP08VPGVBOuopppUVYXuGIdtySez1cfzmYL7zPHlaBexHZ2cyyDDv
DBOKGh/G4X4Qq/AoxeNRTJADJ3+PLDH+WAfYxfqre1Jx4BHjlefaN4G/k1cXFVh0
51F3rYWaik5yqDGWgaeiAMhcpTOyLW7Eroznacnfml4N8tlCj+MwIGEsawmPOhN1
6YELCwCwK8PtmW1OnxIZAeJXiFJ9J1HgrDevXA0T5GFaJIvnZ2zPN4Fx3OPwQGII
CQpTFrzimW4OHWWSksMgz5GFBF61hgSfWRlRKVMkAeXuJnu3PxcLOGq5bBoaW7CD
cVEyw4rFnPulNAXZfCSNqAYR3/Xzsqga99JvhewPA1dolP8dupEtU9MCOrVZ0WV7
3/k3qsplfi2G5MH3jm5umdNBCnoRTNWifbezO6Z8gkWQasJ7xn3wntO3K6yauAUw
DVCsnfBtJJFHBvyR/5Ha1rKDFggbqaaSEnwg2+NP7pW9vRCt5UeYTBktwQzldKYZ
3kL0+rP7UQ9bJh2tSKbj+ANrSwUE27PkFSsT9jeW8eh8Y5cfX5q347IpZYssvonu
VAcX+IiinJQwtzDAgDSwHCbmftPbnoTjS2kjp+TsXHtJwmxffJWrmE+W/S8vT7o5
MeEtyh5g3K7aPuzDZpxwQFVEFhroUiNqJZbL00OjkklJvix24ehFYHzMkrZLnEk4
kHQ7mg6Y7/x9uxM2tK11T0tEyzk7rM52SEEmdEFCDycM+3xKQhDwNWIn4TLtpOpb
c5iviTi/uO5GrG9ywwB+cQa3+jZs6GeIrS6+v20DZDDRIjVV3fkb1rIohkNF6ONp
p6MZ9HNuP24Qh6fSFHCQWA+jiMp7E4wQKMlPMBgpH5v29+HttBCB4YgJWuwSXk+i
t55MUM0xFdzlCznGSkVc+SZB1rbaSdnb8aY9h9k8jO8OORWyuLPWGpcdjcPXCY/y
ZkI2wo7fqyWBYN/q/Qv0ouAZoBiia73p+8utCulwwd5pdgIRSVgD2Lz2/JI36Tac
/edOOi8KYjrZmJlfsg3KZuPWqMigAEDgwTQUb+1QnF36RA82lr8i7PiTxrjSgT/i
9MDZAH/UF0NPTVm1HNCHXVCr0zQOAdDOBAU7p6BfRFrioXNm+tKrBRnG4mWeJaC5
Zf3PvUokCsAxrrcdGGEpOLVa5yFKwQhz79aQJoH6e0btS0c7/qML3b+1mCmoo7qQ
Dz8VsMKO5Vd2+NfUGZ4JaTF+0d9FMVVY4e2JPn70TPUfezxMmjeizx8wyJZzeVEu
KQqVL5Jlumhbi0QCTbdp02ZWshvj38VbB8to2Qv7B9oR/ZXphRbCnsun9GfTap85
ypxaz+QE/8iDGDy6vtXJM+K7xwiJq4mfqkPpAqlub8Bh2MX4fRe4Pthh9N8CvWiQ
5Ah5Uxv85IMAPJkadw+FjnMcIivoSyZ0y6UYxUkncDRv9uy1uTLYTeeMbvKLYWLt
v1w3LDCXURvqL0CIX+VuNQy3tmwAAwLTyp41R9GwIOg73zQEzDRQHb0zuqzDaNmV
k7GB6JS0XDrTl8aMGvUfNcdirJUw6/WHEv0/QCH4zCfUIKf0hoVSfoL0IBWgDPRA
iS+CtMaGFzUgeLcus+rknSHRj3I2aeOpIR8/WKjQkBf6oaqzFwVUNjnlGG5awOjp
T9V8md3UpBNsPWtHoZWRWWogoP8drI0i/RJrkrvIpOE8dh9zdrC8ZbJx5JXLqKB6
qS91cIxHuyodohTV978GmfjjNkOGAMU27tWacun3LCPEETIvm/x5KN2vE5GMbExL
kiDsyoz59OuXayWmAW483wW6RRhwv++4VOUY9jzpHJ81RBlbJkdAh0ttl7af05uy
gjOW/KBZ6FVGjqYwswuE/Ha0eSsvELSK2tV51pNOi/dwl7y+G6W6JWBF2Cmwy/c+
M70abSYW3qSa7cVpZXwaJCFESI1J1+V1Uz5pBdzhXOia/Fk1qw37Vj8F6HloFuIq
qO7d9fJ0NYFolaS8dQKJm67TawnRrR6W13ciqgsuNyjSA96bzHPwD8YiOiSW/hO5
4O6WskiIqrfMg4Va3lVK5N7reGVDqRJQIP0M/ID7Y/UDq3QAHFvxPJufx3Y/9Czr
2qUxmFnjdjdNc3o5JHgk9B1A6z2x395ey3pBf3skuYdfinnj/t0Y2cYwHdBlGbhp
+NnutRvsenLew525lYEsC/F7hEyzeNn+vP1zlTEBPZjVf2Lfxh+T67g01QE0qjo9
wbSdCC0Adizis8uDeZwGb1MyfOLM2D6A4uBROKc2SooWhKqmsd8zWofgdEHN1gVW
A8UNZh1naPUDpVhaghsL7roZcbMbLcLSHK0mrFi8TYu4XurbD8FpVhrDSlr+ERLc
vg6qQzQG9v63PgIJvlvoxmZicqhq2eStV76FRZEelc0ZvwLzvyULpag+ssYNTpmK
OuwNLp+uI/YMiZ8PpLWpwqokwKmRNyqGlec5xzKXi7I+e54lpXfWQxmS85YuGVTi
euVRqKYBzo26JbRLyFJKsL/sAlafxCtp9JVockGnNysPQpTZNiAJeSJ2jHkjFdz/
XmnyGBapaLlkNqlNkwTJdihTuT5qRazSepTIJuvefWRort2VJgXZ+dArZKzwkM8W
dDkClGbayf305immmk2S+N3Z4YJlhbGgSc1R4vnwhdlyP4swlrKYieLqPkLUcEmW
DYFdZW/FBsueY/mAkqEAi6d9DenjLlnAmkMEOwO5fZVASpi74H/40mnwe1jYiWbs
j8S4A9+SiT6aeLtBgatq4d6wrneFp/tVwxwsYTE8wJPvozCtXJK0bdU+C3FkYrNi
tADouoQ1ZdvKEbY2XVBaiLmlEHT23Zz1lLLCqFiBhKhY4hNW/O6G+uA48tXM+bjI
82KrW/KGpGCgQbhge15ITFlfe/CYHta73mjt7SrCkMjNgepjLufz+ngUhW+EASqO
bF7Fk9Jkiuj4CfAmG3Yh0Wox2AvLW6Gm7lskmDq7D1DfbYaqkfP63/4BYBPae8Iw
oQB8gfSbs4ebb1m4PKeLaTEP/DOyR3TXyMPpv3UxAwqrkZ7WiT0TThX+WuHfEw2M
JWuWe/n1/l84WaknGtiyJ7TxWgITrX+mPlX8Uj3YbanIIPMyQMNKQ5ELkYV57wMu
dXkoCh+DHE+m1/k0hg+Dt2dnJBPCbph7h8cl3q3PRD5/YYuKwM0sXHNeFzvAcGq1
2PNsPsi9nunjnk6uYYL1xfNN6y+trzOtp1JvWbfADa3INvoMFBiGpvpIYTFkomWW
DtTvC+a932Ms7ZwkakS8gx36ivNeqOTyVLoL4pHrC9az+Xpv+bq1ico9E/n0CAnt
fbgOqyjhnywfe6+exlvoLHesvESGXInt6cjrdzZ91axwCY18n2suPpqR3BU5arJW
BLPJL809UvWtxZoxDb6gMkJX/GvPoiFGdwzpQYQAP+6sRb8Y8Va93hfgFD/SHich
ayNb1Qou4IB6LnpX9hXvOBRbfhxkasMKSKQuIbIRMohemMlxOezyf+UFni3K9JUe
7j9rNLh8S+1fCV8vGdXJkEctoz95B/vX4qKDcGR3Q6KD7l0gEIB9xg96K4ewlvQN
AOqYrlCQ6gAHGnq/1+cZamFomIQpCCv7vHviMX86BC98+nz8TzQA/yo6r0/GOSrp
aFW5lygsQG4Br9WTeBwpGjPBD8OLEOH2oGW2kG3qCxG5GuGQJGkPWBaL7uE7z1TF
KKIUqy0cIemw4dhHKnUR07CMWT1kaWXo3TzAWNl0l110NDFWPhELmrq+rtaVTM66
MUNYTfoW8KE3C7m9ipDW9O/7M6pnCs+BwgxOQ5bdHeMv+i3wkcV6hKZL3minH+CU
lgAmaENZ9pAQ+9mhVynKUjpqwxiPGpSzKvKD7JAY9X6+DKeWPkZZZOp1Vyb0NErl
Y4EpeMaL6aRKWKO0GSkierbYlt+edLt8fawbRPBFeBchyB3n1CSopt1lWh5KsBuc
f5aTVjyjy/DKprhoLZy1EGx14nKLCdqDcfGvgFAYp+rMeEi4VBneQC5gx24kXa9V
MKgaAne08yF2HC6VnRUfIdIqYEf4bjm+jxO7zRLkzFUVNKHkJgrOCfTDzIQaZHzX
N9jreKir8AdVFKd0JWHafWq0dYj4K+KBR6rs7RKB1WEi6394pLjukwHZNtrjTZII
AHL9ovTQcM6s4ApdvUYyPGxPa5jpkbmD/Reapv6MqWQniJe5r0n+3UxJxOzbs7F/
OS4/kZbv9063plPYzSRScSl82T/4wNGG6kA32msQlXBlXBiJRIA5T7h+ANZsb24u
IAmpS02HGoJFUmfKuyOY240xSKwwQbz/y3/yrIxOKkm77CN7PrVJ18CBFD+3ePKj
SXZMz9vpL4QJm2qbx8e28ug+uFwNASWiqTZZsMYWzG6iDFjsAwOvKKyrcTfFBgOT
HKrYWzvVbUOcRwHiia/1au4yN/7nvQGGjfr3/fMZlfntinspLq54JI0f/R10KWu/
xAXvjZ6oqmQ65NbV6qKg+kCmhx4QifNsRY2mAbynE6ykKnYx0oJEUT6yEXsUOIUE
FpwaGeLeRShbL00NfozKQdkrE7YyGNp+DivZ5zGmRLZLPZk8UaQV10bO6LJcvnRu
aVmpwhvKiOytASRrrWh3sZG4nf2oTFRFHGX8GgtiE+0qvuxAs/DHthk/iebq9bYn
jKJVnigeCadyuZG9jcTW+rDJY6y+JKNJaZAFVVDuRRhJVQCYpjrrs9pc6RPfcBEv
3rwB7M14HtHxkiYpeGe1F5p/EmjxHHK9wFnOZl0gGRzbzo8z1j3kSXbg3avegyhh
f7hUEOmzn+dgawKeQr1KGnUArTZ43EY1fpdF7G9NaQ6EfyD6ykMDxrBDXees2g4L
1NjM/TRxx0Dyn5KBNNkFYqBMpC4G9nysX9gBE1BkggCeZeGbm5H76h8G5aURdVl4
0HoHZTA84V8kh3ovCDV645Va7QS/2SplbknjFyOAHH4dLeKxGRDxzrNs3Ta9d+Bb
cedggMuzjFhVIKkPZDtX/AqwEpwn0GWdlaHJ223Hw4T/s0GPkcK5EjPkpdG7KOX2
S3x2JnNXXndA+hjUnELnv8ij8dl92N2bYxjCVGqm2UVe5pLRsVCLm1cRfFR3vuEZ
T05HL/fubomckSvmcVyhXtGlb91BtMEv9b+E6Q4rJGlhgrsFdNlZATXtb4zoEVLl
OiKdlSNjG/cank+7Yub4+vu8w2yMcrzFzy38ttrnxBD1QlQGzYqgoUzdSfPaeGKx
aH5S6lo5WRJGLFXzJLXG1rc0/dTTLdtDftnPWVcad8rq8oCv2poHNtK2xMb7TYoR
ASPIlt5UhWFv1gAifTHkLjBoQ0CORhyFskKS2qh0rfVhfBllJ30Ndksa2S+g+Fe6
0HYbXmBikB4OS/Ymnq3awj1VuxnPInq0pjbK/sRZ+1cVJjKk+e0Ng6mklEBy187Z
lPOyyepmvsoUFo7Rg7Qj+i7tYY61xZhW3D0vfdzejhsy/N1VDdugyX8U6BAgaV8t
kzQ2CEziNvCzBevN0vr0wc/H1HvDSUll4ELkDeoHfxrPCqE+miwwNw8meJXzqGJM
PvMA9nU3XsOl7+O9dGgKm1aYiAVr1HsuIX1U+f/s9e+tb85Mz7AtaFZP6HgaCJ4f
RdHGALT6r2dTWG7Y7r/P39pzxBNI5K09kLXdJK/vvdLfxK0bW1ARDyslqSAbkgiy
hh2DHWRlaq2suDZ+9G1wU8vHQ20z/9GNFPRFZo4+YqvOTJKnPzT4QirdhKROy8uK
uXEbiY6JL1mNdeFgeWlwmF+nfihiu2SjjU3EzY8QjJQpi6PZq1QobW5TDminEeJo
0bFk4ni0+WOtLBsdaz92fV9dKYNdtYtY0ytiLX0/OtMFeZjtCKQz1ggE5vSyFFNj
uA7LOwV6dGur7Xvft1f4ICKc919fX6jhJG9tYOoDlAx0jXdqKA2Tpfj2oA6vFqs3
UIHv9RkzHM3TQWG8LxUlFiATrBCpJXBSbA2kfzz0PxRwDh0kmru/Le3lHHsMXjym
9JztFwAj7fom1wOE4ufkYBQfLUiyq4d2A9VOYNafwabtVX9o++d1zFHcyEv5iNil
4caYxzn0zu+k8Wt+n/osjD1FlOnIJgd+a6KEk3YJ69923IYtkRHvdK55VvJF8iWn
xuPu0RZqp23lR6sfjbh8yNDzZ/8dOtnu8D4FbjSx0oot42dZLcaTqYhJJIEV80n5
Hx7oTwUno9sb7o2WAFjfmV93Lg2FEOr32IMtBI0TqkiiwsDe1W66eG48tr/IDb9q
GYBV1RnaD0iVWtjwokK9nrXNJyra62WQ2Vu2Iuqba+vLhVp+9OUziYEfpWKzcW/q
LS6d2q2TPJmw7fd6lxE1YCkttRu0yuvVmn+E4WTDwNnaFNMQLE0jCY8tMPgo3/Mz
HelebLRwomd5cIY+2fOnHz+0Nwclsxudi8gd/ziu4ZN7wPKAufdUUGi2+VCRgMrr
HJ3+lf2VMwBdbGaK8Ba04XWB/j0/Zu7EipW6FFgTM7Yd3CJDomugHsfQ3dOWQV+J
J+tf85LrDkNM1fuh/jZxtgCNBrg8uP2Rdsa4l/haVAE684t97UUO0JBVWYJUxHgL
XUwoxOYFx4lauy+SqnIH2DHK8CuW/7JgCCBcBl2IZgQ2jCKwLVUCjAyTWfvyDsrr
QHcz9gklO5ctcND5IG5HqX/dsaDrpeAXm5lZ8QD/Ki6APjqmwQCSB6JKM+qVeIxN
LwPax9xlpAw7NjlImqPYfHKiqhm/SVmw827kC95y7NlsUc6pj8p1ZDcddMOK/Y3p
E8qJxMkUNgVg2jL7yZnv4iWHNUcqyZKrnPlZMcRm/CP0lXRaf1V/hwyrCp5JS5LV
hPGxkMU4OlKSnG/ssWjp3AfjJcpFSA6mAWNzAftOpKzPbCwjoed+gYAayKu44vjC
ncCciGzi1ODxabhscgg29cfx/Ir8i4oiqJePKtyZXzv1wfmvjSKdj3BiptNHod5r
DPxrWwlicaRnRVNJ1+tQY1xbY4ewXj0ubWh9eVDEuuUZn40XpSqHlRlYmSB04QGJ
JJV7ygUt161IBpBqSExNzrMd04GcGBbZGP9lnsB4fnevMjsNnJsXd6bKYSZ/9M+C
UKjFJiSBcnzw/xnWPpyg+Fjg6rZmJdY+j+k7/I3nLyfz1O33QvRqtxKaC5mw9Twu
U+MPDhRTfk7MZ0RGm/nHN0Ic1cBmPVE2lkkClM8Te9KVPsrNs/5h3GffgL1NGdKG
i6Q0cv7Mw4micMHUe3XEIFGT+8RqgGvy593DBAbNhanVnKPKbwHBvXM1nhYbRX/K
fedOOJ5PcHpOmkRp2mrnz0iEhtTwFhfC9Zsctd/B6yqOU/814HQjCSREL+8H5q1E
jkXhoqfaHbReA3DOlRHYdI9DyUhvHNfdiriezlvAdWe0Y6KsOXffvTNOgbjLbeiS
TyYuPCxd6nKbSKOC1G9Y3nN/ZgOFW06BseHU8SKidqmcyemmf5QlriannyrgcVbV
z8NGrWkqVT1sa1ViK+PR4vAdFzVzxH41qlbI6+ug+vuYDf+VdkvwSwuyR444V7YV
9bDQ/kJqtob7JfD4cL+JytCqq3qB5Bt6d8SJDisG4PKNS3emJjLuJZICDbFIJ3+P
o/JGl2W0UVFrGxFYrVQ/ycvXacleODbQkt1DFl0eS3bVkc1VEmfdY2HXZtVk+WFR
GvNsVoH2dalHI6qjQTgOgc6wJGjMh81uYnuW9EUo6W5kLxdR6RvkXkP1oOoxDR/z
ezW0ALMx9LsfGHH5IDlToBDxZigcIEOBx3zQEPvXDvh+1k5B93UuCT1UVXZOmJDv
yg3rleDTZV4jXGLd6ABfDUZR3v6Uc94P0OOWxrat+US+/iOPG5e1nUT/K1r4F5La
549iuw1YCkB4KvaWlM2kT02WlKXOzuZqZhX7fjQ4kpsZ7fa/+f06diFkmxWT4dqA
NKcJHk8vOWP8FsJ2MU5QJrg6GLQkChTrVxcirTjEX5pa0DeU4IsHR9STLvvuvk10
sguqNqyMVymZFKlrKjotIxxKPmmN/VTYQBvGzeFIu6YIbN4eZssNqJ2So9iBxLKj
S3iywHnT8vqa/CBP6hGbBrMH2fVlmUIoVurooXiY7ErIcsknMeeYN3ml+76X5uXA
D7/alVcwiebtqzBjXJhpMpRAr22NzCm6ZqfKPToc5w6qsR4p9ffBH8XgdOcUq2zh
j7JGALkpmKYl1N7p+9lQzVrExMt4co7PSjM8cvDdnTRa2pZJv92lDxXifZNVdWdP
qk9OAoDUTsStVuCaOGybef7S1pXcnxmTBXIWnoIUS7iprr3yQlFRS1C7glm203ji
LsDIrNTnpwRAkgoDfasNtPKro2PdSEg+xRsB31xPmBKzqbbQQTugBrzAlxt6EEFx
A7WYOYyk6mUkKMT55/jr+K6suqcn926zI3GkHX1wdH7HRhyKsytAcImXhvDgsUn8
Dz5r7tMuKXtVeD3epCOUsuYsKKh8ZTknffAEVNI8RLDMkimgbQCmFnRZecYf9dCg
mNuru/h/Ik0Mh668Z3n5BFNuIYOAanespYZRW3i6YToSwsVg1kagvXCmcSy1GR3C
8yGkF+zb4itKB8MovHizIPMA8sJkJVUBEnVkVTxpQK/ZuDC8kA8KRUHtRWF7DTfE
t0ffnCIPo3cF/RLb3B+fhSvk8o+PbLHRxLgMawtKlLqQWvX3gxBnvCKUTkrTpE9Z
LzAWDiz1NNTEKq1BaTuqexraqB1xxzi51ZaXFscy28NZm6IPEtWhc5LtlCT/IXZc
iUPk52dwuVwpuLCqS/MQggLgWUwPWTFAgpO0XMOT+fVsJnIj3vz8Q7eIksqtTTjc
MBUo/pcs5pkR6vHUHxkZoroC65zfciowc6XAWCw+dc0D/4nkxT8vpPje3c+0OOir
bAdXk+CdXiZRZ6NrCuG/sKJZoQkZ0aBnVinRkkfj8bBrTlYA0nUMK5Jhabh/Df/R
RfMpNP+Gal4kgCS58Bgj2rQO1CeKya6pg+th93Uw7MBRl+ZY0uFdsgz9IjetMMDx
zhkK6BiZ6eKSsjLxxVgpFdj91KZ0kWl1FBli0UxyXJq76Rh6mRL//admPJtTvrIP
E1AB/Vnn6HSKtx4u3UtE+xDgTACO/lXxUtjkUv1Wqu6vFfHLRgz4uPexXzK99M86
inzquUc5ryRtCU7hEOvimy2yFVpuuhfgtFRbjVn4tkEFIqtYsS+oXMSLBuZ/4Epa
+zDMia6Ae/bua772g/xJ9wwFelhTm3N7YvfacxD5mzV+pFns3anxM2NTZxv/DOwC
0R9NXAZX8HFlyooEiX1ZAR9Q8GLYSghMmd8+5UdHWwkAlkOcUajNgWShJv1xzTdB
6Trbwg7S/9fvZm9feUaJiDX6RAiv8ODOfSgkLTwe7xaia9l/hIyTDxq8aqjdxYNc
5oWOnzLF0ui9syTnr0Z5xg+ZvMxaEMbwaw91P+MbubjAeoDt9lR6i+bh6BqPKIkM
8v35c+Cq0VENcFVstJjuR4gLrI2yO6rQ2O0HOQnrTyLQ+2L+TpS+pA9Bq7UlHDE9
eXCEewT9YhlGJLPalsndAYtYXQSnXMzdK3/NlprHKqjU8n02PGS0k0f7qHOZgfP2
Tp3ajrzF9k2Wb5CEDBKpYVBY/aisGw4SVs6K/0j26n/Evlxqrlfh56CQWkDLnKSY
bCyA/kxuW5g5192ogAmlaDNlw8i1T2RYFi7Wnax4XCOJ93q3Fd/SD3b3aL3hwfgZ
XZMxXyDjvG/UON6Lfj4+TmAxLLCoAKWqsNqC/mex6KfCej3lNfHy+xkOAnN2T9rK
ovvRAPZNW/Lv/3mmjKAaHwnao2jFHWAUxTNO/Cj23MHaAJadf2RvZARmOGcA5I61
PcUDrY+dE1g0Owuov6AfQ+5ZFCtPhHZOww/ODTiKqlFfD+h0xAZq891VZdLkqnnE
HDV9aaD3pXblPQnhYz+SJtLwO5VvtaZBXikp32+OnT+YvsBH7IZGiTQ2vAOvmyHT
Pd44MHuMkihsZUsWofuDUMH5zvY1Ss4UaX6TTFOumFd/jivVWOZ+77GvvqGxJAPf
PhNzGnHrdLiF2wyA/yrPtxnYnQ/qhQOCJzQXVC5gzSt1L/zlJw/lSNrpWsUX/wwb
fEUAVEhDxpMoWGmCGhL0q7q+VbiLVZVO70FFc16hqN7Y69CwxlunMC7tlMvj/gaH
MUtuv+htOeCxV9y3w7zzuas8b8N3jrv2wZi1PfTmnRSH8bJb0JFGZEle4yz+f7kh
BM8pCQg+OAwLS/EPXewxRasyIXaamlYNsnbTe9eSbgR5U8ipodUJ2RhgaGBOx263
rRQxOK1StHsUHxAIXudK0fsT1hq1X5/AbrtRUCfaR/ydsU3n6X3KU7jTkw0962oN
Cutr//cGNLXB+AHoBM4a32tbFO1WkUQ88QOWsnZ7avAQEqGHDgIWSYH7f69tNPP8
tndvasli662MFsiUagdduggDpUe+/1D3BTVBL5axFZWkJ1wMWhRBpY1Il/QKHWPw
+Wnmkq68smcZR0WKyRwbYGieIfJrRY13La3MoF14YLo3npF+g/GsRoXrVqzRJ1JY
75sz3e06ovpN7mv0nAZOa0aLPDGmtEBTq0w3oTCr0Z8O6047lWXV5s9z1zfpFwv+
0hPOplekcwjdr4lxX/opUmOyDlrgOeYa7Dy8UHvWgkGAE/LLFvMfbchTDXb2wADv
41UXc3NVr1cHNIjSTUFjY6mELUf9bXbKf9DnsEEsHNzF4a6nerRnjSOMrC9WdEf6
0vxWwJ0Jbdw0Hds0pb8qUpg1cFHxdGda8Cq3c9yhOrnlCyUv7/ZgItSBpQ0d1I97
ze0SyGW5cgatQ+YZ04Iv8sdLB+dHMqPDxfXxi9toEDqMAhSIbdaRPmP0ErJr0xjQ
5HcVbV+5MDSgOjLj+QzFRDUgrjq5RDcOPPOkS3l9BUY0kQaxFkg7l8V7FP/eMFFQ
n5Q0iQW0FNI7g3EeXFGG0UtjBnf6MHbKZII+LzOUbu5SIxlqgPiclTsME5Rw/TgO
+C2zCW78u+2KuBgsaQxYUkohhS6ZZttROtwl2PatIuCpSUmsiXt4ZuJcHoF2lgwb
XP8IrPzlw/1PVg8wzccIL/5epsTjVq0CS5T2U+3E9r3LPaQ6kzkfPHkd45rJ7vzu
PJ/Ey7DxyiPT5Rf1JQ2whpRQ7E7Aj5wlnRo5nKtRoePHS6fXkA9DmoI1Mfb67+JH
hrLSbZ6Bo/WUW65MSsYiED/43xM+Y7FGBxad+VbZm3CZnE43u5dV6zwzdk9ugMVV
HZxRNA/ayaEQpKULmxBvDBSUVGvSSeMwpez0BeqkSzbHL9K2FnlQJMRpWt9n8KW6
p+kHmlVoyz5CQfNazR2vbfi8YS4lQjKSVQuicRL7AMyQH5MNYUS9w2fYD2dlwtkz
nPsHKQNy3pOBpOHs2oujtRvWIKah4MEq+1U4OBpRXFII2gxqLWCUI0PLKgq4LQHJ
v0J95+icLJU3A5wPkdDZQqxiC6LsA87SoklVAjjAywLufyTj8Q4ss/k88a2Uynfe
MqAsGli8EYcALaIbbGZ6GuszbPKS+dZnt+NIacBUqp8HAY3uSg8tKF/erV5wao2f
v/cQ/9DVaVQ8wNL76OsV1dCHDAczotXj1wiidQkNkVFt1rHTs95bKmGT5DNfRrBo
6C+BTGlSgpfYuupiD5QaIJvwgASS5veGqOiePXuW+FgPfdQj0r7Z3Mh5DADH+iI0
Q2BoTAJCQq7YynaSMEl7FYZmJ/lhSmTTcZpyMjHwdEys28mk62tmmlZruNIgY96n
2j0Wsx9+nK+xzHnjzG7j1KeJCom7WT668TypH1rV/9DNg0alqLUgZHS9JVOx9UJ3
KLRAhKXXWPGC/u153G40I3hYP3tsIqQ2SnWhYvoqx/f15vf22nfimneKXM+zTiEJ
aRJ3Y09f0VNBbHpMdHi56vg5uPOVTlVMgNsYihnJ236VbVI/TAXVFemTfkDTkYwL
e0B1840KsxTgLdjoaSv0r9RsWClu0rTlWXW5+9cTWAQOxw1U57wTuymqBc9kiBS5
sQuyqPECXFK835Cs82crR0HASWkBEWgpNzEzlJrf5UdnYgxqtSCoFR45jdk1EiqA
JyRQxDFjdNLPFaMh+inTBvtFPl2IuMfjOyDL829La/fv9UdybubML/OsIDHLCFzi
v+RYwXUudbMH/eAFReiZYD6melgGRe5v2aANxE/SQS02F6L5MVIz+jnSnOTMMoSG
OKnSiT5tfCFQn3ARqE3ZYG1Ob62lXthd6Ap1n4Qvq2Of3fGk4Cgk7UxTuKMyVQ+7
HMNAEzfb/VXKGT60Rk8G66MXMq0hS9JBM2nWRjcRD+knaUxs/9p1N6OwQl2lurWF
HXt0CLX9iwWFFKS/1CQfC1SOC8WCbiueAt5U31A49hBqc44WJ7mgO2ZLnVVUrgmc
QhdNFdz/WP7/9S/qu2kxv1NF5MTVQMIKB8MFQN25OrNp/65KC/e46DKLxZu32gHr
Pu8TgTTfBSLASwAYxLMKoPTPDMV4YDW+C5NW/Qv0Jvqr6vcXSgjb5JXRQo7pZ6c6
0xg/y+6mxFW7zHYnAwOjqNb2vual8WNMHQlb4+PqeuCVVejTO/PMsAOerDQHq4NG
QJ04bmbERb/mMYNNQ2844OO22LnBzjmzT+vcjiRrzbihd87HUdaHee5fKG85kfEu
vM5b6+3uJd7S4cy2L9OLTIGyCZu8oaVviuxJsAIvgJnlQQheBn/tiY0XO8zGp5G/
YcHLC2fkDlTrKcWc319kyuxaOoVYJPTUI3Mu9zf8EgTy9bQQ60WNGz3j4DwU7YWT
UmIe51izfslPl+6m9WPOLmHpd9U4qpYOP9pK4rjXDM2jCYbnOtfajlRtlB/GMKQN
a2xMQY1o0UWPj/Ovu4x12U6p8cp43UWVKTWAAOIXej/H4CQdRsfHNPV4NSiOkwob
wrmf3i1Aca+Bpn9VuO4XlPpdmd68UhZgoruT7xewwSyxGRaE89HiWBcgwVmvbAbd
JJ2HXlL1i42FokTtM5TGRJhMguq0CI7l+uISQ0avfq4cZoMIyL5lGYZEJpguTMZI
BqYsQO+c09x6Xp18sw/dzWHLXJy8wnhLnwJzj6PzaBXRxXtMdece8bU7dmACNdPh
pqxyJKXuyKSWVcL1ww4oJb347vTlKYgBwTnbfvMXXrthVM6PPOi+6R/qE+iLpIf7
bts7ZfwLrULABv5ph+PiTaD5J3p1XFTfU6XnTzzf27DJal9rCP04Rs8O9eprHrCd
U80+13dFbcRup41LbIhzeBbWzOiFZxrJpz2FhmjjtwXtEue/GbJTJADKI4tZraIS
NeJUm8JCsX/ESBO4tS5XlxByKDUkS8QxdcPFvSiPXtr1J132YosFDrOC3zbOhFAa
SafWceeU9D9kA3EWP92KColFGyO5TtRCcSfaasIh6H/dq6idH7JwP9gA3B6DgksS
RECvtENdYxRhY9So4JSWUauDFgXFelbLGYGp8GAOTlP7QbLjZovYEs0sYkb0tsss
ju+A+yg9M7w8prTyZnnUojFs/FRHAWPP1YHIi5Mcvngh9UFjh+2Wtsc/D5v3VrcB
aq5RqmLJW7kpp61wlCuYHXQijJt4RF4Zw4Shs38m4zQY+csD4WqgvF2SzWA+uMnQ
bDk3Kie3FuIHlTT2kNDL2tgo04/J3O6ZT1KCTA0B+WRF6gvDazua0aREC2exudt7
avQAJXYMUjrhVqh/k6AiRtToQnqkMKPRADvjXhNj2xU9D7lZORTpcKMNOco/OjdM
yckbwCLtVHZLfvR0zf/qjKP3Ulp3REJGSRDbGh3oex6m39U4Jat4OkWbgG8e/Oa4
G6fWO+9cPoSjd2ggyx9HDAyOaAzwZZmFnMdXu6cNl1SqY7W8WwSCbtTgYUEbLlmI
EpvvVY70aYePrXk64O9YbBAgA9bSPcOA+vz/b4KZeOg6oYeVF1kyxnQep1hCIk9o
63MQfljxXqrIkZsg4S5tV5nfUqncjOx+Vu6BpA+2n1mUOKK28v/9q+LmwAqoLAWc
t+qt4kLLERjFULst6GywfNRoyOestJmkbfv123dmz9hgR10ed2aolEiMX9rT37er
2kEcNWcnmzqJUr3cpYi4lWc9gUXW0wc0X6ORt5gNFwnzwHW2KDRMiiwRYzT8/hs5
XNedWu7+ZRgjMxIcED5iQ+Uy6FJS72thOA9C2aQJlvksQYWXgJvjICioEGMSBvP4
OKfIS9S7wGiq4ntU5LSqdelBuKVIc8FH+9cFriYSIxB+Yn4vTMeQF69QYYtBNRJn
T0x3Mbb7hciiULnxxxPZ/AaQBzB7DFV84MxFYq8c7kqMun7ezqzs6SssLnhea3ta
vJzxNu1liOSrpjV9ahrc66fyp2Z0JnDY/HyVZ8HKIIe0MbK++sKRoyoALWeXqFvR
Lgo0kzUA89++Qsb4YDoaCVSvKp53cfdnzDlq2kX4HphCtC9e5fjEnbno5deRsStR
CpQWOCKAAZBbJz+uhSYTKFki9lWLKcpwowaLo+Pkp6cdjceUQYFtjEfODvp+qCH2
fjUXBtFVH/XmIhH8Y43RMx2DM76RpOAtTdC4LhrkgIl/j4yDq8JEP+DVSwzpH0mu
enpwEN/ochTjWnwkn2P/B/O/1FWGUHg+kq3sdwnbIOxybjbu2myxt+XUXg03l0HR
FLd5W2TxhtAlDgWGUL0I2htjuq+fZmVwz95ih5jDCLEdwVWQjaUPfspAFBQcAhJ3
fr1djy2F4HJ0Q3nN0G/u6lxOj78M90fnwCiL3ooDdbqT9EuKCVyIq1osGV8ubNXC
7o8QawN658l1vXKn+ukx+/tDdaE9Us34xo9uAJmIEK2q5A134OrQ/fDXaPGTA8nS
O2NDlCj3j2O4vittC2K6MRMs2fWoByX1MxzV0LTQ1S9GA/8Key2082K/7LTfOX4F
SkXS7UwIQDeH24pR7aD2eWBkiCrZLsal2oLb+P994yvkT5YvqwpWghfA0KLXT1KU
YYPkv7nD0LKbWBbkCpBR/tMlg6AREdi69ItWkCYvIXodwg2gJBSxhaf2qWlf2HoC
6o1UA7KN9c4JUb+/RFZB/kTP9Ivs9vIPQSbf6OWZ10/xuGkRjLp4DL7ZX7+9wbXl
pIB4Krn/6xs9+Uh8PtISsQZlgsy2B/5eEN95bp3aiVc2aaK8BEWo8evPyx427nMp
PEg3EeB0P/EuE/mrnqXQ68KtxyXydhjNLJncqDZIw7nsC4DSrXNXIlHq5IZuvaFH
DgUdEvOSXxil5RrDxkfWXsPqMbMeLUmWb94GhOVHBY6mD6nzVv3+afeLSfQH22vM
hQcmJOXF1Bs8eZdoDmTZZarsufM8hgKlZMVQpcCriqamSppF/eZujhLg+ILuTHKF
66PVT08P4Buvg9ZQ7Dsekt9335WNqXxHbL2qVPzzYlYoJyq3f/XHtfOSDAL6U0rX
/1gJSyvyAI9zELu6QkCnV/AAnZ3gh/CcWOsdQrdrRmTKSqCAJcbCG61L7Xoh619a
h3XO0HBbjyMrY5Vi5utyRSBdjD5EzcpEifN+q3XrgKdpVRWdLxe6ZyTc4vLh4ABd
IWgltXOJAqClKGBsTiFxxy4ahQRTwc3pzLm7J4TM+4LBMcGV2ASCYE38bm0cpmwA
F+7vjFyeu2TD0x6W0Cbro61Og5mLy+/emYXQRIkQl9DrXvpOzresL90Er+EAVFIO
EqLn7PqrUj32j9dXiJS1QUBfdBojDDiipD/R/205LCrhWO9VPzgIID51CZqdn8v1
uFDj2sm7HqCYKn7HWekETfBMQvCDdgWdbXDjWqoMoU32Xe/ELwAR8vUvYOXMwzdT
5Hy5TLwS0KC/9KvRorWPl4RixXYkpRZyuVg+TRfhamgpnmtlCIThHze1h7NF1LDx
15GxXSk7kPP2krs5UqAY6Lp7rlNcbLOmOz5NQ+CiBLrDtjJo5KykZwu7kGAPSVAg
nN5PfkHO9tLaHZk8Atk/IYZ0kS2tj8/QUFeV2XbhpO8fW132yqwPde+KxIIfuDia
NWyMmFhBbai3vO27hdg971XHw9ljjdFW7x+pMjnZDcGEl8o2b7RzOURmGpxEW7KH
exBTC0tGMjnUkwiMXTHUTUmA7RWQQGTrEGZz+XBxEKJu+9L+zvDJLd8ZnrfN/XFD
fjynHkRlIDJAYPmiQNZFdoXAMzA/gI4dRwYolkgfevRV17rweW65w5TWPSZML3xN
gNgPB7534/b1obfHTC61zffLpsY5AmZlrntvn2IrePxRUF5a6rCPSp4lNaqTTHCA
5ABK75TnzmX0XaJe8+yEOVDWmh1RjRcvq9Xp9xVo8AgihUls3sNKKZ8q8s7TnvMd
5AMPdtUUVEICXmv0vSJn7W6SpNqu+yyJbeVGOdMcFQnkPqnQ+vkhPp8YNOw7luYc
14aEjlmppxbWFbHUwCOB3tVtjopNr4EMQcSDM/Yv6KANsqQugfwaYGUjJv51yULB
KXRS87XbqCBFCAULVKlPXceTISfh9smpa8ViG6M4B6XidQduYTH/CkjDOfGF7TIb
`protect end_protected