`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 6720 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/59UwEX+aE7FohaWu0/8IpTj7mav863zUNIsgIH2BWb
Abd9opeuBjbGF/waQMI2vMJTwD1ie1YueHc3nSNpEh4OXp8P5ybZFY89uyGz3ztU
W1EsuUnchJoQgbHZ/sLbgtGRgsrAFn+ZoIeGN1d6RAF2wAESJmYP8zw+p00RvjZ5
pBGEHX7wooDexzkaqKS5GwiU4Jg3m2I8/4ahkf3CQVcN8V3jJTt4zVozcjllFZAx
D89J03jg42b8qgTi5NS9ZNGOydaxHBEInQEcoLNJwhdWNYcKXIM4DNkqGc4gm3cj
ZIqVVEx1EvJyy4jN5RMaiRgZH6OFK9PLEHITBa8yx+noFG8wTekirbFtebaFB5NG
qYMdJgy7otqbZ9AmbCCWE6BnUBnR5zwE9fta7znBEMnqbPSwdE3Umi85laL1KbNI
Uv+yM+GhBK3ctyLyilMohSgxfYwMCTL6p0mFY5Wu98dz3Z8ZNY3kLsVxzdObTiqx
V4Q6FPVaSp4oZLwDx7e59AmPOp1PkRt5tn8bt4SgJKT6A7NQRirmxAuSKD9eYg6K
EC+FHNNzt0f9u4o0MgeNEbxuzYAuiK+oZaVH18kaImcUCDdBXykxL+D6xnqmReuC
bcN/H/L+DPmM4HHKfAt3Fpox8FX+exHgFlCK5qmbfzevG5GAbXOWFtiOz5tgL2Vw
AQv7I4v3KftreLfLF0xL9PdrDtTmETW/18AQZ9f7Ubd16QQjne4SqwxMQaWjTG4T
xlZVNFlwdVSlk5p09tV7bhe6Y3Mi+5IEfKFLBACbWkzgyGg9xnkw62Mm+pgjydJr
rMhl++fTARL+HYU3tN1fVouG7diYe53uxbzlvodUdTOR49L2ADKGxV3dLC8ABngP
92KmLUMuy0QouMS248aB9vA6JKd9GtasjRnvVWhZjc1qYZcym0Dc2hZ1UePFmTZx
EBV2mDhtOfiLpnXCrIT9naQsK5lPlCljqvYw0nYmQt6yo7hLZrz6l+/Zdiw9pNNi
HjC7qfO98XrhH+IBUm31zxD1UfPkinMPB6BMtNTO0Xm77haJWE6vBZEq+aeT8cHQ
b1OWWhjra5EOHeEoFW1LblRX6c1YiO/9okVZS1cDJtnuzj0cDlZWMIVTZ5W1UQHz
cJ2MStqBOsc84PoMvpaDinXEhi734F1HTjQdxtCvzrSK2PISPci6EXq1BMc+QBuT
Ptqq4hm8xuRcxfXH7kzJFH+vEejs88bZ28adB9J/dpb+q/lVmBrvYctqFDPSI5pe
hnWqLs6B3Rn3HyOc6z6R1hxAMODuthwTgQy6cAImNuh5mQOWm7pbVF2ETBOGCckE
hc0yWGkXTc2GrB6EvZZ03WgHIUDtJuxKzIOxuyZyHjcbdXbipACwPE5Lgq7w21GL
XkFrMD7z/dhf6NV9daERHF6S7apuVcy04qmW0xaHM7T43bvME8u2y+Yiq3UHC06u
e339kvZreWavGqUVuE3VNsQW0RLMT99obaSrXW+nr/HxWxog/pWbK6hcy4IceX1w
810Wmsm8WYFOjYG2TzveHPC7/pnWI7MooSdL/K7ozfcNO0VrryP/HiAALmPuxq8J
qhPbVLwgOGkQWeSks+vqFjLkvs6/3FD5acHyg5h0l1fB+UFUa5RyJ2TEIYrWum26
WuiHKEEL1fyaD42Xa8sXzY7u2sGBqzbrViuiMviY2fu1kOP7Jz6QPbviq2EzXYC7
vR8WDyYIIKsABjx6+Lh5RRdWyY6+1VZ/yolkTrgvLvCinJqN+xshMmKfiFsFMfQB
xKRdsqC5ZCalqzIN08X9TGfjACLgRFPwMXi1hAM6zr0qeBrSL6t/+wjJGt1jqwd0
Efvw7a7qqZ8zAbLJe/jj4/TpIwGD3Eeu2IfhwMAcfus0HkFHDeOjnyuztGYOhI0+
VL2nOkS45PHzWOnPNxq75lelKe6fp7yr4ECtBMsO1VS5alM5m0wx0GVzL5MA6dE7
sqdltkXhH88f0q3/jXy6P3At1ie2lZJIp8i/VZ5MhVftAx5Gev9hU0EJbhxpOZBK
mnk2UE/xUs8mB5Wu8t65C2ncQ17yinF74rImTwT9cafmyvqHzXHy/5lz2wwucc36
EmBkM3ccn4HCxzSodSweLZU6AaTo4b+XzgyDXnfjr9wciKMRvTYs5VpcO27LuOYr
/XsMJBKPdL9U8TuN/QucYmGE7he9mBXWwNNO0TCk84s+irzZ7z8k8QKPz1LGbF6z
xqUQ4qA2bo3EfN3ziB44KVZ9tEgu8xj3cw3+17RonW0WVq86U3bBLryQnRy/WTh+
aTD9xMO7Wsti977zWLrtgEmRwzEYdVlXpHd2fBHlBHCVq/t8vRBwzhVB6Hi0xLJG
oAPnQ8uyapbgzJRSIOoB3Ow9HR1Di0F21zCMKmL+Ck72SiDJ/GKPuRpZdrmL3KJK
RK3smoZ+zhGuOuOFssuxFror3AkFOgCoNOe/ZAUVyPsh30l26YicaEE/yvNNElYv
ZHvyW0xSM/dpEefd8yuHt9Ea+twE1PArOeAtw/c9vfT5Y6mjY3lBKkJCf5KEZWDR
hcUj4JUz96ugVW+r3OmlyzLQ1eO5s5pNM29bnlGvimCvNvkBhL0j5hmVilfcPa3V
7Fg1wvyae4kSq2laKqJQzBdBPffn8TbL6HKZKJTz1K3mK8OO5Vj5LJWY5mqK0YF9
8RoL6PAL34wjtI9v9gYxmEW88Ex0PFJmFded9UXLWUWENCpS7TzwhHr/dlCXvrFh
4d9BqCSX6U1cUJvXn5ci8Ove5QqLmr9LTyaVpo3WIVs2E8b6OZqpVAP5oPZQuWQ/
hp1oFkXJOTX8r2t423d0elUIPU/S58lGT0oSdFo53yRiaPFyP16jb9wber7lnE2H
EjJ7KvrV8hieM3AGEyKbXTU3swWWPTRO6dhk1G0B9fGUQAmUaM/iHO5aq3FZ7Pw9
nKx6UEGKwl3pSqfJILuBiUMhWuVKTdpBeekMzcwh66XC3OweYEFnO6B2MkG5rq4f
rTEkuPwMZmSDQ7JtpM/pDAWpvd8c/MCUq7BPW1F54pZsB8vYGLtgn0UjCaQ6IJNF
YTZtCzYcrM4RCjH3dcVEiRMofGuXONGfO/AVWyKIonF0F9UAhk+H5Hsr0xyqbmLb
YqhKjbaCs3zwjBaKRDGlKM4TdLuZlFTmLzJwIwUXQZ0ifuenZ76hcRUywYaj2Uv0
A2pJ/WPU/RSpN95gIBPEVknq8kAdVpCJbYX+khOUfKcp+ErIL1dyREzQSbGRYf9v
yKFdMhNJ9hlnBObuscSSw2c5XA5Zd6xjhbChK9evWZj96OonTxRG3Lz52OoK8ZSZ
JL0nSQZjLQKC4OG7R9tmEDl0NBUs1FvUipwFjs8UJfCihYkAcmAX0WkQkjRgGfZ0
xVmaM8ZRvo6NbI0tM7AqR+MvKoqTHeAV+3spHfVr/XLgQW+Vjv+3zdEyorZ6PeyF
Pt1dXokoGAs5E1mCoGO3WJQoiROTA+8SddJSXHe/VzChHzV/ooa25txJUhqHxaQF
xUu6GB8dBZBJ8YVeamhMaINl5M4hY6JxpeAX0J4RRWp4xNJn0ZbYJDXZQ2C4vDb6
20IAD8kq5tLkbqYN8gv1D+PNoafqA7qupd/GhKEymjZG4gNZKJwv8M3U1LsY36tq
iUc7wGox8lGw24gL40ET79emp1FQng2uheZOQu+X2Kn39OWZfwbhiTeSZkR79B9x
1tKDjGliAUPAgiYTaQL5pTPFX7jgWPFX69NdcttLuh67tIY2/a0uf8jHwhS7iIeD
j4l1cDGp7Gt73OL+CwCVff5erKiGnyAQn1dUJaJUiNcyaDo2vVfrC49MhYtiaxRz
kXW3q+RVoMljCXqFVngV6YljRfLoddt6pYA77ms8g0nHZ05Kp6ZA0+b46n0trZgQ
gUmTt7421nICx85ZkfG4GXOcyTY1LnEEmAq/JSKXTQ5mJJj01bxX7Hug8f5ZTueM
tRV2ZVIzwBK3TTMmc2x5NixbYW/PzK2ikRb9/UGSn+1orf5cR9cYb4jrEu9r/0q/
XWcoxrBnlmMIB8ignVnk2jLxbK+o3TYvuflh9Qug4k4Nt7pmsluqJ2ksVnVLLVJm
2XycskIKlNQxcTaEfEoCM9RcdobcH9FLLc/0fgtJ02+GPklq/Ug08AgJQbbM1hFg
sN3CWg57YJOdVFW+Gu+HomtugkVLBSLO//5Sl+22Nhs6wQIA58HwqLfBVOhUYXGm
KM3lysO3+0XuXALsCvJVKN8PU9RnwSqWI8lD0Ft1eJnPOGA7nQOeaoZOWDywMlIf
8fI/Kncc4ZhYqTl0CQG7YQr7XWDoFJSQUBj12qVRhW6XQohjnWFqCzV6f6ZDo7gG
skJu7G4+4ATwM6HEknt7UrHZt2lReYud2t9LriO2n0w0R/l5FlPf+2gf0OX88/Cw
EzNaWVfy+URLQL1orZ/Vuw+yn2bvT4CxOTRPo0B7f/GDEFdXUnlPn4bxxAA5aRdI
aAO9D9vtmJqhizy6o6WRSEoDnkWKBye1SZjERckMQp9xyfJY+fyk4cWnV94Mu34W
qhajnPMrse77Il++AEpxEBBo84ALrMNYB2F4UnQuUM9828QHYcTbF/6HwWCoBYQF
lXDUSAi4rvJYbCusx435D4rmrOWdFLFNX14hMxx+N5FaTJe0XJjhxMsYITG3591i
2IB3nvRUfwUfKk4bV0/Ouuvv+z+idjPzhfZRvdXKqHdywX3eerTIxzQ7OPUeBb+6
KHX/BLXWrEXccveNF7CwsqbzQtioW/CzsFvafJD2Bf4oe2kGMNfR816HolYqESy8
JwoWL5m23th2wsxYX+6NbCbxEy+9DBAJsCg41Ase4snOf7sBwZdXHYpdtBaZeC2l
C9xWVIZHtXLnRHdxIkr5xymKF3+BrlxC4HihZKN4Ckc/T9+tEmj0PkYTDVRnasyk
Kk94cRC03zNaRm+72v5odTUSBljJXXDGxTwk1VtNi8++UCTw7+kpM8HEmNufBsii
Mk3KalBhDG1/3COZ5dqZ5GOmnmcr8q5WJ06nFLRSdzNtr2uWqKJ4ECbGi9D0ocOn
c9a8tkIE6Kks24iQxTPwpsgzIeFIu70D4wyCIMqtVAJTwU0N79O02OF8GSaQ/D++
Q20Ul46wjm3Ob4PIpDp5jjdSslwivPEGG0EBcL6+P7LLw73YHg9LmlYd3ThflT/0
2HMNniU4A4bdufN49mhs67yha4R+j0ay0hKnM5C7BWTRCoI91MN/9C0OwCjXeQN9
juG5HoXbBb/yvPIyuTke+g5RS0l+NqvL8i/SZr3YWaDhsqWbN6f2LnHGHszDVFTu
67yjb+4+adQNEeRHahZtyMbSDJCsHKp4f47bUnPWVgj88YNVY/AguH5nWQUfhvMq
HgWNuCCL+SAZ9GW8mCoq2twAGJEHJorzUdMG9Ud8jyCHnx0c3+LzA6uqiQ5q6xbC
I+9m+BUnK2RL5o0kcGK92OJPSjPCIwzjZ/Fi8cEiT4WexRCSqsmJYHzrG4vNFn0C
c3RgcFkyO4haPVLDO01LEmDB/fsZrDnGB7Oiyt2ljVkbN+dGDZQ9MPydlHaOhSsg
WCZDbwo7EvVJxVB4/VbqCgXHofoOn2S1fFi+k6fMs3ox4dv8/wsFCiHYmD0zzQ0k
bc605jB+dPS1H9rp4DMJU24kVwk2OWXFuiWbN/IN9z3dthgYFlpJOKstrdzHSNqw
dnUzQzzRF87w3xutoLGsZ9nz1Bc3Rhn85SHpgQ3attDMBe3WR4om1/hJNfK/iOjl
cSSyMNyUvWm4rj8IcTUEKAMtdyiusVvlJqGv5twanx8IdkqzS9lcooV4DqRPCEkm
xtXJ4n/Ky+EjsNHQo8a30iSCGJClm92/BHmHAqSoAuJjRIUlYMmB8vovt9Onw2Xc
97rIjQKD/92RbVaJS5NxZY30I6LRKsZzGdNL3qINgSzfID7/dN3UrWZ3zbgED0gY
D09197ZY4FDlu5VjNTfhYF36kkDOtJMdC4KbvMqAEKpwHcv+8lwIYtbP4XYS14G0
nhw0XNMRRgalGlznqdEEebc2CkSCULHAAc7nIDdwdseEt4M43mHL3glOQUVR7e7k
JpblQgO80m3irI1X/7uw6mDQDhWMT3eJq9OeI87Sd2Dqk//vlkqtr/qEau4f65yF
gpiM8AhW0+ZSg4EiWTZL2NcdJl9SxmqltnzTeS8+iyWarCmdzWIm4abDn67ZROdz
+oVdWbhR03LikJFWfLU6uvcQyqrgmb6gUVW/3Uy2yhAkL72/A3q/FgMTU3z7WQVL
QB1VLtasK7sT5PWsxwT9708ngkbhxdi1Wsp/SDZJyhqhBgSE11rCQ4VhU+RYoPYs
JqLrE2ysAbvA5UaUw5pdnOHLSb+U93cObL4nwi2JFVYpTWxGfyvbN67+YB8TXSA+
qHnAESA5TY9iWM4hPz+90ZbZTN3uJ1Fh2BWJdTF3HxVyCI4smlVOZE5ar/C7FqGb
/Bl4W0AuW1tfUZL6gFWgp7V21QF2l3ruLT2r0/fiOupHh9p3RPq2j/O4dKBPbTN3
hDvHwEsYCyspkWxXN0hrJSBdvlM4v1xuY3wk8wZm0oBK33/n8vE5jEc+neQqSl/5
owdL05sL9PR5zqiT7fj6s22/6asTXO+nntWPBS3mAQlXHxjDlUUVr/cMkZF32t0D
9N6X+jZChSvrJfV5/JGgra4dhAcHJfIkpcVCTjreHkYpOCwQQGnUlV9F+eWkfBfV
308/A9Uw+uH0mFPiIlLTgZ344WF/daMeH5igzglspDAVe31eSyqB/frGsh42GfMl
Mse0ommaNIo6VlkruatsN56qXmSRYKcm+zEACw5cmTmWPldFHtUgHaYoV/TYdPPw
6XNBgkWHr+m48so0ndE5sG6rLuBjBWN+JTCE7QN4wFXGU6W0MPT6+BUNi6Mt2tfT
a/Km+GU7wusXCJOjg9BqIcSAsNKIZNTBoSY8QYf4vLtfQeQ/bqR8lrrtyxVWeNrJ
HedBds4w5fvd5oM49BvZVQQOcgoa8LZgtfCfhyTXstvdSuXYyEZwYyF6tw+1vLiJ
wD5SNgY5n/8ra4OrVtMj8/hF8U0nR0r+ghuMqXsxZmzfJpb/fQz1Jo62jLTGxPT3
wnLgGXf+F+YDAoXedLaJjm7k1kKhq+EJTKMpy84MZUR7Viut4H+162URYmQdgpcw
72OUPUe7TemcL1r7fJ8zk1iOqVTsYUSJ4USln2JNjP6KUrI+d8R8tcj5Z81SX15O
SZ84AmSNeu/Cp1WpHrBd73fMTA7VfDnXV3cCl2Kd/laCfYWp+10tAbgVogLRCZIT
RU8R5Y3FlOw9I2dM6zYoJW2la74EuQn6a+o9FcJpPEk9Pw7mKgqzwMoiO0VIwWbQ
a0k/Ut9W8mGQvlib0xBvqzaZhZPiN7fknj/fyHlyAclg+t6m+onTpMnf1+aFW8tA
FKRm4c/yMRSXFx1TGz42Kvb9nupwJUAdr7p32FFVzSAAi5GgeriUOELhjTePGaib
aw8A9t2n0UdZwXQHm2uQ/OTc/yH2A7Xy9J8AZYiTiEWSGrehncMpHfPb8AaxtV0m
NZr5DshfOpXZMs9XGiTUOwatpH2gNsUGNkwVnfDaraDpCoi1gXvvKqwicBEI2EhB
2yUzjZ6m+Xo392P2MrmF84i3dw4QaCOvy/QXaekOu+azzIMHLcGLHyovQ/GyqdmR
ahJ919muxYL7Gv4XzPi8Gt6BSNJAyF3JIB9c7BednhcokpnE/o1WzDUjm3IK9xLg
/Ze6VLb2u8itUfTH+ldOHbccLvAZem1epZgwxIUxuxMIHjIbHjl2tZqAfgwbWwDa
FPJ8J2cy1nI8V1Lc5Ugt2o6LR3yVwjTqB4WMox+b8+5fiPecpDzhncLjMcE4tOV1
1mCn37lA326MyI5firtb5m4VDjGV0EzU21snwD73QRjzHyK1Gk8K53/r8Sx8wHAb
Grh0WXvPQzBpWP2GNpiKdRnik24YvoKM6/UFNc13K8IWe0cdTUL7+r67MajjJo5h
2Hvxq386iGDYf4YCquXGEsj3N1QE3toiEee4biZmCMYoG4w/k1jH78veLzPeTqE2
QBWeU98Q5YzM/4PN3iPmkLUEDMFcg773iIA25A93Ys4RByRDbjn7gmbASM8jSvf/
EBJgW6NCMLcBd1DV1AK7W6a5RYLOZ45oNfr9G9Z6mA1h6Ht/9GNTxpETKB0Gfmg8
3edZ8e5altDM/B3iU0zVOypDAzjJOshXWWBZ1W7QuqX8zV/8+Ou4MznKON9ZJkev
ufJM1kdntNccpPMRaxqWanllpJ5EQ9OX/TkVVGxkVn5wt3+9WsavqeIl4UxIwfmW
U0LntvRn8hbDJsKSxoGcxrlZq5u+Z481HIq5/Jc2O3oucBhi8faaw22w5KleJW9L
9+pbSHLVJ9YukwuwfO2qelFRlTOVXf0mpCTuBonH4VN/5Hb4uOFqPUKGEU6rOSI2
UZ7KsvkvotjQ+BztR89fWcp4ZweWqEPuITYZ3nXPLgLqtk+psCkaW7tUyzvyzThp
pfN1xXTylRhmaUVmHl7G3tNw6KqKH3+d530VfboFbXqZ7H73vHxpKll4HmHlLi93
HLKK4QIAHzaGZyqHQuRaq4nIE36RewDK70rXqbhpTJvSjJ+Yz9MjAf5xj8LelyMv
8lYHM/tRn3T5FmJYIoMEZlTm0qyZdr7zUFyCoHSsSw/HXuOS4s/WoaS9/Svd4Y6X
cak4zEGDrNE4ZCM3v5HYpWMuHTpUK4xV+XhFAhNhB4nL3CtIA/Gy7oTeqP4mxT8/
Oogs/9rtheDz4qka2lyk87RnBXu1cMKW/A4YLZn4hfDe9DrFVbBF0oRGhYuIpnWr
OdC/PRL4Qh4kM86ggma6Ii4qf4lockSX4a6fl/odmJjTmuyBnaivYxP1mIeW1z8g
LAR/bnCN629fjf1fq+QcMChhqHHbOuo1pnDPFrethEzcU/tV3aFdTgVhD41oWNzS
`protect end_protected