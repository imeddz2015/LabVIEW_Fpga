`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 15456 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/9huKRhRMtvnNqb3Z+UU7TahEoHV+T8U3P3ufru7l1O
3DlgtZzb9QxCbOjthp9+wDkjygH0eUfDrEl1ovhZG62FdHaxW4291aDlGrJD7R/g
emfroTsHLU8ELCedAOTvD0d3CYBsXg8HLMSLRpkDA+f1rexRvcWtlpnobBKxEsRD
49ciCA2ISZZ4wzeoj0PVbqzboFs/GX/t4BYHJRPIiT9VPenZ0pGsGmOXaD0X8e6U
pQyz3DdO37HdYGF4RiUoZ5bt/pfc5xeojFy0Td3QJ6aNmA+U6wlqL014gAGsUxsz
+b2728Q511e1RJE87/6YCrmSN3gOTjnX/guF6HqL8st4lwndbjvcP57l1+de88Ev
mEpv3IleayBPvj3J85Ds3bRZjfIE5ZTVj79wvb1XR898cMwLTkhjeMoVWN9M1wIn
MzaSqKPIs9MUTpdWPn4iDGdEflG/+pJGkrSp4reFkp8/NgLxfWkuj1ktW9wm0SMs
qp7SR7Wh3Ss7fDBhrANfuKI/uso0Xox9T7DT9u+nDrt+fcD82jKH7hKcGV90uLXw
RWfnl8mZYySmCZJS8T//QQfbwBvcNMgmsX9FL4k9EtcGNlqXas3G9C3jBPcOPI4Z
G9rqRVJJZ4c4QvCWH+rmCSU5Ar7AX0ETCr+OfAFN7IPNnfNQWXzcfwjSL8LwlC1u
48qCl7UuDt2gpxC35QUjr+dGfwJ1Fr+A4NTA+vf7eWiSofG9kdtreDMVUEzREH//
OjVGTBsB6YyYKwNrxaXPbvWTVb+kV9roQ+p62m2euz8bxKdCDyH9IKrzEgF15YUM
Plad3LZR1SzKn35R9NdrT1DsShkaeebyP2e5G15qx2bfoKjs+mhwogjKGEBgCTLS
dw2j2RX54zLQW9tvLkTy5ldRW1Oi105WqAHfiudzKOoWsUmG46Ov2uNDyToAJYv5
VZpg2ZKF1qo5NY5IFUcujFuON6GsjEL0Ge1ckdXFlth+yI1J5Xj9d9CScsSi5GeN
HRuYUXtObI0t13CqWPau7zqA5Wan0We9pYmKzaghu7g/8gkW5ViVXHhu9eYSyurD
YCXudyQBY6mZviwPYkVIXr5x9txp1upGsJA/IjhHqk/Eynef/1t124BYOyX6gn3i
ioZtdT8om2a7bJI8qFuXwGW4DKqYi8BWVvqDWp1GnrlqGoXqGO5DgnlaVY4LFZd8
BZDkB5q7P21YzoTymheZPOxjDgTiDccE/XsXGwvKe4KgwMgqnNdxima4ElZUvyI5
sfAOCHbohIgpU7nhfthKP+ghH1jHiOg03AIprIeVW4oeEyj05aR835Fs9kv71/OB
XvtQhN+r0IXZG3TJT4BjqgzdLgT9jd5T3j6qdIvyNX4QIVgiVzMd06GiRMR/+CM+
CtAF/CETmSKxJ3MJhMUzk+tQw5wSXsdDZhtpaZT6Ty0RR7kyxq0+L7vDl2EJHsF7
s1Hs9exdVhhVb/tqbYsD7aYDbkGqyUljk73AyR+S9Au2qlHYR0Z76RO+/OJY9irX
VHoLhqs5QkYDgXpPcj/JDKZdptFic+rMBn5NgnCoJLYw5VZ9kQCuXMQqyxNQbl3+
iQzVzSto8IQt656+zTk44VuLJiC1ljvjBnGDGiJJUHEW6bRwUcLy2WUkbTkb8/RO
3oLT0DnfBa7Y4WYz6vHxgzpRZ8vNqMQ8tiaZ+d0BL93Fc/MDMhi9fI7vmfImW0pl
VTlj85w/PpXA6L/F3Y/W9KZUUdxk9juk5fEkopYuTkKFphx43T0Kvg+oizKOsnA+
ZDDYrtQIZqQ029XpunvEx9Qt0uWvUDTA+8w1JyE/pl5hkaL4h/bDNRTC/YeCyFja
hulIaEfY2L7On9O2nSazzSsNGcCKDEULRayrvkfqvBIEoPvTD5Oe8Q8VATai8O4a
S1aDYIjQwbnSvF7pDKQ6XCsKqblwHIPJT7kFqAOR7PqRfCkHsQpRYMgsPhTTKtJ+
x3LQUs0hwu/NlgmGxgiMcFhGT3+NyHPZCjaHvvrGdP12gG9bDJeCbBGCM9D++6Vb
I2uiELRx9aFImCF39IbFrHf0aAvfVRy7B5ETk84+k/tYU3luOHLX/a4/rpHPON/Z
vcG2MEwX7S0CYqHMYSZFjHJnw8kQPgUQkdSeuyiuC4XqWpDo8hYOGt7lyXoJdIN5
jC6TiqlWOP4uwU4Ogg4glEAx0X1FRgN1/PFmogYTpqlNRlsY/+j1qKp0Hd7daRK1
TmtRsFfPM010ERyyPseVZWhHQ0ld5Z8jQC66b4EHy4ceBoPIaeD/NDSFqyxdEm8j
Y38IS9EbwicUtbS8iqEo7PxUexf2X0X87vbcm5y3l3ddTpREvz2Bmr7ha7DgH/nd
CLdOGyV/VKMSU2QaLiXwZAYLejMkkIHsc/mUQOF7wvD8apIxtvCaj7scMHyLOSFL
/CaY7tNKLY+CWbZ6PRQt58uc/VUPR3AamH4jCI5bg+SyV5Z0rQGhkhQmYD9+5JLW
PlpwjaA6swwXRsYPkju0e68/yFqcAATTrmJD8kcXHJmaOwI0b3k3j+KRlt+Tqpsu
7hrQWk5w+1W8uIwiPEwhmttuyl1maUPae2ryQzfoFhhZzG87y4ay6GCfRtrVARlF
Laug6X4xxoUUKJlMalB+aLyTSKIcJsUa4EseUbRqD8mcNNYOeVwbCsySykNA4gIW
ePdbs7tuW7eNPnF/pXQCvjGNqcTUwalAwBXKb5cD61rFXA3HFU3jm2qd0do4p4po
+WpoGEpn6edxR573WU7JOMOvJL+YC29fo93TBrY2V69p4b3Tt9gPtE3LUlFhOjlv
Ybc3ZFeQXBG0KFtmMnQSsay0lQn8DgSkgWb0V9NmEY8DGyAkO8sY/2oSo/APY+dE
1rgeFjKt09fUkMBX01/3xmKVMBMJN6BqIg5sUuI7pY4eMjQ0YEAt1ncVpCZCb3dV
okMw5sQFy43950e/E5y356hRsIiQ2YiTlH7LCfjPXg0vFhtsMX50w2hJGXViEe9B
Ylr+0qOHdZ2XgDnzQSGPNFikgR3oOcYKryxHeyf4p9SdZ6iyro/lF8LZ2uOFfyBB
fY4QP+eMI9UpIUdWx3FDYuOjsbAF7BS79nEYC6TmIWVC1zMkdP1Ag0zfALfjCXLW
BWRRH1Ijo5zXj58vTRH3hrFb6akbWee/1HD+vQbryNklGRclnZix1AcQMsMyc/bw
sNfiYC3JwVirtPFHQsO1AGJwE2lB33XUVMUIJy16GoH8Z1AsrlR+QkPYoLnV8J1v
gav/yjYp9Kj9na8WdWABuEun0LrmGrTg5wq9y9VZlbqMjcO+znyU9MeqZ5SlvB9C
WIpy2QH9uOUbjkvlkgPY9TlJ5B2/suXzlWZOQ8Vt27Qd+zkjU0nGZZwRrd3hs2LT
UA67pdzgvC65apT4TxjGk2mSayn2FNwpkOKWwbE3WIhx3Sb5Z/zRdYL6+eJxWUFl
YSjo7cGhxfMdt2oF/bFNciA0Gp7czZKeY4O+WcDAzkcacGJyTtzSHlyofgMxYD9Y
DUoiyzedm8+il20xzOv98UrB6IpT2MJMhXoZbPfglr6QvEteoCDoEYvx2v7ZKkUD
8EAikWU4uiQ56UYpqGxHaAd9kXGCEoA3cVghHdoxrU98XeJoEUfUr1VN4Fq53YY1
s1YktYHGuspRNpoJ+0e7j83Vw2zlLBFpj2ho4qCKzJ5vMHChoAlUh26zgR/jQI3k
M9ilsi++f75w5qYr7jtpBTCnSJPwQdxrD56xNHU23vzk7v6GX68cOBnQQKQS+qgV
7vhx+5YidyvvQADjsjLy5qBEhP/C95+16/v6nUrg7yAT1Ey93RohP2KjzMD1xDSo
KUP5Gp1RA4w7MtekZ+2SdcOe6Zul+/1d5SuHaJ+OWSiUfDcVMYILpJ1gnrzSyx1F
YJr/B121xHRxv50XBKfpJ+gcCnttSHbjYWCdVZE9nQ6clFIyVEiUDag4nIyvTznS
28bdV33QoxlKkuuDld0f3zn1o5zkgCa1tW6auw3yY9iEO9J9TRJ9oUJNGOgFPf94
6Sx8zN1xZCUMskyQp2XyIFuNgtTR9khXm2TjVO25F8hixQenuaRPSWDsJS5N4T3d
xdWSBngaiRPNpi7lHX9gKKp7otBUI+lMzrUMVCELAnanv99NvzwJe360wm0Y292A
1UOeISPWtlOUBkoj4U93/cHu03XVGE9u2sHAxJI4ihzn2FCzBnyqD1JNX0H8Vidu
M4o6I+o6BJEoW1NQqI3rQhcleV9bn7VkL7IGGPSOSIpQP5VIGFZBRQLJ8qF3GLyI
wHTz9SgxXiA9MJ0qg0lkQFMDaOJ3ONaruUw73hDedQOXY+38z6niVOUvv1ELBJQM
kYj3TqWXrPBpKOstpjYvWfOTdMLtSp4CrRszAbNbIcOzksREzTCqMXiVYl8hkUp/
X0Kd6Rq7o7bv9S20TnTbjesqaJvd90oLLzLMHRj7TzKpyumSTTDZhunrbP5RcxNq
JMGvXhCP2oov5D8GPjoshWxMj+U2eKDJkRC8cJJWwaVkG2if/lRfin1Yuzk9D08d
DKv8ntRcCxiVkp+kBfJfekZ4jSVceh8n3Omq6BBjwXyziMjdlBqfhrZOOc82E9ZU
uMp24YbQWgvcUyzOx8z5tIKAjlu3/cVjzyCSS+JVZph3Xnc75eXkvZOleb1PVPOJ
Kc/XLJxmG7txapoixm6bQBE2+XkUVvpDuIYHM5mVqyaAFYSzKKx7ovhXocK7OYF1
KCZPkMp3LLYDDdwVSweogM5hnMRUULReC7CqH9s606CF3EbG4XXdzs9ijCDVvK6C
+GngOOkheCQv2KJ67nxUS4XoAnvrKKLCoA1ebxqeCQO17cD7dMfF7GojxddCPDJv
53X69n+F6yoDv1IPRKXrosGmJB294OFb1FD43I6wKZ6IfwQFICQT4mY1I9LoG8Zq
VepaC9lkcjP2G4i9Dzq2ijOn0+Pgkg3xE2nmDiM92nexWn1zgvYuFoGCJovLj1aJ
LQchsRFJmKfgV1JP6BQq7IcpKYeZdXU57V0CdRjMKPe4WX0BTgp9cn+WvzuJFtyc
oaP5F2GW/FZIGZY07Ey56kVkjssnfXoEufH0VNawCH5wREepO6KwZBq2kzOGyrEA
KzTZwEIx8XgO80YV0Z58iy0zkXiqhvDOXsUbLk0cRoG2BY2We5AdrndfIunU+P4X
Zb1dBin31bCZrnHBpC5foL/tJfsHO6EuacyKYaOFvgKTc/oBRLLiXBMuEFQDduXf
1+6NYm54HQ6aXoHRe4E5Su51pS38edSXPSCNQnoPl7seGYvz3mDFIVTdPgx8o2GD
pVMTILR89/98uaR9OM1huKfAW5NAdpNbfqpxU2bEbE4o66mDAuOxukzMCycMQpMl
mJgbzgzKuTdNG5y3cZCylmeRhiuDH4T7R0zO/EXU8SQDpMGX4DBz/FhS+tfXpydK
y2GMw7sayFiHHca7uz4TGN/MkgCasm9EDVM4G81mbvDF2apzH/xeJTxh5kxPKMHN
9yFO9Mvu9wvv0eag2nHhfRpdAq5D0DYleR38T2UNFjjRMw3sRhhZOzlaKF8Od0l7
JKlzmpzWsbYQizwZn0ptin5HDS8d5e1T7LmGdhYYe5G0ZPjG2jbSgPLcK0JyQpKU
pIfRX37BqbvXBYaZV3waj/5xcxoETLCK7IDvh0q7LbgfqBAgdUsR+JzGOIAn0s14
2e40aEVoaKI7d1hACa2578/gtrjY+nC/hNTuP7xalxXLg+qPCuc1CBPWiIYugEu9
CA7j2eUQT5DVRGDKD/HAmEACPkfkWJUMtd93+MAq2UzG6LO4sIbzt2WE+Spjj6WH
sNTU6g/H8qbkWtIOp0d2B3B8BkS45Mq9hfObLg/mdlOlu5SgPqF/Kq6UHvqSkfWH
pUUJcrYypVxpKOGGxIRWYGxh0FjWq9vV+StutBLUOFSJYGp0OLCmZIUy6fY0m5a1
HroAoI/DX6lmi4VaIQSNi1M3vgiUAz+WUxZ4llXzwPBnx6Dv2bFDRKzHsRDOljuw
N2nKHldftB8+bLp0Y76OJ4kbXZEAbqFhQx9YPUYCwF96Rl3fCO5w8U6RRTLE/zYl
mnnRGfNYK5suxIWoAyIGoCE+daxLcuoU9LwPcrCoF+1ZtCgasPFtALdcRY22I0Sb
LbhWv3wUeM0DdUCuOUKuSZBgscODGavrr83985SsYlDejgbG957udH0AWuasfyIw
M41dITor4lsWDrJPzu9p5D7GZ91vPnYLWUHj7PmDM+VJaFhCPKtxIWU/HUiUmfRc
6OTkpjFBALd96q1KzD3xG1XW7tGcCkXKEJD8aOab8BM2SMz2WcxHhW0bh9f0tMhw
CcOopYvX/bzHlI9BzrqVlp3/IxN4HfCLLQ2b24ftEF+C+WjqtYcR8cTMGegVSpiD
rPTWyN118qOTevG15NEIEVdO6W4YzRDyUZpYUagITKknVSKZk3pzDBa2OWpVIeEn
boQgXg/PXOu+Ac8qe9qQRK5FmrlKoajZzV2kMT4Mjlk96ADXP2uf6oLX152M49g6
ym3UCJmXRQ3UMlrBUTMk0XMGxnJ5TCpQTUJoe2yCpCseBVdh0oiyuhWLMraZkVgj
/MnrFiTbhbRKWC/PJ57IXpAuefoQaxK+oIYLVj2soPMxsDOmSoSZPSlNE5dJ4yms
v8q3LOqACyq7uJwgfzysjrU2TnC8aAbOYPaLM9PUpljLs5Fnu7ooHoqRMmqFbN8k
tZq+GyBIDPOzaZkSkUbskb61kl0xU0kkJcrVMyVgDjaiSbUKTnegxAteCvP24x/4
NHYjkwU+QPnCrMJ88IiSbUsCJWXz/tXWzYo24rtpYXJcJmoR6gikdaYALRRe7SZa
fdkyz5F8sBCNlmETDmwR8SUyzSD3mNqbHEd3Gnc7FB/jLWPbF4LnQvqalXOCW/ke
PCHkmkKQ1YPn5w4EYg2fPA7clwDLikamzbbjhWiFQRiPVLaRZOkqauu1x/TEREfR
0o/CiSLFFRP/iMt9MZPcr2ECFbMNTEulQb7MwAP78+UWfMYaCitwRHPZyoywHGVo
jbFzAiJbQA576/TOoauGIXRivtgY29925BHLMlm2yg4lm2+0F1EJYzgiUU0cZr1w
E3QXJdIT/wUgRbIsa8C1G4gIvxTUpA49ArDLdcJSsp0tfBvh4dwBW2N/TOOL9pBw
vw5uqpaV4a38vl3MA2aeC/55L5eDDg4PUF2yLEpiKudNiWXfmNygsIeU6YE2d4ji
GTMwCZ2qEK9LHtuNZ/KlkvwYi7fdX7gAY/ntguuWe1LX0yK/vA1YOazbgz5EYXPV
STledOnLEJZ/DYCFczi8nqPxYbim9EiQUbQdoY6jPtYvyJIk4PrVC275kUU4mH+C
FfZz5Sl/tUokPEIh7dCKgSNJD3Y0vbwFhQ5dA4iMBMx6KnoSS4zBJRHz5fR18oT3
Oe50GfVlo7GejCO3eUqinD7scP4Mr9qxBOd6mYEdETmzQZcQaSQpLhCZ4GDdfaMV
iWEr4s/VYC+MQx7HHBhB28fnpsj013PxAsjeXoX1oCz/zv5KevoBRTyf2Et7mopV
H1fA5aPyJKCHOijN0kcJywBY8QvdmJRsW7griXFAMLyYBUSebecLucO208sdBGVo
CJzlJPmJOttIWINPTnhShar+e7ZV7c9NGxg4HHxRKVEZQvmtOxMQVyb+oW40/7MJ
RlPs+dr+/rMnp6Mrxjs2Hzh6uuv4TsVkKfzhNB/fWhl08GMmo10sgvgd0lTp9ote
eram75EMvHeCowb4tOYynCSnArLXRrMG2M4vTxmgHsKDjeTpPRGteB8VmHfY01Yy
ycsmblR8OoxD82cYENNEgsynjM3OAaC681GGudypg2ahbxrx36uRBY8LMslyRmtF
PpfD1tTRbHHG6FuVaEo1O5lYrZQ83gv6Th10I4maBmIVB2wB2vSLbjgJ0zB/udzG
noRfG0kumw4PofboNxvtp6GZSYfdMG/eTH/5OdesA3+x6j9hoizxPg733RQSVC0f
Bqh4KMHOd0qg1gIFVmwQDz3DxVDU7ptUwDvfq6TGIqRtFh46UlrPoRXvFsmXwzvv
8JY02XKumHlbPfq0fk24FpwqJVFyHEqNVi0TxIg5eyUd/e53ZW4r51cxdnrpmXlk
6LhEnjTk6eu1KhFH5nx+37Z+PPPeEgHTNOQdgyav+vQhS5v59D1dZvi1BRP2s8Ly
oiDwZ1b4UdNVe8ezGZlilAqMvA5fdhY2uPX5sBxV4oWFA9+ooeRFnvmzQklBFIbv
xwJtoeQuwcFM01AXWEA9fH9YsILf9CYuzLDgQxjlslCnsm+VeLh36TtxVHgHxlE8
wfBmw4RUNouyubQOYmRoGjFcxvE6P0ihtz+GzwENE1ZUeWid0G4tyt8gexqmRRx0
Uc394a6zZ2YF28SYN3Q5rKdIXNO7zFDQCQT84zQfh1D3ey39Fnn5FUTRpURqF+kg
JSxCj7MVZ3sC5zTYQXpD7i6sFhMgFhgAF+Hp2ZKcmyExhscZ84+vWnjNUVUa+K7L
/QxsSYQnB5WD4b6z6uKWHqRLJAsDHU4E/GARsdWJsovw01+kxE8OJBGBXcbjDUkI
BGcCA7719s0Ks++5QcO3XaTjnvf/hS6XJtUmYHTVTvlp6VkMU1wWotEZiV7aWMX+
VrNLi3fMrZm8VLTV480Xjx8s+QeJrkOkFpVS019hzQ+zHTcOr7UWIULb+ymfHg3j
ojcw46zeWElaifPvbu+w5PK9g3hM2XBSPWrkjdpHxDmX3/9DgONZOcSMfjwlNc3R
TqCSRmNz6ZVtu2W7LB6Aoc0XIqBsLa4Uv8R3hAwHmpuonBnVyWdrnsG2NLKwDYRx
/w0iTuPysm5oBcdlR+NS7SBKEivu3tNqXUrlvl9jdDk2ETcblh31zHuXj+R/2wnZ
QFjNms/dyT1AEFr8cqQE+IZV/2PFCH1Az0XU9gKr9sVDUV79NeWmwDq6ofNsz9uY
cuvHYqTYxNG9TN+z+mmh4cpEIR0aaISBcOkk+eh7B4ugdxGVsMo17sJUUZ/ZGCsx
dj6DppHOS/XfwWswobmytYerIQVTGa/Mv55vR8klg6vTLGAAkoL8V+1+YDyEODRX
frowNTrJio++OBxiX2UALDA8aEUkknkl1PQUFjDHNA2NxkGAJnVFEj62IRkGebkl
BzQZhObR+Wf/k2Uul0smd1TUVeRGuhCFnwMQ5Nc3H1SehJnEDkJ/5OSE8MjwbKR5
u+72w4C6kmFtHt9/DoJetoZRsjIQe1rrsAfoBKm4qou59CSlOa0ZgUAPhLYXp06e
qFaMN7yCrZfoc+sniH39FVM6QjDrgYugweuktIbzHm8bBg4OixvzDYAIfrKVwyVk
kJsK7gr9Umn4LBjiHERkGbQFMfzyFy+2dE4IV+8pCokzal6sr5e2aOlGrOnXz6fR
UsFr0R8RHwb8q/BfNGi9wJ3DkMbfsHTj8wayXd1IPm1EraT121Z2ambyddsb8lki
STcv31fDo8Ik/AX1bdQbgDNcJLLRVwlk4G2q0x9wyLoE51ux3vcgvKAkddL8s2E9
Ru41aUEESqQ7MLKrhmcNzaxaBiXNAw1zWX+1LumQFfwCM+3J2+sgciHgZJ4B5Bl2
a0TDj/1p6UbrvP2Gj9wAdggMaRX/+UzjEq7qpabTXHrFyPBdFw85W6rLsUL8kbZn
OtRUItE8QpB8JbNB8MmpDzjRFFIIaY+LdPTyh/qPlnpskgbGc4h9EScVEHk+FKcE
2zqn7DQTggTaC57qTYjgpn9yOg8qsHnf8a24R1JNlRfPNKw8errGGkjiKr4QF/Iw
prxJVW32D2WwT9SF27lhvAu3UB7aTTqYSB3btSEAVb7R5JpvzSx/LoYLPzjyWKWK
qyfnv1IPBrzMiaqj0S0i0/63tk+kk9oaxiEgIzNXIud0F6bdh3MJw9XnfcMHHTQP
HFmjK9dPFaGJNn+ozUz4Rodg8e4OWJ5yOHGPIUX5SkIjgDiVX9BKnPESrEjW3V7C
qrMVWlmszoEDCB73AHS12Ex8xtHfqtXNF99zvF06jSAfSldHmoMs8UgW7vVryEKH
8t46dGaHnSWoj4oc1dLtu+b2CtqkA9FMLp2nTsKzEN0hBIHJqMeUqQOYdbYE/nre
qzkb+x98R400YfMhXxnKF+3CYCEfqqZ/MJcEXh7/xoJIYUDtm3XSi1G9n9Zlb/Y8
pBXDyTAi0OYZNUCktdtwE31n6uPGXq/+pRaYXdbND5M7E9DfoZnpg0Bxc62cq7dy
f+LKWjPKwWquvIra5ZOrghfINWAoT2ofI+Z53enIpM6CCVW+YNUH2pUdzuVJTmON
zOTe+HCvi1E/YlUC+LQUmfqWUzTQ00+18Js4ntLrKmFw8HQ5Im1ooWyMi5J1C2Sz
IGriCUdF1TsBmu8iecZI3ccmXqggD0HwsvrtHT7++KEgaJpqgBYIqtQSSHmCZjxt
wcgFkncozMQ6ZWatIwwxm03hkf7cX1/hfbbNIUVAZ3+SjBdV0UEHUBdHyxWFenqX
lbI4qEOkCurqYy/GCL6R0cZ1vQFI3uyqlhWgayKfX0vIZtGIjG8lAJW/G/STn1MX
EplME3zo8t9fqm35eaJLINNllLpE/+pXmYE7vRWseNcRshmoJHX9eAJKTvzBMmMJ
f89QM0BZ0VuJbZgZcSOG7qfa6h7hGmnLSH2QmblRjTc/DSYYiy9AKKinRJ8LxYY8
2SnnnqLvBlVxZtPV9PU6SmNplqES/TVp2pvtdAxW0Ik58fwz9e3k2U3A/n1x+S+j
fH3NnBeBXHRrvHRA/OYhM8Gj5XH2SQAuYhV5ZQcd7QnpDOQHYXG8XsOv/mkyMhI9
hMKToL5nX9JgCd8xN4L3RVES28OKC4EOxeFOyJLRlrLtYVRcArsKcY6rarhOMKtz
4pEaScASottrEuC1P4bdwVtUSbiovG5D8YgrBI2YtwMsH1zJd3+7/dcp/wYGBwhS
6NjCRKZJjU5liICd8+6CFHw89aH1Ss+cxRF+Hepm0OLo6LG+VWJnJkx7ZqmeHiR5
3yTq8u5qs7eHo/V8vhLNLYx1cbxCjD2MUxzac95o1qdqDe/cNP+a4WCoT5/9zQlP
iArqO6WZMA+GtvcM8RewqGcCNIbNix5kMrSahq5tM3uTom9zuSTmnI89hhp9o+HA
sMh5JvhhTjp8C8K7evQXFHCSCyh9vHk3UGsg7uOG5AnM1evaYW8jPv9JOG0uCGCJ
aSmhT6C/z40zY2gpBu/KYfmzjoC77sgZeQvJpOhmg8hq/SC/V7gyCV4AdIoYxtvU
PhfmiLHWt2xBnuQYnVXu+WbtCB1lbgJpvwfxpLYNzIr8U7V5upEldgkprhOKvATi
ptPR4gOuxHzp59HTX00j8/1n9KvnIIwL8ElcLEdqoFbdgC8VgFYcSagrn3PS2Zvr
TazV5uqQgwQTjZegqMU/oXwOHmwD9UZkVeEowjQF4EYZkgLeIxKZay/7zaVkJbl1
FLWC4bbbDNrLw5hxARccqG9rMZcj6/3lqUD9o5qDTQVotCA9HiIKSqonARNGTATl
7pGXsCMEvIj6yiiFhrPfv5IniR1mS/qem06Z2P6HwDjiV69nJYEzyHK96j3841uC
WJni3zeEBzL0L0YN/XjJcVELASo12iNJiJ7us+v7K3ddAgPLyIEPbbpMF7HJccFS
GIflckCn/1wf0/P3AVI7zNUz6B7MAhPmR/hj/Vs+s9nTIdAm5G82B+7UrQYo+TWb
/ki+5f3IbiwOArx5URPN2jqm/ualCfA023/pG94FOGiKUBo6kwxMJo6lRkbLIl5x
SVIrFRNhH+RcbPK/YGeYUgTKLWQo6cCH9kdPE7u8thzA0Zxr6F2qssbOKhSkuPuj
dXuzKE6yNZybyp6F1VlXXzGdottcsJ9aPZwty6NswpTTUlEAL2/nNv8PB+m8voVr
Ml2NUGoH9gTDIJj5BOgyY8JlDwA+0yEoGUsTjoBP4sBNhp2j/GSl17+gV3OaEX3v
9PfKh/kTyqyf1FXBjdSoW8pUXPsbC6czfqearRhBM586Afg1eHGSdDHaPhuscDJg
G2Zpbzj06fekH/OZDMzgawjBlM9UpMBkofac3b9ci4jLMbdFBnSaLh1p1UspG+1D
5jFyUl9XGNkKHvKxoHRskRxSaVnJDNBPOKdkdPVHijuw+C0pN0ZETEy0FBeQGAv2
SaRQLqfQ9ILVsJBFSQHxQgiL18Wq1d+yQtTLmrsOB6PYK6mPRwYSaysLlfd92/dd
mB12c3L4jzo9q2zOgwdqjphO3QCQyV0eMLfmBiL5WgRQUPsOB3m41uCuGJCAUClA
vwd6/1U0jUC0ZvSdPhoMMbwHkYc1m8FqfIcnL7jVkEo3Jmub6Mfg3OrE9QINZz0n
CBFqkMpoX+TP5h+fI0xSoq2pnTYHU6N7XlNuT6IpGM9iY6bS74yStMiwEgxW+C7w
73LKjS2XxpP+CW+g5dR/SYF2JscL1aIhb1rRp6CGY/qzoFsX1+0m3utTDIP1Yv/e
AGHyr34BCTJX60MvaaTclKv2tEe9/Co2nraCzpF9OKz2NEfYI9HsO2UIZOhZhPdV
pnthKD+prnSVPy1bbQjdZOCxjW+ubNhzGytfitu4+o6QvdVBmFWrHIBfFwav3Pyj
lHQOvp3VEIZ2pKoWCJsAL4EkxsurvWYSudwI1taREkgzQu1kFsR6tE60zD4JXw9t
uBS29L9FCaSaaQMqMnnzXH/IKDP965mLYxzetdbGf7mujZS08E6TpjowoRpBibKu
iGPEQFJSq48A03MUJaLPhDtfwgfJMmfrGompfr1f358hK704j+11meaUX+hlLX1g
xbmjqiNz1711iB0yD+P2QA4bhv/GNPAZ8KEYBKeYHMxi3v4wBwcmygmp7GPIw66y
x8J6ZRP6YURfKbf5l/YBo+/rrML0gQFkRcR+3Msw1mn8tM7UIq6iAjobxFZBNOtS
2UUoEFYuxzPZi7CKBSlDQIpciNDmApxf5jCAiciAFqQg3pjUVxUL65xfe3VqvR2G
eaV3K4gyxmoKeQ0GkOcv4XAghCGghmWezFpo9y3kGt18AwiYNFWepqk0G+XksTJG
8+zsvZhm7wZyIdRQoTmrNlrIze5z8Sm1n5lalBLq+84avGsf39+A3cyRvjKRMCUd
uthJ6uZ65jBygCek4nzIfYDuN/gaf3eRagT0FaGV9p/97G/QQiy3Ba2t7l7grKRq
bEW2mKyzKI/pitf1oCp+PBF82evFj0j75pUTEitlk0vQlNjctFt6HWLPz2a8W+1z
inw8fJba0DqYPsT+h4msCFy3lxWDf7DbERem0/O+w2UtkX5qy+u9ety0wfzpPRXV
ZBXNP2LyExC8I7H1VskN+/FEJNQ832BObY6xbpDlHNVxWwMvZTPeMZj174waE7y5
0eRcOkkvr0zCRuFd4Df0yPCqWr7MnUPjWwh1vI51u0XCfFRvxSfNftJv3Vq04tS7
pdeZCMUp1Z8rtV4KEnBI2cmFJHogtm51B2oOEc/1ddyrK6mg7j/id/ZpVbWU6/eQ
0BuGsfMKkQFRqiN1YTRCXyHpNr7rHY1pq+OjnXEjsHOkqiJwb9vXGluYWzm2+g8h
obGYW/IHKr1LygOB4AXC/Jwil4aM93+QW7cNgj008BfaK2SxPDVxoDGXdpNnNutp
JH5uZsUIg2YxTNzrcQ1pv2Dcnsp6VDX4c1s8kMYWngGVjqOpP5LEt53oRYsPDaHV
2pfVPzfuSUE99NYtHVTPm3/kKIvkBhuIOGeF4uZn3YqgvNap6PfUlUUkA8MPBS+2
i0ydHUeXdXxH26M5Wpnj9AlXVYRGAtHapQb9g6rAuFLXmKQkZL5xj7UZCvhtX6oa
oa3LQ0X3n+CqnoW1F4q5ohGDNjEAKGEq69t3Ag3t8OUyScJCvtRUozaSByXNREWj
5VVFarYm3F6eTskuhP7endhozUWIInTYS67VgJFsY1aM4ylDAHng6UwRT/f1D/OM
KxXo0bex0hAaZt938GthXbSb2nGe1eszesvSMoFN9KNUPvDnCj6IfkMClBvQStUT
ATyfSiAvIWNd1EVe+XUeQv9b+Z1toFhT4Bvtq8K7fO0vCzARjDM/AB2lCiKgY/jf
bkdk3D/7+YlufQxIE56trXjkKjMsLCohZIiJU0uzXkgVO8kSCyrNzykGUKkUtGZU
Vsj5+z0wSSHVdEPnGUd6lSN3BvYkLzOBydyvrfgvzUzTBSw/wbwOQVg2xUzIl/kI
xJKacHmaejuDGg8mzGNRUT21Su+xYpEGEkW7bcEYtkgL4qsLrKA8W2hIgJgBpsaD
cUCe4o1abALTUAZ82JsjTuuZHf5KcmzoUyXxb3kv94lZMeF+6RdFScojT9tEAtHW
BdTofoTmZ6WPWE5XYP1/rfIEOe/SqKcSFH5FZRo7cmSjZE4EMeN75ZHNvuJl85Ha
rd7bm4TXfqDh0PWUv1vwjm4cVqE4LlZhJ+sMzbk7ELw/0iBQpJRpdb/Wcc0Xj7ZP
WT4bVEYef1rPhidqan/SNAznJiFtBqAANhrUV0yOGnrK4rBz3G9Z0FnFIXU3J+sy
eRkKZ2YU5BPv28z28yDoz442X31pAq4MaXquL6qLpfbQ3uiRfXC/ABjYsCUD8A/o
XWrTgM0f8Nu3mZYko+6etgS98oiKq6mt/c0voo2/U4K8fZsxrh8VlOiTaYPtgvI1
IxtzsB/C56/OmZk6FrmHkw8ykHfFErOojsxamDPXaakgfAI+RU1GA9YaWwWlx0G8
xOdrddRmMaXcVgvee9jvhhrSNniG6ZGyXaHYB52aMEwJttZcxskS78Q1RmWn3hBO
yekiMElKLGi6FWQkqJhQYlYg6YNJEZVxzUZK7ZmCh9zA9DaclLzZa1sDa7+30H0F
sD0/Tqse9se/hSYmh3Eulcvnefyrfp80mNQLs3lAF7MHuvjzW/oDmr4XO+j+yDHo
u9EE+JeCV1YaqBFsCQ8fdpN49hHk03OTI4ngD0PlF9Z7ngVhj/bjYK8LolYQziu6
NLW44KadMkhQtbTcYvvPDN4ctH3xnxgh54cQsDqXnzTzNQKhs4sQKkXoRPhd6/pA
vOxzIufFa5OJN7OXFO7e9MLCRbY7+Yf/XnWeqPMxAstEFcPXVIazNVeoHcIlINvi
Yee6ALsATCoU6YcmvkXrKfQfBe2Ptuyxv2bK5Mgjan5446hBaXomk9JA4Z19dwm6
n56tnIsjADYvDamTvfF7Js8dy6LPHdWfTO2M+L9srHakK3M0zRib9dL8ZBtB7eIg
ptUG3wfvSriTxLUiuyEdoQt47Qe3OudV9XXU+qLgV2wzwXHQEmyhgkjBV0iFEegy
48d6SLK5lYgjGxv2bQ3WQ+eAJ3SFhFoaQ60Jwt3D/+mB3KEgAAq528PcmpwtpfbN
cCShsI4ERKM5sVKM2cT7HP8PAvV9BOaFT+9k80Ua/58UDy7iPv+nc8hmCKE4cdxE
rMnwNeHcFwcBIkMicU07zWKC1Dp69eJjMZbCUxUgYCPG4mhRomD+yBHUO1r1gRXH
Ixm/bFpbNTdvNcTp7ODqyKQYCTmnS2Y8geTPqZXr2o9aVquDKlZ8c/vrSAr+QmuL
orXtJfQveUDp3f7xj5oM8WgkOMABfIFNOuqQIze1Pk1mEI3IBy3EE4RpQiD6P21p
kohZZsyxgxBe7boZNinXUOn0dafht1I5IAuWwmdNdBGIgAz4m1TboWddWfNoTw1T
W+J5+GjuO4h6/xT6+YIssDucnV5syHVNKJzp9C2HTM4IxkWzGLC65/zd1JmUQlgA
nKzjZTX6kLzLTqUhqI/Q91d0ECpwN1Kmrkjb3GR73IQPiR+3OC5PrG2BXL6SU0Hj
8eeRM+0uvis2SkgrnV3QEBhocIVr5phhW6Zm1K6zitpO3LWn48cqvPje7ZIe+3J9
MAs9x9oLF6uJM0R5dhRDyo4eFxb0PI6sm9H7Mmwc2qKFKDSXPTdmzBnq0IAbJlWw
U3rF8G3g6zRHWeHbwAG07SfYYfNwQBhpHuZ1yAssSpC3V9s4ndcJ93DVmBI31SYe
FQInr5He3dIzGyo41/GjKATs1z7JCSdH5/wYDMfbr03HOMVYm3GITu1D71ATQVKz
JRC26fjQDsU162YfyaSj3lBOXHIbP2xiM1K1aRc67tthGeWIbIIhyRVg55LOaJW4
Ur5xeBrWqDvthBnPCu2XsRvdDsecT8PUnMCg/dPUbLBjq3D8Rzdz0DiYckSA8vBz
PCtBxyoRgnc0Onh2V8c0oT6qQr/giwAy59OW60ECOXc3j7/nv7MRSh2gVUFT4AB5
G0XXZZ8xua0cP53cH9DeawLfd9Cm4arBY3Il8xfmsNKBWAY+3n+fbeue51yAD3XA
kRYdKmm8BeI2/EaXEDnraiYZE//Th0vbINPKx/eT1PcaiC2O/iVwaHo0XWsjBLPv
3VLQZmKNGYvqFNhwLvR8KtBNZskWFH+tsyCps4YPIAuDdN3u/jVwWWuYLzqp/AVl
BdKpRtE3mPCwwtHcmQJcAlYhldBSNKoWWFiU3nm2sueQUuuodu64oeo7b5nuXnl2
A9sHjjnHoD+lqw+ULgL0djSGK27epOmDkqwxAZDt0oTTgV36D5EiyODsfHee4H9X
wOJZPDX6uxTJkcEbfuVGqrctd447P5voALdrYVZmAcY6SfYLcW35PqeMkprkUzPc
4RfB1a////k7CMSbnANYQTv46/Xntbz8qIhc1R/w040ykfZJFnsZmFpP14yxt1Uq
60ox8/SR/fW/aUER5JDIxYOCnHQRO/YzbwFKkjFLajUyW93QNRzhSpad+QNnqlhu
9cv50FRFjODzEjPkAQGvMbKcDMMSJp4GcxO8OeiYj6LE+z482WpGq2aSolDRCaql
rurArksIr4PGxmySqssh3jexAfSdFNGD/HIVcnMxx7FGqgvtavonWN8K1F8bfnS7
7Eo0aK4MIP2k0+ikonnpkuV/4vLMxg4Az2eQt62aqvxG0wKdOD+VBmupz+FxNXCj
qgpNh6boQrZZJQmrRBosui0/2KHiKjmEQeEQXvUdEKgMAP1MvuY+XP3ysrltY4X2
+2jI4XMiAisBZXjtigFypnBG/7TILJQ3MUf3we5Dw6gAOJrrQIVgt6w45kR9Zox6
q5u80X6njrL74LlkvtAQA5ic0jnV2BFQx6O1UR7B0YCBssu7Nalkv9pMPk+xmrBb
yJrrMnenTiqM8jB/A4TtBBs9B3GEJXLFOBSRsMUDMIhDN4aomeXhqx589DCbTbcJ
ZcFpGiznpN2H+EMe6u39tRRCeqChCFes5MUk1ToqHVFBEjVPzZ1QwG16of18hDTq
u90kbfw7buVluadH8zyAktt9KZLDdPn7CsuLJLSrZ+ZkPC/0Ah8k9bXh/z4OMQmc
8QM6jAjfCOkQR+Wb1O8hrOckPUU7M7WYXlqSLD095cnjf4UGn06b76h1+usA94mb
T50XylgFNcDm6mGT3YBPgzBD+TQV6Avt6IPipKxKhuDL7f89A0EBdb8K5uJgrKOa
RJ++v0RiMEXcCwJ9gFAzX+UBWmPyLd/1EF00USnXALHvxVhEk/NCC49yrSP9HMpC
pv2gc6Xzh3Y+3QvrDCW9yLYmvgIUlSNobxqMqYnwLrFrfEzcjyoCwF9qy9huDLii
LAvjBAvzge/9E125aTsjHWSiKSVMe0E5MPIm1Ud26L6wEV7JPRY9tbc14cweSfYM
SJ2YVzZpZ27TD2Nv8Lwi3VqaRQ/RCPTO/r+Ot8NBpPuskg5zNrB+4jRmSc3BtbDl
9U1qF6VjVgvqYxap4RrRN9A5hCZZup6oamInn2i2y/tEE04jjZpUSXD55HNWDNM4
LedO7CK6eDRviIBuvinc+UBHCo/lrgDSJBv1gFwh+BbJg7GIAwG2l8T7o13Gp2cv
UgMmlEN1FTRhV6rqsOnfr2ORcJLRbeud82DZp8dFufRu8GmzB5URHvdGe43vcXGh
hqo9dXwC0B97f7GCbFb1IryXqixtLc0MGevMM40smyrTeYeiNFKLHbGcEiHXP0Lu
unEi9O46sJEHDLoIqCaxcEOErkjv0KQe7EEA0diztVa3lcJHca7PZDJ6boRvzy+E
NKH217Cz/rp9TUuwrQJEQMZ/PK6Dwahhhgr5jTHD8n5A7gcCWKwugpP0E1qGnbPv
SWz311apfs5xiTzUBuLOR1DCE2CEcnwaIBbdodsQZkCgXZKCWsPdFMykDWf/eSnL
WQZYpP+cWAVwgyq6LXvy5vEtNXdBcZUzDMCQ5LQ2mzsPoTBhx4ppSbEVmJ1Wyml8
p0qXPcDUqRdt76ne+mr5DlHPb1sM/uINeJ8LuJrcjA5caQvJ6bxSa2Q3gDU9GFyU
zTwhfS4ZpW/KnY1KRcYrPyRNkYrJjhXt7AGlihFfk5PRuohwSo1ZTLTkDgR8FWZd
fzssyWicOK668f8szzQBLxHkmHtKReESZcOx687adliYhTqTwV7TCX32oQl+7uKo
mT41Ao+dvSuxGf8Rp5Zl5n2YqVm/suuDWgA9sia+Ikiw1kPhhc/mFcZNW9fiU6Ir
LYbJHCymqGIBRCGOwPlyEiakZrCP2Yu64ydwlLoLkYjC3KnkvKRDa7K5e7IfbO9f
2O9i5UpBPz0cMnhO6rmjwNzGllOct0UFFG+yOl5sAyz2n0awrdZUWw0axaZzUiH+
VijKhgZrCQ2dx8kVENbXXJtA2oMF3rUlOJjcsGhavSsZQPlfvf3gKMRY4oB7FbdZ
6Y4u8yfuMQqwSy8D+cBh0Swioz0EvT8lb2D4wBgMiMzwLZsvYSNk0/ljfHjs0zks
k3NXR9/pCY+CqLKhxp4pjWojzkK63j1wWNfz5Mbp0T95tDw4nTf82Yom08RrOLT4
Er3qq4bUDqiM7gifrZsUFtB8e0QMbfqAb3yc6gcYZugi/CVJXvc+xGnk2Sts0FRX
qTqRapi4XixnQFPHYk3iy1TSPlflm3QOSeXvPG8PE/24mit7Ahh2Z6CUmrwBHjOY
2/JRos8a7if5mcRAwHn8fDGToG3QGjVKV6+ozcFiwKj//8+5tH1m8H6Sd68zgRwa
BKPvEI+bN1FfkHwnz0cjsH44k7GmchAx7/Ay9hQnHMXm2oOKz91dRr7CXAn3twz6
kiUGKbl+PXPPDautqj3T8Grvcl2aMHoALiHOGCwB/Myw85lPmSxEzqcj23q0gEZE
V1xur0Fj94e9i8PXpv3weKSGs/eLoaL8qSfy/xl2xG+gLAvrtudYyxxrX8tCPFaH
7twJbxniRKlkFDsK1ordHzUMJphBDOnvYWOiushNZNPu/VA1EDeLsVzByeRWb9EQ
v/o69/WWUYmNzZGjDSMHOiKQFVvx5fSABlT7/GRVpIzF4Z9y94sStiBXVV/qRF4j
FqfYDR8MOOYe9b7dVeeml/Nu2BOrl8QBJMBkuBQtR/9s2kP62FgHFRbc7VfOdovr
oNAdH/eNollf85pH0b60XeRSyYm3wAYh++1cN9CPWxPdvuaGHJ3wtDInGVj/DN5G
BBo9+1Gp0imF3+uJROl56e0KKPBb3v4wDKZpbxciUCkwYMdiD6p8AdxLQW3GJyaX
XDKA6nnS/7YMH1dXMKkuE6SELBrg6G95ZuhH13umzmEHAVrnGIyx5Cv16+Ao5bm2
/MtjnMTyhsE+TA8doLnKCXMydWanWHGEO0Ia1EBmdGi/QtkGDvJUWCIJAMZ+8A30
J0rFbDgxWolugP8M9IAhSGEi+q3q0dqwQTB0yIxIb+PDFxzQjxGX6uhRXkf/8flL
Du/GM+zYUAhD+6QkMfYceAkKwVwj09RCeyZSz5crwzs7M0M7vVl6Zv8b1iBazlal
23jT3Ei/1+B9Fg8MF5Do/zryGyawnfHO+yaIlhiADjEDEht0MNd9PvW9Ixmvy4Uv
RwipCOjz1pf+WTxhlnpjaDxQjsfLd1ONGoW+jOxW6a6xjxafL3j89Hywb2f4Qm7f
qMbvNwMjV3eoc/hP1GXN23BwOSphX4PLEYnFnhoJS18t/mQvpuhwccC2Z37iaNNA
MePXKuBVy18ByA+3NAKtr43iRza/PgDIJyfdCG34PuH6GoMftaIdX1nu7dHiNCNT
X54Wy9OGOnUdAlRWHetNs8Ugv6Aj0sOo1w/p2ZpsxwB6AUr1mzkN3GT/Gp/C96w+
0a0E6WNRdT4lJwcz4gEVxZD2z0wnjFRLk1+bSIbSRgVXxtPWtYZIrUOaSOM5YBrx
+O37J/zPEENcx6FW25mhlyHj85ECHfR/JDTFJBhmlYJ7A0T5IF1NvI0mnPgdyf5N
sy+Hs1Sq5w7zzfzouw1/ZjWyKEhHWGT51OwcZ05xJEiArG2qmcJ6h8TjNvMpYPFI
TAxPjIhZBuVER0S1TNg2dik/2TXR2QV2U3MhCgmxUIdFBTUGuepOHQm8NdWaTxpV
TKiSasNL4eM1vyTLQnR7dX/KEYl8jDEy/DmnjvOcn0YPUH1HnmG9bss9mvyXYbYH
1+xzMlj4RpeHwVofQeQAtYGwVSRSGZLjLuBORXPByKhMfMdExpOrDBX1jCmTRUEF
x4RqkNvvFBMpNrEz634TjC2Kt0mJb11hrPf/opnch8tEy5l2Av0QzNul+o+tcfAX
LpfpOiyidKutHI3RSI365lI8mFqD1RscVivTkKBIDV9nT8wFdZLLSHuJvnhmk2Nc
`protect end_protected