`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 50416 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/9huKRhRMtvnNqb3Z+UU7TahEoHV+T8U3P3ufru7l1O
3DlgtZzb9QxCbOjthp9+wDkjygH0eUfDrEl1ovhZG61qMVaGOv0dpUNw1ENtMfBW
aszjOfaFjp6xvAa9LghAqKWo9GaW/axHgQ8SWy+v38SiRvUcG+JyYGtp2Y4ZPa72
8BBs+tsXUrRSrqSZxn36yKBvkqwwNm5/y3lwE9Zrm8QVdcvmjEGdL8eJAVB+tkWa
5apm+nWoodvvUw05lZQ3i6n/uF/bXY2CMcwvuU5evmJs9yO7rsds9YVVtfcKaQMr
PvJb05+VqiJDjQYWNW6wX9ZeFNLl0e++VqtoQ5CUshzGQo/6QVlY29xQv6vrg+4a
sGOPX2neonAuBY3EKWMtSFJwA3AiWJcKwTWXb/h2JM1cCqAerYcpGfrg5KYkOieE
gNrILfOkXOZDyrXllp+G2DIxaZ5bGwyGXU+nyqtDK0YpP/P+Y1lXrG58EIMXiqRU
VAc6FJEiVIOBUFXTXeDE/otbqBsqX0+uRdCyvcx4xTW0ThWPpLeohNg60+sXD7wh
xTuVK32afzDqb3jD1NZPNBtA3u4xZLlKeRe9pxHnrOj/xxH3Ob6+mG4SK/SvkTlg
XFt+ieIeuzDG5BgbIkDwiYk56Hlpg5r2ghkfU1+ejSOB72r8+p0V7Je443wff+s5
pZmL7woBgO9fO2UvbMzYsMM5aiq0tEaqa+MR++KHDcLCsGbZUgOqBikd2Iq9y7lH
57mnk9LPNZCdQZr0WzZjXc7Szv5tQ7nOVpkj6ov4Lma6agQgfO/Pwy4EmuQDMKA+
P3nf+51DvF3LXg/mPa2+i+wBiL8d0h66wuj9Mlq5EmFWFPKM+XKse0kwMQxo1uLR
HhA4RP03Pm5KMTnQohw0aZdiOjU26H7FB/vlhTGSCKZfiYr9PKFs7XqfaUrKFO4G
5iLgCAC8bOiuTPmHqxT4/j13SBnMRQTWNYWoGGUrLPgYXkdwmPlofwpiGhO2Y0kE
8j9SqyvNNV3GHCDxWXeJTbBwnKelyb8ftcvtIjGJ3v8VksTuEXqoglu0+xippQoF
YD16DQ0MVVtspuFJKN7jgyIAZvE6NNDU3lIj3/eqpBPXuH0Yq1HqBEUOrsvDfmye
49wapSvai5hLmq28zSgx+r3jA1sJ0kd6CCKB30Kn9HxCiBnkWtAopudtEZIzYT6v
5TiMR54eoOpJ+yn8xoqTBGOaJ5cL5q3e0VZd+S+T7JFLS1lmea8JQz/1nn8oh8dg
WTDGtUHWBJOQyzMwcnWdMDiKx2L7oXnTbSPUhepFMKVamj/symMS18pK2GOouzV9
TboWyqY/Fp02FU9U6wH+EV2B8lryyQ1VMHlEk+Qrhb62kaSvaqLF1lRzl/ESIBka
MQP6nMA1HmLipgoLsBRBQAEAWoqAz8atfAAiVT7Rh3iFGNdTcJWCNTsTsxzgpKDa
ccpKs+NIazKh/gIb3JIeqcnYKXHFx55Ur1oiFcg3LbYyWHVgKYPRW2DVuDhfVy1I
oqRazPb01eVSKVfpaOQYBEYc1BFYP0mNK8X8TNVpS8CGo/YjotoHRRb/yGk51TkQ
6hhX/dVSlwRoghPHxk9r9GxqfnwSnLLSsa2MZWfBAIwywiAeeFJZ5oTd7zGzwNSf
znax1wekPeFhyAYYzRU2wcEVbTn1f9KEstuRfDmklXShCjbAF3b2WT29XNC3C1yR
5m1u0Mvtb6t5cmzkeAQ2mirsUE1EGbVI6qRhyB77S0ITnWEbhGon+7jQuj5U4KF4
SDOrmnclQteWKIcuFs9zFWjeBQtXP9Tjb3ghF/roiFk1/tuL4ZHqNM4Q1oU0TOUK
FqgYUay+i0WW8D+0k+by8A/uOUT9chq1+6fKDfKuGHzOxnAb23XRKHY9AuOlzgpg
2WuPFF0I4rouNeoXztuZslgso85qsYhdRprrl2Ut4mt7sGKBM91P5VNVF9G3UWSi
LSjTbXTXeYI+UGFuBnFbEEU2nYgtWtx2ekjdqDQu1jLq19sD20kGBFek8efjK9tC
xf/iR5pvnXkTpP+Uw/bNaqCESEF+DLczT6oATgzWNE8aFsVhsb0DXKAPcJNuPajG
koIAEr5VwqLILvrwCSRiUKXE0440PTUhz0BnB8sfT4+WCDRxrBiQwWeVmX0dyNHy
UIE2QoGuCejTwmb1yMOmfcjNR5iyuDnbwAP0bZDjLQYNT1D2OVtVTA83vtn6wmtd
jSy1R65t+Uv6UA4f+qmxlEQs5KNFALCGrdZxlPUY9YM20i+mkgLlTW8nT2Wf2xmW
oZnCzemC2jre1PAS7npQ8xrkWH2hOmbX1PxvRCK9lVFDT/rKD2GOYVoK+rXZjCjy
CtEaVvueVnIqQ0UGm+8cApOt9FBsrrQmE9x5+/OHNpyFMxzilEGtP6S2DJTXiQHo
6v3/bZoZRSjDtKhPMDy8M0kMMBD1x+WnfYU9A9cSoH7lvwYHU30Pz/0IM3VH3AFR
i7y+H7WksUBJaUZ7Zsherv4ADLnoaug601q2hS7serVyVmXilqKceeHYqVp2AptK
0dhvLbesP47l2vCl8GTWFBobfhwUuBKg6isQc9uw0yFP/eVzPX8c7Y0ylS7Hgywa
kwpfTIHAwCPPJsSAs8J+JZRn4ioks1Ou2oFZVXtXCSFPcQo3x2ooxXEMUFMLQoPw
3S2arNSXkEcFxbKsAwT604OgRY06z7EIVJWVcx9lRvVASpz8H8KFqsT1m7wKCTX7
qL6W0lJLf0kj500OmPrXp0pC53aw0rOMWpKJGOi6d6reHxGmJBtwhcZUSmU27zyb
UU+0AnIIZj02Zt3lGRVQfX+fEebzV/cRSyHavmVjZfz0ocgCMX1vNyAOkxr5G85d
CbPZDC+w9S/6V5FowkAFG3j3wey0VHrDGNJzcm86Z5dg/q/iZDCsz68lwhJZ8T6/
Q1FsGDCIWbzHl5kqP1yDECmnH3iwreGCCU5OrI6NyVv0nQaAAoAhezLMky5lEl45
J6CTRZtDuA5Nr0CMLhJIAai35oSymnm76uNHrCZ/rAk19m64SPimMXBYLCH+O/Ol
0FdqgVeCgIQPILpOw/j81sNZ5xFM9AC/iT9HlF+J+D0o9guJjsSzrBNwwi6vro7R
TUV6i+3fZzyGNBTNkR7EUxU9qmy/6Rpw1VQHg/wesJzlUpisHTpPTizIO/5yWE+5
CdrgNSQDl2AIOmbhwf/Z92CoDC0qyFSSmaS8oJvObOrcqky3yH0XrxY0VBEoLu6v
2pD7axwLB8EBu3MAu1LbEty0qlrs2VW5yShcYlFfdRTXfizEZMj96Pkpm1YicWPw
flnZ7kLLTfkA4jsv4NU0CZSkHWNIl0ETfjmbnUPsjc6y8VYQryW2KnSeT9QjS8yX
5x/YIHEXUCqXGBGkgWwcedknqHMGpvp+jXcpKnumG/rcCcPwfM1panA0LYyPTjNz
Kff/+pCiCNjNa1zkit+BpmPCfbZODOczhNBwxrwjKqC8sV8x0eMu4aBD5DaVHAHT
wAe5QR2+P2lCpmsIs2BYje7lWezTyvNYZ/Fcblu2byYXj+KOLVK6RLJKeYF9KItq
HAdr0O0zeQFH7+lQwg4c4pYh1IDwA0Vnz4rD+qU5w63jHzdVwX8M5JgAFwiExpOE
ZvrvI7sEO+jpTTDy7vUh6PNENcYVTHIuCm3YCxN/xAu21V4ZVYeKIfrZ1hhnpWEY
iL3WfDoBrOjrc7xmkP6agEfewk77lowFxWKPafDoCKGMZX0cqkVT/T9VkjJ/Mbd4
Ogi8m4aRkABDMWXKgnqZfnzFJ/DX7cpaCD80/P+5UEpq/m4xn68I2uKxHryL3xOS
hsPEgAWVBqj3caNXmnfwzKBjSczeF1MdtOWMuIIa5kvVjsRWlJtsCSEC8ihsBWBt
ssXbX87rn95kOUhpdPW7EwbvZwCf4LXd4fsZpgPJNERev/kpeNR31dZSaIvWLftC
4EZxd2g2KBlUzmvMuWCrzNVtU5KNBWVrpsHtRNPml69mfGAiWWCsnyCVjK1g63+N
HgqkF2jpkvbVM//RlMeeRP/G8S7Idpi1X9A62SlFA+wfcLp5E5Hdh8SXTXWatFaN
917BMhYilbYuLKafe4YXWHPas16OkcmA4EDuG2kfAmRZPEB4TBRRCL/5Fb7oN2/t
EV5+oRmKa2+iTZ9MGqpKIVIQqm2OtU5JOR6gS8vftpAGd6QkxnEEQ2L7XvZIPICC
sKEX8UCfrypHZv+5bCvb4Edp9HjKgh84aa3J6UTc8qNe6Ic1CcT53u3H23gMVsXm
GTUvSKwETbD9byjBMiHTIOEfOgemBk7xKlEhTi7Mzhya9NH9MmFwr+btgrYu4Vk5
ujkt3Hg6Ofo4/FTIzgJn193hDurArOHC7ToC+0EZoB76Y7pD5TZlWj7plX/KuG0P
W2Jfgg7nIm6Kkmt5SWCcmmMTgUC2BKwAg9ARWIl8VGDOY8PZ3/2BQoeZSBEALv1Y
5fNq+B/1BtOKq3pXMMz9dHYJvdLnj7uZBlPLt88le0em8VyAV0HO8vj0aGhCf7Nh
j3yrkkGJ6kUx7zsWPSIR8zgyeiE4Bgnm+pRIuip85ZHJRma4ZpcxY6PA1qEQ1/3Q
u3FIm7cRfnZq8tv1VF/g6JBMLunJIDPuyW2eAITTieomhNnZwejK7Yyd53FwKl0Q
i/IB/gtSdQ4li9rgVUkNSV2MOvaSbe9KKjysEkYZQAL8q0UASoQu3ICaGApGDkBK
lVQI0/dUWvZItewpUboTav2D40SKK1qmJUbpzNhY5voNvt5HmarGwy75LThSSYd2
5bAj4eLIPSDeJZjjX5bwHHDv/Uh0QxlQOmYyr+pq92fzNBOD7PRWudxoh0rGt/iB
4tWG9sSib7NmaavMaTJ2E5HNeSdLd8Z+IgGlBk5sdSMMUQoIoBaUZ6rfH9bsLueh
LQbYv/oWEHmGxBfaGGy1InwsmnANC+SSOy3zqNUdFD5463dJEPnWyoVao6QZdrOv
NHTDDHoritdnSiZ2cYAJKMVj2t9O7Ye4Agh991CtkvfwTLUOc2yNlmpPXFPQu2P4
EwXRdtO5kiUqCjJD1WX4FZ9b1MwM+ow5mmlZ2ZUxlIcvzfe48EP/FuQqz4qq+eS0
dBnzqn+ZGBPpDIhdgMKnGHR303hDJ2Est5DCBQlzafT5P3hUs4NqZ+wn6j6avKyL
NLaVMg+/DbAhqURKQoPqucEgtj4amahOlogOqUHJOzuKD3ecJL/O5Rfv3mLfyYjS
qufH+o5AyfNvW20svybyZgTgYWayxBvtNF3hgat0PSzAF9o3rcQYzUtVHAfVcn6O
EHq3Ci0j74BFo3nTgkgU6HpNTRXb3uw6gkeBFwx2WTPDOa9v6qUbqp102vFtSqHQ
RwqtESDfcZM5dIyoJx/eOF0uSf4gaYZScyUMHPrS1Lig/v7bp+5vAtwFqBD6ibNz
Yl7Kfr7wqDAMCne/dm0gLJCv1qK7manp+U0q2px2A7R1H7hlF02Abr4HCOLNS+1L
Uxa1JIw/taCEebB9vmaUOZx7FTgpEEiQkPVHK40Wd5lBwikPUn5pTQpGBTUDnoiJ
tsX0RasJyCUNw4CcUPN0i9XCMc2yMfa9H5v2u0ThA/QRO8J2hYq6jGtq5ch0sm72
rtpv6GAoTnMvzSoq9gbPxmeyMzXhxhp7BGI3AfMiQolanremjEKbyWEEikYc9JZl
G/rUSzcLG1udPMd6fzE0WANheDK8Y3MJh48AMKiS3hFqD5lKrcXYIG3xvHi4haXp
61xCKIfW+FNycenhah7DK2ahQ4nyDYgjk69mBVtNDMpzkXeenU4cg6BTrz5UByWi
oG+d2oayViaLDoPOxathg5zQ7Eq6lP3uldF9pwy3UZfrH1FxGG1xqDd1UbZrk6J0
N7HF3J0IBHhAn3O9S6fLj8VCEx1vmFbRCN/X+2vsNSAeld7OnLB9p00Iz18XMoy7
i4Nmu3G59pvhT2mua5WCOvNpmsYyCqe3b33HRaFqb/BTEPPtdClgHdMkuU3OI8oX
ZynNeYoDPnCHp6s/PfvN8YNTpPAkjh/2DfN+L152BFDb7Rjlihe5n9LIDlEl4Xqd
6C+r/dMNw5PhskDpXSETfofqI7FSKr3utTrI+VQaLeS1YfGB+W8Kpq8/pQzAkNod
FXolQThUP8AkRGeCr9KtXxQ9v6jVu6ovQGn6Gql2vPaqX318mLUAo3Yp2kijrU/t
JwkKf453aa5+4OEN/FHlzNpIsjWCqJMQoQAQlJCjDYQZKL28eyMjMlAM5LzgQU+a
9D69Uol8PenF1WGlqKy9zqDxYXAibkjcv5l/OTteu3GfMUdTHd2SMw9k6UjHMSIl
5Cn0JOp8zQETNdqCf6I1tDttJsIDxPehg1ovjr+1FVSj4eNalNR0yZRi3+u09DBb
r+5xU5sQiUH3YoH09YGd4ihhVEMcVReYWtawa8/AzevLMEEgb+4lil+ZkfYXhtoP
S6Gu4C2QctROI4Ov7qYEOT9N0VmA8fn3TTLYL6Ih234fjQX+/IaeeNwsLuo2Cmhz
Iy7Cld2zAbMlA5l2d1nG0Yj8yd1eFQfjrx0ukUw7Sx/qU13SEdKCjO04ExwifJkc
hSlHyudB7v7bWWTtvuH0CYQZ8pP3md/wF0me9Yyh6Y3lXoRFWG4MnuAJH+R1/80p
EEwLeVzKC1h5tWOl0QvZMtcOv/Mzb2NtP0KPjT7RRPjkYW5DUfkiMPY2TVu+6YiA
AkRAjsrO2ZZzx5tsaDLlhthUkGbsJ76e4cSY0sgoG5R3CzEVBWXvEro0+IaqGrKU
o2Yh9OvA+2yrGirU6bCVFQCyxtBc4rU7VTfTrRK/Jrimy0NJTwUh7bu8OJXWXN6A
XAN0O5NCvF01grLpk48aq9LQrxk/OWLx9+5QmLJdvdt2TXr9zn22D/f7YEWMLxVw
ynsEOyig22ORRxIrepQuk1v53C/J9DdCdX5VYWNVjbSUDy5T2d0P6uIgR2QT81lL
+6know54pNnSsfm5QozNo0TzWcw0AstC92J7sYFHs0jhuQAxkwI6koyCuzUBkjXg
OxIzxaoftq3eXQfPsGRu0Hwmoa3qxDYYWkIBQK3niqNAJE2Vccqhp30HFkwzorXs
RabvaPMdxU2Hn6XpHlwCAOo+/6NvrAgyS7Ff2X70uj6QC1Ll+e85oeHqE50vxGq2
gg5spZWFupRnmrrJlmM2ZCJQu/WV/sAtg6aKtYwFfMZlbyZZmX2CnlUjwQCC6oSo
B2hBZUDUIhON73CJFMidn1mW/hPFmcXuXnfO8ynVktOiF8NwVIyWAtq3HgUgmfSZ
DCzVzwV2v7xtE4QEbl1VlDWGmv3wrjTa5+Oozd+toiTmi0u6KriiJ1oCAdAPaWNw
8p1QrWJeso0dwndasR9pWpbPGZCSG27qZQ7xGANTMGU2Cn8+awMmDNGz2hvV2Teq
/GMKHaWvpA1UhxR+8m6VfaUasuJa9NG8jvPl/4tXA6kIGxuEKDJSCKnBJpHT5siX
Kil59v1k6mUtmFKKnZ2+v5QyoYGx5E+RdvJeuKsPSnkeCvz3I38hhghWtSIz2xR0
x0JaYq+7LV42ppd6YZnWVtsC1xXQpkDPP3t9rUvj9MILWiCiv888k2U8mu6k7wtr
S6NRgJBCax7euDW3mQKD+Wzt9x3a3cBIq0tpm7Vl7ECkG8BwzzJBBHtexgVaCLQ9
WnqSAuZrs7OI8b3XdEugpApEPLq5yVepCnh7tEDPvszSfQEh1Gi074/yH1sQpugy
8zNlhb6IltSyHUtHga+R7WWiTfufTB9EKw/hfJV2/WRr32v8fDkSIJIZyt+nSZs1
cQxozyloazdUaBYtC751SOKUOCXOLlh1ne/WwbhyhZHIt5zd0woQwea8pUoszVbk
MI3BxysGrGvatCbcxy3b2/RoYh0ENMLWRXV9E5JDQOEyPrXeeqwRvLvQ6WAOu3zk
tNh5LKpyL7MYEiFLOUJupX1i28/8nVqVUadumeCzU1aoNA+f7PMfhdhD7B1xuN8S
Fx2D9HctUvdqF36KOnTuaeZHU27t+niu8b0zRUt1UHkb3WJ7PvQJYbj4I+ViVaEL
ISY25ISfzC2e9erP7OYZe4t3seEaxAdnS+g70Ncfzvmt9mmFBHvuunUPY1KsSJRt
Hc8TpTHgT5ycnZJeK/Lqi4nYFpN3wYmKu0WM4qmWrUilz25s7Wj8/ZoGM/PWhzDo
lrx/KYeJJVSXrZu2qY9Si5yBgxzYaAbxg7FKgJESw4Aw4D9sTf3Bs0WyRN8LWEdz
ahnbynA0jJZ5iEpEw5FkdEcOyR1+yFnnf+bMR9LYA/zHYDZDgt3/cffFp8k/e//i
b/RhUPCQjI7AlcqAP2vWPL8mRm9RWGFDhzA3h09dj7P2PzQAQTsjdnqUwIhwF8j7
YczzSd1G8HtHRRUT83s1u6/ovD065kbrBNJiY1E667/ismITFR2l49IWVF/svWrv
wf9wfgOdP8zj2AWeETpTf+5g+A/dFvusTQxdFz4/ET1b+G1B6iXedDbDEkFJWS/h
LNWbmzq5c0WCL+tsqIzuJJ2uJXYJZqFsy7UejxegLAUqO2iZVJ5Rg34E0YyAPu5Q
IRDIc2peLIvg+nlReFm1O8Dg1divkfb9iXcX073/1cuRm4L1p6y6/uexFf1cYIs8
ZEMLV06EeVTjf5veA22peOFjer8PXZ+a+TFdRYC5Ujzz2cI/9C9T4Wbfgo7V8Y/D
644mUkpreViAFF0ezaJ9UMR5D3lQxRyyAkea3eD+xOTSJZUIRobqRChnS4bymXPi
uOZIKID+AUirnPkAKycevyovqVHUVFlEaa+JrNrtlsMZDn+2BB9R8WgS1gRQXxfH
NZB8BHgI5AY0F+cZ204ULrC0ik5blKsbwuIOdvGU88vldrVv0zAQG5sVhaEfSkqu
43q07OQgx3h/hFqn15b8PRTsUeISUYYH5hDkm7zf0dbXKHB7jpzyFM39BVNDndTh
7xXg9PI1HcuUJI5UIZI1/o0rl/74CXJip13B9D413aDO+ACb15mKKL9kL+vQToT/
EDaOrUoY0w5xbMoIVJWJ1yu5OLlsUBV8E3bObDMKfmphhlmDtBWQ4t1VTyAkcFMn
Cyx0Fl/ijKirghriMJOgvQhZ463UY9ovXSzciEhCewAQc04MHeuKmp/owlwlmSBC
3XcBO5SExgLCQqdw0QU/7uzDmWnOoLwDhm8YHclhrAsYG0wF9HKQvydGO8NOJ/bY
rFb2mLmEm2JSmrQGXy6lZB2NRhAHhS0jT6KF7gUNCPHzp5w1mhREQNZx9x/fmwnw
q0NVt9Q8NufaV1Eloijk/vNFVszmV0dRx5aFKK6EmiQRYSOdlWDxoHEROB+uBtZh
yUQsd+gUEIVrzCPJlLpJ98ueY5HAEJiFaA/6dm2YWD5KtTHM3akRZttlTOYjd6YR
bzdYooEEC/iMngspBQS8Btd7QK2JtY6IcMg4UCB4zjRIODJCI070+oYxpWB2nMkr
bcOANWQInj04k9FQ+NUBzkmThUVV8Tg1TYioOmIO88omRTfMEa5Cf8h6e2278KAZ
qYgGwPEWXAmOEW/KQk1w1GtkasGYqzZku74I5HQboFBA+WAJB7L8B00wGPJixWoe
MtRy711suuaXepcGWfrvRg9SeqFD7Kk1DL8QyzSPZn87SpXg/mzUKiNpDKDBOZid
dMDgsQypkGGtNtBloO9c7zcrHb9YE3zfgx+YQAPRdJbObrF7bc9m8fKQA1XxBr97
bqMCqm6270GJ41p8zbLZ+5HsDtVK+P2eqtvS6gG8K9xk5G/8rpcUMIG8aml+pEpE
0Va/vbluQCRI1G+5HN3pOIoJsYqBoEv/VZkFHxv0vh7n3bJ7X3HHs7J3DOOlcEgM
dP9E6LbB/qcthsaaIzEoA9ksARkmjOwuQa5EV9+QEhAxbsAcDMwVBs2Aq/Drlf/k
jMGb00LeLSfkxl7avI3g/Cr4iI4OnFeZxsdZ1H3F+e0o3L54hZZBpoctdfjJX3Ql
/80HNYtnkvUESP0YpVz0Czlx7djfs5lDl2rjGLbE1nInU3ea4qeGm+/IFoiZz9oX
FnO6O+0BKyDx7Tg7ycP422fkiCQ7TzbLkbukmt7SrPlyIjG8MBFOMHBN+vWmojWb
XGVA6Tfz35jKpW6CK1EDExSkngRMBOZqL3EqPIeHRDof91Tdn/ueTUIm3xwnv2AF
zMT10hxYzXm6Z+nSoJn0L2OFOSFACPjMEZMxp62Cn3p8VyDe8viObv3L36PQxX8B
zS+2FDb161hBEc/6xlkimPkNKrai56E43TKccpWvnyrtRojass6+r/h3bZUwEKLl
/45K1TyHv8l1XshKot1virxVUZGYtKvcDMJ6D3kBoO2ypa7rrVHRI4Bru5SnxrUR
3H90B7HzssIYiR8rURZ7PqP4iiX/wroC9vSbEf3cfjB9nDnS2UJhJKwkmZxZysw0
JKzntOQzkEbbWGAGyAHoz+4oHqW/rMqNbyPzFy1FKAmiaQGAqWtfvo/ArfrSUezx
QGhfdYYaBNdJzaSJ/BUoInbaU2tvXArq6fgJQEcK1ijeyf70xpm9SSeW9hCkHS+H
q5LcDRD6OmjDe9B88L6L6fVRb43BeiZK02OoQXo1M69+NuHsqeg/wNejCamJrx7j
Rx2HZaBQm4hEj5HMo/xOuByGrXJPSubH/jcjxHlXRyrLGlRZ+UdZlvjF1Nk5Ng/C
FRHacR5T3TvSJX5RMLLuOTQgP0syYTyrrtl0vb2d65edPt490OZxxrIEvsQpdKWQ
2q0ByobAo1j9I6mxVV0ax+cHxaf1WrMet3sI/uU3sDOHq5mh5ROZvDPP0RK7VoKg
b4DI6bN0SO13/TH+f7wGZIaEcUJxbAZDn9csZfLSlNdavsfAdjBP4uGH2AyhuW52
9O4/7QgDnSStI5f5Y97++DcA0KD/oXN2nTCiTU9QDX6AIQwQYhd7VZaVM/tgQrrP
wsSn/3qLRcdn4KkmM0/132bOIyGGuVn019B4BbMjTJGSVXOU3eRRQXYuUnlwviXB
z4I/gIz6qigw4GpSw9kj43oRBTSiU7I4r1KnHDIMVHctnwFoO9cEhNXULZI0i4An
MtJsFm1E2w9BTzx8wyHxkBVSkmlvUgoaLchoOXm/N2kLJhYTvsHIVc+Jhc7r6ga0
MQnobtqBqcOz1C+dnG6+2IFYbrcr0ZjMrXXEBMpIJ1elpmoRd/HEjiCz2/PaRHk3
qrSZMLOrJ7akRQV3hnNzDEta/bOkj3KaseBh5IeE7ZBgyxa7K361fBRk7jed22eX
RxLJlnEV7AFF0LrR4pr6zNwIxZGQSDEyPb1uXnGgCQqm3XPOtoDYd+PctwTbn3bG
CHTG9PCYDw5DTMQdGUBcUFrxAAX30xNoC18g8QZru5YOXElzAozo0qGSqsWyTTb+
aGjYOhyVS+GRSUHfz/r/tVKVS1vbSa2YtuWrFFH+5vZOdXB6jwLaG7Gq7nM3m8Pe
A6W4EvBlOIMlsK+1EgFSoAinS5otF1XJnbdzs2DLqVjvvrKogASisVReaOCqL6QI
iy/C5Sz7JhroBMXaIJEmS3dALJol8F2RBnWYb1qt4FAAJIkNCsemR5zZ8iosczqK
xKD7JrQ2g/sIdFAQ4IxzkdGc5GRz4X+w5S6P7/CNudWRKky9jyCg0VcOfB9KpQg5
JGbdyj/6grPUjCL5wn5j85CXUT1ZppBaWny676skCt0oUGtnLplafnT5b1Ntl6hL
aTFVXHg6SsiSAlfqh5AvYIvrQhh9uXdllBPMJyRrL6h4kKdr2GLQi50vPpk4eyqv
KDEf5I05VUcFSVe5Ix3SNeYTqbGks7UtH9SDLltAU2YQJVLRHYCrcT0eSkHQJjqr
rNaoB0kk0s2xAPlVatVBolzmdyizIQDte49KMay42mRO1OoBn4wtpNSonUN499gy
1GeJhA+CG7WTh5VxnfkwX7IOgdJ79dZvrHh3Gp6pNeTdqKibL7juFKchp358JxT9
zrwPe8JFpG0EmvVLaZLZewk/veJUkA3hY/Vpil8pPs6tRlfRw80TsO+8aDrX5WI1
0Gi6vqiOcQMEGNKgcfFyiEyELM7glWpoxwGHILc+xC4neUJL9tRb4uVTVzQcCOED
8I/EZNGo5k1k3BGARN5bdwEF6YPmInpNZIomQjbZgZmbUn5QZI9XthyIudbfnVs1
wLgVn5XtB6nNOLFJf0BKXisDf4eW4h/3aXhfKE3mwJqamqKZLKJMp+/xKN3d/Udf
gFq665+GBIrvVTWTgmT3owt4BY2qYmzTAz93fPptSHaY7qa/sjforVFoSBladqjU
/By4drzl1UavqZSIre10SvGF5K9IqYDKKe+dlPUPHkFdABVnl0n0q5dmdFENEFqg
hzEP7DQoe7JXNSkyXvVljZHQsXMrzCKRZ+bVh+Hf1tndndRHCi/lLjsJ+ltxKP8q
89naBLPB+wW1GmUurhjRKARtUFlz6rLYnNMPYcJKtx/Ly35WtneaGZfcFYHCBnsi
xaW+8aMYIhltTrI1+PO9Lu/6K8oJRSMQ6VyqHddRGdF52CzvqEIxtUX9xKawsz4i
VbehL+ceAhQweD5t9hHiiErjfW7dbvaYsAk5AtpAtH3DUtqN4soz1sC0jIN2/+Gx
Bqo9QLcSlxnhFALjbRMSZIWaRwq+Yv1NMXX5lgx8NZAc2GAKZsYe5rTSdTqj9/5J
yN/+UyMJ7vVK7RaA1XoHyz9CZbQT6HrlaXD0e8MOfhUl07o+KawG7JLiYDnYJTn0
AIFdnC20WGYx9bN6CRlTXwnm4lh1Kr98iqlK9QjbLNNq+++tpcTbOfRF/9u2U9Aq
HnehmmnvNLPg3XIx8f7g6jYCYka5JD7JuygalE/A/t3lyiyCXhHburMgowgIhcrl
86rFcJpKtcU8R+UcYkovXyKd3xOBSPr554adh0qXpjGl7biXN6NWDRa8m5MPcX3y
mphkBIw1nNg3i04PO58dUiK5rSjQhOjd2P0MIGfFWbUaeDwXBSzF6px0I+B8/tWY
Khece6Aeo80XRlRG754OLIRkQWjyYOd2fD60NNJTcy6o2lWXP3JSsv9I6RPoa4gC
qe6oOPn9aUomEKnozpyxSKqIDb3ssqZ+WD09BLH+EQ+Veo7APmP5axC37JsfJrho
erlPc8ePPKWXf8xqMUJeTS93PeS5jz7QdzkdDdb36x2+PWzAPPLI4wIraF54aVCI
2kTlYFTNdUpSmbo4NGbbivFXGYKafYmYNluoac72juxQmi4E7iYNHXcPee1NPe6m
vZR22NAWFUBMhyXgIE/EVgMKZNCQpqSFoIrtVVlvWp/8LRJ7ZdSkvagRrhnI1IHx
yLZwP2Zhwk4z9Kdc4NQtInJ0YPTjieZs6xXzNuXYR0QsEHHZpSbEblb5LoyvAJrs
07ShuxbVtHkfkugGAp883j2rVzfFlpzuK/Y3+oNnfYsqJwefty9FyYr8dfVSQKqz
wyQ0my5D2EgYstSMA1lsS09Ffk3u0rnYbrJrhng8DVbKKz6WcCd7F5sFUpSXOtgC
O/5tWeqxulmgL4XFHafT0Gs07MaaUAKmJCt3rCuE7DWze1QG+qCjiINAfLFPsMop
EYUTOVS27RERXRIacKudtjlkxfo8f0idMNOzTPTM97VDkyQL7p4yOmraL203ynjT
aQUPHsVEDayS5CVTpNMliYdXgV+9QHQfuYCw3STFSFKsbTtLEaKxhCogKhfivymG
+L7xpith8Uq/RMnR7gipvrK2IkDfdi9Yn/LFqIouYUaE3uWhENfRkU/WQoDNX98f
9eXqpYS2yTGMSQD41OJaNdUL5mOova0C9z0VqzTfLIZEbZlgKTwXQyGAXw2O4H3p
k0+3jnOnid25UNH694903RfkkXOoZSzeS3Szayx4BYzrgyKa4ItH6Glanq8du5es
JyIBpUuDdeXX6DY2W5909Xy67HQwm+wJGhw/cYqd6oXpXsQEo68fF6QwfHQNNmOJ
4PpfGKApjHNYSN8LWqARG6Uq+mS74y93mFnTSmuWubjo1IsBOU+tSgyf3IV9/eTg
n32oFmrhIOcgFHUxXUNVemWRJZjbw6J1s445ekJMDpaXNuEPHghet6DKbnXQzMVq
WWZ98kgD6Wjjs6WH9Lw6o0nr5pE4huxiSJSH5kZ2lNcia+LSKN+oNS005AtRqgXI
XgGlU5elpo77jPJ61+c+8T10oD2beBoMx1fBL3RvqsDR8UOO86oGSqnZM08Bi/Dv
dg/No2dfhjlKcGbe4LwspKxRc9YoP7rokH0sKVOOpyC1nUi98eqHm1t5/9CtYWt8
Zk5hzngt0gmgceyx/b2IUyTIVqghVkpOWu8mE5ly+M6K3on5HOPQJi15GshZDhpJ
/dBOBLZlRvbBQV4AtrLr0WbNebJFqV7Ed9hwFa6wg+Z4sGBtPtm+9PLai8S6ZUeO
XUaIEkD7JBM8iDGE52woHFeNPkQKS5/qEm/fk3+cBmdAeEjJjXF3kD7K3Fnjh0VG
hDof8d+Cd7CFngWI0jV19b+6Turp4SPde9CbMuV8l9k6lHP1/c3Pv03eMaEwFR1u
EUKHUZhuBFD0v7WRYvg4TTCMnDRRdYD+NWdLspwEep80QB4RUrl8uK2CKhKZCTYE
NFUd/Fgq4v874Cd0AKV7E9LE8yjS2pQzmTaBzKRYkD3feiDxhDhiQD45otXdZLuR
kYwb+PKTW+mzFDYmK0dfiZJl3MbavXbI7fyqwGoDh5BTO4moij6RV8OpO9by+Uu9
TrVoTWT+2Vp7Tp1DGo57T/Rzy525Eiv+34m8OP67h0BqesVgCe0sKpPneLgykUTn
lX6pBc9VnrmOGSjXiSUx0g0/NZ8ul8H6VknL/cCmxDdn9amjD801MXx1KmqdapD1
XKInvVwrOeJWYnCzVqMSVcB1zlBRlA6DJRoBZIYSnOY9R31i0y0cfamIYQcBMbhF
GmszdtHeVEmWYVsF/1l6IcOmu3012WZtEEeAaD7g9x2NyBqm112QmHZjzICYQNGb
a2XE5SdrXBxTYJeKagwiqgtZNpQFnm8p8X/Pamol9LgL4PAUaBAgGcMo/nDKm07r
1beDQdePJKGB6tF4icq/Met34J1xmv8+GipFeXOYRhQxfKvPfX0uammUgEEnEmj2
ax+iaFBbE0ceDxRfu2Pj+heJqlngDm10cm91Xn6bthOITqY96ocziAnvXrxPzuVA
SOQ5nU13K/B13L20763cHOH9GNrf6f4hLoWN+pa5nuw1QHTxsDV82Y4v9sD3zUi4
TZMvORLp4qrG4q9uMkbZM8/ks6iyMJ5dUao8WS74qsp7eVcRxOgdYiDvdDocHLJf
NpnsWWWiJW+4+XgdSX639etLSJPuFKPM8NlIZ9/lugvXEcUcb2y+mg9HqwYoxfns
xi1VAAXL9SOyQWjWDgA9eqjl1U/AavT3FJq4Eb0d4z0NahS9ifzjtCEWXOERkYXk
NRVl179t0yZBQ++HA4qfQrz/lhox2r6hpVXnDbxX5XPJPrHrrFs5heCW3F88sGpv
DZbHUWXx9K7P2SvRIJ2U1IS/rsXzIYi11Sj+ykPgtIT5WKb2Oczu1BPx+xnWwW/O
BAX0/AfWhwzOxsVblgKNfzE04vm+6qyL7dUMS+pjfbrte1SpPkbAaLM0lfGnTKnM
XmVKa7KTJHlQSemXP4Oj7IfoTdqSv1gug01/E8AaQILYsUKXREXstfXUiYuNzCFj
aoYqRe7CLXdsPw/mWq9SHVyZjMiHHGxt39r5Rx/vW7Aztn+0SND+pyBJBOPkUj3e
+aa10kghDSeoPWM4xPjfyJd0El+ajgEgU+JEQdVT+yJ4L52RIMrCoJE2NBxvFlwU
CR/a/mh4re3CxprwpdevcSSNcRKHZHiFAKDov/dKSpavq7F5kg0ioAXWiFgDjRsR
25G7os77r8PDyoX4jCR5ZMUmJAJxPBfr428IuMgt7LMH43csh+lOOxr9hzCF7GZY
qLKeRiGr4oF9/dVQtZ206n8B+ZeggWQjjoYeA/XW/0MAptm4200ZDkl6MQG3i2CT
YqFtlRAsH/pJr6WwrBx3DcvUl3DY3bVuzOOy6t97GZyddVDBUo14SFkyET5PX51K
1IoWiXC+lg5t3wsXCb6pucbaT9khxmvwsWbr1CSAoCKOwwUf/ssF4jb1e7axhNAI
cT3xbsOm3v7jUazGuEs/F3d5hMxf3ySoub2QBheZC6vI0a6GK4ZHa2lTF1GHjnJq
anBnVcV6YnhMObwWwJtqkn4mTkGvu2933emjvy0CGAOlwf+zsYzVybL0uqtGC84h
D9G+TOiuSWjXJPWuGklnn+EQ1yKGoXtT5JpJrb1gzHBMmM6sOKHJqQEUWa0x5ckx
gcrBs6983Fd0OfSq3ZYucIVEigZAIKxH2cNBzNjQSJkQe8Kb1Z9AOY8vjZAlipXs
LixLlROCiPH4G8jVOJkARG/gkWsW9vHJw4AZrVr4ju1hOtLdhTjQz7ShqwjPAPpN
lPx8BmDgskNCcos3E9NFko04KLes/qSiiZufNtF8qDvGhbXtzGPpJAAbuY3P5Liw
ZaAMao5vQ5TM9zlF0ZSK96wP/C5Kh2+ifLAYuestFRjF7jJ/+sFspmI4c+vzCqHm
SJNhHa54+Rk9hD8rpUGz/O2Tom/neGmcP77sSjT2N6NSW9/k6rCAH2yEyQMUksMW
Qxa4BwbfwkvQGMWMXwlr5wdMvuytPtwHoGInZgy8qwXGbz1TKX8NcKbg6yxa8FBL
XpmfT4s6nRw/XFQWjwzadZIyVTqsQaBW6f4QNAvt1HN9IkpfsZb71v4CTtsSPAhr
bgRMYkQBF2ryXQDc9jTnqSNaNBGQ+P6yRYLOPULKDHXgl02E6vcdYR2CB/g3Qyet
gNerRnnfJmLKPObtQlZ/aEuvGwS/AE1kjLFM2ZiLgAIDXbtkw1swZfhC7PAVN/5f
MXRZHwIuHBKeDzHzncsWX3W5neJ0IyOhfbXnI1Brki48efIoF+6om2g91Mz4k/VM
CFmxNtRWa7aQIX9KzCnoRiIvgQS+v8H3xgHmQZEU0C6Vy9zt+gMwI2E6lqd+IWH8
bXT2fv3PwkG35072ViHcNO2E2dNO7nWuLflkcBfEsoqq1n/M62KQg+ozO+aHDdUb
N1O9z5/hMg/hs4T8BMKKFFmcH9S8YtTAsdWmKpi0Yu160LyilBlQQPyRqnfmcQ/z
KZmbmvWcWOFtC3jVsbuS3XG3HoUlPUPCAka7sG65EsNBFbfiDLm9hPNMU+HhDms0
iYsPKPXXEKH0V9EsNc1aTutjvInt2ZC4HEPHLI2GuUjyp/81XHe76v71VQnu1iUH
WLoadhEGrQNWtZ308MIut7fM1hj24jBPzT4HBiXOFvY/I5X81vpqrDMF2vTmH61W
XpjNJO5Jy8yiU/7TQ7KlbKSxVo5TPB+bwLlTz3W1pHFy+hlGckiMycvDErCk9oji
I3E6TDFXbuJ+S9fNQzt8a+d5lzblTIlJPJa+DBITV1n8CY/Pjm5O+srihNAC3BnD
DyQTD4qPaZaVJhuJ5EZpaQnSpQzswvwbeRwysCcOEclP0RDrRQofKTtVyDWP87fy
HPB2YSaej/cHgNP5FttoOECxB7CDa09rFVZVqsumwh3nkucYOyEbCOgdJwkU+UYf
jXXpw6KTJ7bj2xgj8hFdu9Qc69mI8jP7mRHm6/xNOzTH/T8Jt4cjdVeLsGWEA40J
+3w+vPBFzNcvGxM/mxx4/nPGHPATPfkf50Oo1FlAfCYwYbyrUNZQ2a9hOSVqUf4v
m7x5QIyiLS+wdzu5dG9Hruli6Je9E/EzLFmMEs+j2UmDbfGdUoh7muqTN7Bmb3Ms
0kvWvaHCZmRMf8BohkN9xiuanVZOoFA03IypAr4bgjbiQoHdGf3kXBWAYbs1OD5w
o8GfCI0lfWSP3ZA2Qn+WnioMcZTAKt+rTQCFqjtmJFVkf1QJS94N4DSf9V6cO3is
gPQbKAkM1pe+J3fuibaRw5h1BPt209thQdQ5pvnXsL+GqHNSTFElXOO9AVSzBUnR
NLJdAuoS+6Di0uNNjBZ+v2a1jVpx7bE/pcDgg8jbuJ2jRYF+vTq1Gnk7fXiFpRKn
NSERjxjY3ti0LJANKTHY5Aw0p16Sh3FHL5qCMWVQ1fGC6+SOs2LGMnlfmbclrQKD
Gr8el/HqlhLYsV3PYXh/lACzmD2pzcfAJVGnQTRCnQ06rjBlYQQ49g+SxwFZhk+Q
tSnP6ifbn2vB/rOfNMog/mD6RMDHAf/w1vRULVj8X4TLwlrBOijNn74n1LwyLyQi
viRgQp5ynoijn3mMQLywueHbRfbF96GeGz2UgjDtzk9cTMnK+P2JtJkG6HTVhSUX
TiER184H3FWfvARTR8z/2cdvS7t3Ui+qAbONWW5u4Ae7Bv+7NqA1eSalCnWzFs2C
Pf3ICi28HoTP5XyP7zafwa5yG+N8EbaGfYZI0wDcszDGgDJI9F/h1E6FAPiaj6UP
Y7WyXY/OX5TqHJfVVOT5OZEX3QhmcBPzwvxKlCLu+JFt+W4fuBDz5XlcYRRZBo3n
wrQHe7bm1F9YaSPdCmBMvJ+vkIrvCGrO8kDvswUOiGP24sflkDW5jSnad1yL59nN
FZnNCSQeavmm2sX3ETaJrq2h4D2s4W5STL30vNeDWkFYjFH0u2DkLyH7tDphwjlA
suHWWtzR7ERE/FmdnJLJ63n44RztwfsxBxR/DC/k8YHdH2YwhYuCj/UH+aBeoh9h
NSgW9YVmVODiJGwwJ5ViQo5DggABdpFdOtLJ6G8WUCInImvYZIqYiPqZomw7ONz7
nzyrN65GeeYhxMFpZoOWc5/lS/tvDKWmlSkKePHiBGWO4iGIbaeN8/a16TGJGuIg
t20FlR2RWtAMzkEqlpMjegRQnP7FTz7QmLZ/PXeuQtjftCeIErdi5VMynobf6lk3
PPAbMtd+r7KJjPHfTj6ZFeFfp48gWcBKtpbflUongUKzKLrZ64Gk9BH/31wPE/EH
TEu9BjLgcEYH/HuiGkZueVCRJ7H1h1IPpP5O+7AlP2MU4+RZEOtf2QFVVrTJ7VDt
Vo2i61/kn3TZ9rjx8qNX53/zB/+8lpjIv49lphenN0s3wzMbvzNDDEBiZEHEzSzr
4rARDYByeDsTaP7NuTePWUfpFpQ5B6X5jo/DP7V2ese7rCfzmJe6s0qur1jNReDU
fuvD9E6sMFGrWtwy3U8ohL3/gp1w7W/1jZy/woDn5dFiNnCwvKD3MAUg5MmMbKx6
+pwSgk53oT3KKcsdJfiPFmdXNYgW8uPd/z4zG6gaSC0R8GqejRRDjSz7F7UbuANx
Jda1oFoO7XzZpefmPO7T30fUpuUnuhzDd2t39G+0tPpKu+9qKRQzj4yxNMDuupsz
Ah2sPKmidjPD532k1wrVQebBAb2aNJZwBensCyrEOGiOW1+RhPloQ/w8D8DsQfA5
0u8ivn2L2nhTJIBckeOz0UbxSS/GWB5OhLM1NpIN5/9hnhUBIB24RFhpeKCWR5uL
7gae24YXnQ0aR1tRG0fxgPfj235hDMhkiluD0Ik7Y0WthqfUGs4aDbJuBxDbTR/8
fixUkNIQE0lWORKtXwfvL/IO9AE3T5GsyydKlZ/2QWWrz582KS9hOsWLQb2WjSNe
yRnSONi4nl7Z/rS7eMcYrS2YINzR4hHv5kOQpf3y+KzitlzJd1m+v4sj2nNjYVzk
UGsjvd6LLlpNWSzuQDYdu/4S2pNAXncsON6XkX4Gt9KmD38RRHoIJGkZ3VA4afO8
YDwUiiqYtEXN0/dpoleFP7lhmOw6jbB7cEDn15XG6ooSIVDv5zCdIUiYOw1hq8fI
cXB4VHzAW866opi68edgnbnvXA2c1/OHW4UyBURYrguF8jVul80SuMspk3zbJMSd
6orUMSmZU/0qZFKPbzhOFkxGP6Q9T7+4Z5ERr/zABS1LRd/EMTegZuXs20yVnxdv
bmeRveNpnIt3jjI+a7om7kt+UwFm4nu14a5bLWwv6IFumM/G3+5rXrlgqIp/dd60
BobK3X/+M3Uny+A7uGIusiF4CFokvXTj+5nJ35zs1WXFztQ1s4Easju+tcNoWPn0
tO41VrmC3CFXK5ZzsnSLoq6tRvf2uYgozsD30hVPcfcP6h6CjqRPPKrpLmy2FOvH
2qAv2YVv1Rrg8FxbLXNaiIpMk4aFJQF3nLGfKgn63lYz4tl7jx+lShxq8Fry+IsV
LHOi8EEMgKeO2xYg1M2t+Zdq0yDU3iEhMklRw+7IJDtjMVaMfoKW1EA7wQTqUrB9
taSHXqX6HKbrMB85O2v9cz8wQd2puRxCe7BCNZ4a6+lfagN5v+j/jtcUVvkUfKwE
692dhqnerAMBj3LfA8Lfl2iBCkV0+rdQsV2rAB60tRbJ5rchuLBcilWjcEJIaR6B
MPLOfdeJFXQBPE6U1oWeMyQ185iIpcJlavc17pS3gT+NI4/zlr8u2Rd0tLaYn6zh
Rs7Z7oVPSEqe1RIu34LV5MJkVp8u/vwEC9ZjeqVQHA6A33zLPg/n0aAKJgD71JXb
MzF5RShoZVK6FBvGpZ+n9Hs8+yCWXw8iUiI5R1ai62FRdCNk/cdpmxDCI0wrfX24
oJw5iBbIAwm/3S+HaqwTF+tvWXHzn3FNQTL7Vx20lN/f3wsB0HjgbGO/2iS3Z4ZA
wUxp1VYgsWCJC5xlX7h5R1SOR7xlysupqkdXVna6xIy5uRsHreug+EUbAkAFFf+3
veuLb+31r6FfaOEKhwQULE0ArP0Triq7OM8UOOBCIyBD3eKLlUFHXYOx1BDQFVKx
S2qkctka4YLmPmeKdlF8WNqfqCZqKKjigvxrGnymm7qNRITo9k5B4soiI6NqI4MB
j6fi4WTdTcahkwX/ZPB0oXMfFVSM9Q8D7PMBt0DExwhmbfmMDORp98Q3SZQXJqsK
R1AUshknnr9FkWyJ35W66F5blBx/biA7BzU2LQu6rlDKAx1DQVKIlJ/7q1Ga62Zq
zTj4iE8bIS7q9WEvCG9TwItVjby3RW51FUQ9IHARVXPFYf9v6yev3C336CJPL/vh
voXQ9tmPxlK8cZfVHeOB1GmRpEJNOA+cU40JN5zPmt31Fm7iTZkf05yRH+7smZQA
wL1+75SWE7AKMt1O5xcVarqE1RHyJUwHoWsm4MuhJ5YEdcgVv4biFIwj//DXb9Ag
T2iqu5xvf4qgB9xMevLiBZr0cLkHjwOntk6QNOeSvDanHDRMyGuuVTKJQGZgyHe1
QTZHVtRDuV/SIxW6DdLqDw6SBonruPvJDr3jOoqnxPJvsNC+r7UHsi2b1mJWqaOp
utZN30cJCzVA5ZxlFptd8o6fcXayG3NSC4hKShlFCcZaFNWW/C6KUl/EKvnyAb8p
h+03S00X/EX2s11w4jMK6FO2GE2jfOpiMn9Qr2NErUke4TfqlZA0hV5Mle+cEszE
/VWvSLcH12JhR7yWnaV/P+RymJbn+nN4wEOeDrJ0uOtI1NgtX/0AHhhytVZjA7LN
ch5RMeQLCXuxgRppAcW/deXVRJzm/5f1h8/EqQmsBQTm4tS1W8p46zcjVuolJJQh
E8LgpAg9aGimwEv7SOdOzfaegSn2z6+qUGLrEgUEeCaWfvjEA2EXC2Keso8Hn4qO
7z2S90CO8gv76O+Szsp5jgysyk4wiRTzNC6T6srkWywDQUktjjTlQxmIeH6fXSRf
aPVA9gHGJZOiQxFM8T2KpqluD+W2aIkUjlvIXTOi2dv9hWhAtoQogclHYRZQznZG
Kw/vwSn3wwiTF9kPR1r/ejoGLg5sIomW0ZI/yy5V3yIVSei0mXYHCl85+sXcsccQ
AUtU1BgYGwYGtFS+Mju144gJlKixEYF3QP+SILvaxLSPq49rCXkyLgltFxJxKDjg
3fLFCdOxomYpMlmcpvvX9aViBSYdAnB7AqgeCWrVZKZHBBJmc9P2+hI6EaAmQWMr
GSsMdxpH/F8BZuHjAVU1z2rOxXd60GRiS9C/aqV9eRe+pzs9HXzEOsGQm1YKS4Vg
U7+Nsq5SpR6TIz0cXw5/4BfUX13QWaanhEoa8ZBCS4DvB8kzG1lzBLoY0/iwz0em
a8+hY5KTRhVRx9es2O6Oh0FQS+uBUCccxix9ERueRZ/EKxxhNp7+5Js8BkvoP38A
4dPgp0oxhMffnb0eoOvBgWeRTQMUBb+BSSJEMNi5tnxq2mwPQvjbxITCIgrt6XwI
FUbWPgFj0XNjPEwd3ACyua0vk5Fm6zPItrmSuis0LK8yP3/wxa7Wjod2Q3Rmvdch
3AhzPaWb+XpSPQS7CNy0ld4ux4dHH+9F8pERrFS/GDRsTW/Gxpe1fCyDzAgWpWMR
Uh6zWjF1aaza65q0DHgZtbt1WZmL0AdHYV1Ce6kk0z9nRfsPDKd3t3if8IY42xl9
zYbvB162S+jK25B7xRHuy42FVF/i9lcFrQuj1KFBuxvsUQlPquBYsc932bcqJGG9
NrRSVFeKjHAM1bWHQJBEEq47PktA3giBQ0maKY9+/xEN2A7aAILvVf19STVG21hc
7QNSv1pRJLmw6nidrd0qLrqvdpNzfyfltLCaWawQCL6Ua1gF9Nm6QdWltX4aqKkX
XOXQzs/ivCAImxK9nZPCRDQoZp3JRtNRXSiAyD5dxaTLUOc5kr9NsD6Td8sHxNuk
lIry6ojpiJhhFubigS+eI8BLI5k8CGHZYRo7vgaaGYAmKkVZytunewW6RVf+m2Xy
96F7nOJWnm3JzAcFd5HlR9tZ6Nd7GL3G7yGAdNOO3ap3PwVdaY/2lHXf7m46p8rJ
zMLAzj9EKRKEKw4jLI9hZxKwjGiXNkrg2LqSQU62ITJqX17qcPaJdSXZuZybD8xY
DXUVf41EG5Rdg05Pox1Od1d+uYhSdnlpndsOVk9LW48IiHjdOQhIjZxuNWJVvVAR
8xy6ti5HpzO5F6fJJUzWg2sEMJ7D8hv3QZBgpob2Up8y1pUWHevDjmQmce0yORML
ZTPhQixe/ugfUsGC3CZA8qJnDOhjqw6dCCLbcljXS/NfJVb5YxUcqQpNlPxhzXuw
4XsqwUxcqcSduPCllUsXc9mF2pWojMJUY9eBiKUFOQESMHSz1dsuATUl77HL23Ux
BTxJp4NSydot7wHAYPBKrYq7CxjnjPLN22QRic59KWneiqqfG0bzYXXF3PQzKWrz
uxaLW2lIRvNIvwG57P+DE3cfUW6+X3W2WxJmiHBPCWkfq2Bur49Vqf3pkoEvy09z
pi9HJ6EyBnlayyhnLJIiiXs1TTcdI1He7SJ7Fbe9nAUJQvnDxRHdW37VHlmtlqzb
I17Sdo8sPzSPDqQMyviHvw//Gw+Up0vRCjtHprfidzgJFIeu35xZxy63xxCQI3+U
4pHRtJ58Ic18TciQkuionYNG9cbPPNLD7N51cZ6m/TMF3b0Onf/Po5Rgg8Ho+aAp
cKxQMY6YwN53P6/MRqGSl1ErD+KMkK2nbi6I2+nmLY8fNNbqzhMTiChSRR7tS/Cv
sGJ2tUQfi573aDd4QV8PVx6/pBKuznoWFGhbxvOaBuJ1tSt8VTl5RK2+XogkgXYi
8LA/9ytvs/sBcYNliH/kYq6VK6by2lFZm88Wn8jFYRAwOnKHzX8JTXnvyLG32u4I
ImUoCJZBa6yJst73Gfmgh4rVrFCZ5pfMDCWN+sszy3uYyPL+sxlZEkDhoWU/0+L/
9oJNW7RbkXf9wePQA6wMpghCvWmFEH3lrYNS3ERXebt8Y9YDfdUEkn+70lfw/2dv
iJcyU+Q2rN3NgVUzODTmtLB/dth9SnsqieiFL2pTEKqN8lhQz6y1w6FVHSXGgZNj
YzJpirGFXpZABs0FMnW0brof81H+yTz0nBxn8RyQ4V1jkMnO6mq1ImQoONYzh2kl
sGsmNugJZiaiH0kjQIbUBzRZiyZO/QEG6yUwFmYDUWACEiQsfoLIuhXh2uJc9yaJ
IHtfXA+7DF6zqhdEB0Vsv/shxXAm75SG5Uyj0d9SzxZp2+B+RS9PrVy36knmc0FE
DCoEK0P9Q905+WLbuUpQ/rqnyhM/WuKMS9wKIfsePbnB9Otna5d7dvZCVA6O4qww
8Kvn8t8N0fj5RmmZOSMEEkUg32mAIt80a70dIRvFc3YKeh/+ObRg6maLK35R8ssA
J/j+Qwy5EF6gTQ7Lvfjzmyt25pPW944gp2KAkptWoDJ72SGr8PGKxCoTqScXQCuS
mDNhrvFftvz1LzV80i7gNN2assruOYNH+59YTSbjLo1GL/8qQPjiUhQsonQGOa/P
471/x5uEreVHrMJVNRcW+k5Z5IcUpji3+ZoXTdOEezARmghrAgH4HUbmbyu3Iodh
VEtmx9fe+rhOu8+hzeW9jQ8l8M6eCGWtW/JRRH9EQoGARwPeNDJtOAsVYuKB28V6
XALcE7Fu/Uqhv3uR6A5US+KFuc6tpKqhrFTicC5JGeEeTZAU166FsZglC2C9BwJG
6N0qGOiJkXk6ucmI54CoJ0/iKdm79joQuFIuaF3aHTovDNfeUqna6lIOG7AtF7Op
5KaEydRrFEnM3IVhhx3Mm9rDObKzBaGGdtCWoJmDi6qbcGFqPEUfswiAU/TbcP4n
rC3Zy31KcJo5zNFT6ZD3bMTtMQgxeWKsIJ3S3meYcX0U341jxkYKq8muwrMeIbqu
WiqUGvwpqRVZ9acPHRCwt5+qkg/UzkQlzTtYVRVR2yG/xhV1T0P0aCpbeGD0E7B+
fEsbnEsKYj6ErejtNmlTSMoSIPBmp9cPLkLkEmHwTwvsWR1UKoy7BZ8nOAxdQTFJ
DPMwqB18WlqWxybIXXZXSCi+ZtwhKYj97ll3maY6gdLz6dTjgju3xQRXI0731otE
OG4TXWBCttn+ZKlOssXcFsKza0mAqDm/RH1vG0RPknZL80W8hqJtxteh+xOGBM5e
JZGemxGHME/jqUbY6MhN/383L4z0qg6+bwcpozhweT9pyXy3XZyoOveMaolNcdq7
peeOwD0bGIHEMFAQ36ly4QNGoR3oq9kUllv2X4GHhFnpQg3WhW/4LEI6tdWCX9NF
Dog7pfmPWYlliYdEZAuPFVFEbuhpain+E9jGe1+oemE23vku9B0lSX+cYFTLgzgZ
LUzlP4TQPCvyjmdJhTCHjov7oDTQBvD8QChivABADcRfrPAgF9rhCwYLsKucwJFu
eNbXIsLqNZdxr6MdRWAxw6Z8ePVDvKH/FYbOD3+/BOLpT+eeAO7Bu2rHwV1DRJls
og5WZq5+T/u81+/CsozuXxFvP9rc+NB7ujx+YHTaVKaCybubQ/HBzz5A2GMLyL07
nUpoZKpKl3E/SHyjsx06+Pni1AAvBw+aG6p6qZjMlGGvdEumfWPe2ZIssaKK/Mx6
FY4uH7ybrw0jOvBySVkMkKSfRTdf9AvcRf5YRY53nRlhiL3SYjJDcrPEhXBf2zrA
mEyAD8WcCzsNxT4ZMMYPc7PGU2rgbESffRiQOvK6rfVl5j3kUhGzPLVFuOXhcxoI
Ssel1ucDNwrzyPH8R11ru3fz3ssH1CDhFhfNzzbEuS59itXFdAWV3Y3oTaPz0Of9
/s5kHxc4Otmr/TEhH4gkJu8qiulG9G9JVVc3dROwyaHDPUXLoXfO5KfbacAKe1s/
fgbRwT2wYg6jruXGsVOMNvPKp/WuVCr05nx8yjB4KKlBpko2oPE/2a5XJ4XEnQ+i
Yk8DPB3kCTX5pi3UGVGoz5Icy9Oyyl0uo1rYvcJd6GAdBkXAexCxJJTIm7+UKneC
A4RrmGrGxkai1kCAKvAZGIRFhrqptNf2RlhJeyxMTQanJap/H38yiVrBmfxEQ7EC
blQhTmWNpAAL3/y8HbtmCyLdUDI9FPt/g47tOnlBqXEiX8xbaG+16efp6P0zyPQY
U2+B+9feK2tNNEQ/B1o1v6Uvg+DWGUvMV6nQG9d5/xcAykmTzBCAfQWHoJEvyubU
QA1GBKRruJD9QumftIzIMSI11t34ziYVP9SlrS2Z3Ig2cG9NhmuPnOZZU3HtmLft
wWlRM3QKXv1tlFdrw7QM3EgFUOyzTx5YTRO8vv+4Vv0nYjDZVwODqVQGY/OHx2Te
H8TQGjQaW716VrhBZYbobKW20mvE+RRSPsOqOBNWORH16YFdlCk7xZxXtPm2oCjf
9mqy/KEn49SgWRkmeptoib9hO8IRRHftiwHZ/GrQj1yQKO/iMvAAnAcRrtSrDaVO
I2QDiiS2+GW3MRqX3BJAOTJm8oz6K12Abl9Wn/3/Iy0EDsAtp+3OyKRIUMf1MiLL
5viGNdNJT3ryEhpqNoemkK4H75guTdcweWxa+LhJ05/ZpzkB7kjKo1AKspTyNTQz
RAmTj53xUsjoMu8byVKzqDpqwGcBBPd+qrvmj3YWHY3DPcRfsFU5tJ70Xhmn6EFU
PXFNyHLwoXI6YKFCIakc6F3Qj1E/9ZokI0Iw4vne/LTutqqrCRrnPzGHWBpD6476
dQnmZqXQXLxc17llKlu0OA2DB/b1lzpSiQOWwjqGZk++We2UcLJQRciu2MHiqYKb
cTnd+/8o6krUulppKu6tJU+bWB1OTNZz03+sY1gbT6oIZvoxBDAWnXNL2Xwe9chr
SWaKWxw3SP189oNXO/QXJAUYTZxquC5YgFolgVCsIqXc49PDFcee5lcnF6WBDw0h
j8Pra1dzeyJI4y0XhjnoYbiwJvoGltwLiiWMcXsP+nnaQwEeSDVqEJr/rGEmiOVs
VA9O2sOQRPOKpwtboh/3jCOn5ulR9n8I9zhmZwoBynM/2uIecXOIjyiK1m+sepI8
Xkg5YTYJSOIHXf1Qv4GvROvn0+NfXuB1HQCK6Tn6oFDlHIg5JcTPi5JpcQmIHPYn
OKC9MfMykhPTE4PSwdZjhExzi3YlnCkEO2YFH5NWZ9NA3Yr8nvP9/k9qfRUJ+9jR
Al+BCdC54G89Pjy7HCndZzkVxENYf37CgVpRXPPZ3TSSay7pQrcPCdZuyhLjNaDQ
OhQ3mSFPyYAgTPSCsXHnxT0mGitptDLfeMSXhrXFcnldNFuqUqIV+KIF82RO20j5
SEX9XAXCN9FN5oLAk2LvDsIt7Ich63bPyhHy5m5tW9fQWK/zELQDVU1yjxMH2h3O
K1dAH8LnBXqDzoRn5MklIYoCJ4UpZL7/uFrBWEEGEhC68/ewCCRjWkIn82rwZX/H
1K+VKTPtKV6hdSG21cU3vQezRjTxAgaTW+nXCNqveOpG2qF4fa3Td6z9/1PVr7Uy
lxn3P7hMr2MdTxuEjYwpvZlT1Vpk5qfWkXcvuNWJ8zOdC52VqVLwTZRBb0BBusfH
jls8gmAjqdy4e0Asu4Ysre6y/HI6HRSj+T5A01cOukdgx8U+ENCSrRdeL2lJFMTw
HZVJwaNYJTa6jS5jUU8f01ryGo8GzZNzLHGLW8HeUvFmJDWqESCkNILaintFaDv8
8/IgRILE7nIJi/J9d0vgW1g+OzHSO2Stvf2v5s2h7xowrDO8i28OmdJ+h97oKvr/
rtR4lDdw9SeSBecC1dl3tb0d6Jn5qoeo0XnuWUPHrm0Mv1RyOJRP2eH5ShSZx5B2
IhnUxXVxHK5d78E4VpfoKCcS61vQCA9Cben4YuODJ9fYmwIlRtu6h4LysqFEw5Ur
+CdutxYPx6j3VZf2cHBNrf6B/dfhlRNJt5Cu/iC1AYskx7nxoWGkLJRHAyDa4hbq
FKafJtNdWpNlk64fZfucfhosyOAwPnhVOHCj7cgOvs/XXD29/+Awm7AG7cXA5ahz
kCijS9tIv2fEOCBTkpk5A10vd3SkTQQiv2e3+FYwacf84b0OGt4902NNaOnWmxvZ
I31wLl7Fwko4YEGmvszXIqVIEXSWEv6pZvNhQlG7HUHwjy8po2D4kQOVFLs9/Wui
Q3HYAArDtiA5Y3HsunJ2Fl2RsYNPXU6PunRshfzww1fXE24AERcZdVdTCBKbEsJ/
juonlmk6Fnv9SgJDLzQhHmfFYrtpgZXYsxqFKtPomyu55FUbrB8ZS1+GgQNY92Yk
SHUTwpOdOQSDlRBtmjc67mZIBLeVxpodMvOCMTWR+7kCL5u3OgbJ3kBVnCLLtEot
b9WWRRzbDDkJhswU+hy3br7nelk6Dw3FCCwfTPIY3nUpTR0jzviehQH4rU0t/kfS
ZHyMPgYo4IH8M+6n7EGbyp7oRQkSXsrMmzrz9gBNGgG8YJlCZB2OGeyMDjCLgmTh
n3cZP+myav89T9izTd8sFBemNK7d9awGKUdmlrz7JmdQ2zpt6GnGVqzlQ1bZ/W5d
i/0vdAERvY5gBtgOrWuMmcbT8W3VrVZqVj8CeRYYqMVeIr6zxZPAs19JMsGtyLL3
g/z/5uCnrInvyF99nfR2q7+8xdVLP+1YVC2zPo2nZ3iJQbikdUcCasz9rrzv5/RV
A6ZVmU2hNi9RX93CcVw1v+awNnyCMcoeTQ5Uu+BD6/vbbziqEfm0OP+8/VbwGJwj
KycDT8OIR2HXjXBLInBm2G4zoak+bBQRaD3DEdtc9m2UMGprtHRdQzv/njliBPUd
FxIwbhFU9b6Ib+ZqKgPuL72ndxpDMgTs3wRwdwKTtTg17nYJyY41iLxBIzCqxDBz
y0pyE8vSB/74nD2rr/EtgJE4w1POgX4oJguziQSm44+jsBhX3EpzqMoPU71hQKK+
9vMPfwp+V645SuO0qw1W4LJD9xfPnETMWOBNw3vkb3vs02RtL7ukPqfTgG7oRjsE
6D1akVdQNxotLBHnm5kYnBOONQQjwUvNW5soxHJopq4hiAaGK8N8ZuRdwpZXdjWf
S6rudM8Z+VSJspZW9xxcx4a71+X58ongf7HjBYIZb5qzBusPknzjmH8aXHec0hmN
3ZJwgCWpCbZiR985rRPa8pkZKiv8GTYBrHAFQR3DHr2xIuswt7dH4mrjSJM7YzuO
LMnveW94wQQ5T/zkP6zbmOhCAbw4CZhAVl9UkJUelvYzTl5izq8k33BlMJMOchq9
SjdzdbdaOfPXHF3ns0MRpdltXfA4b5YvBYnavR23i4se+M5Yrf38v2Knj6gpyx36
cjSJYm0oz7fJ9LD+IUXggQqR96oMHgPtHRUUCmfz7CykibPq7eY5hJIbCkCIxwPx
T4VVFCtgCWnVABsUKBgA7qJ2U3Or8RgT5mEeJGOEpXvn19GCjkFm2fgy//pCDPtV
dY6dK45OKAcgX40UTqPYYRxYMvOqVIk5BJ1XUmTQQjQP8s6nv84PT6lLLDC/nZG9
K/MFLW7LVWV0rVFpL0oySW5zwaM/y9X8rBRXVZZUx6rxDBCrrU9rjaGGXpbOCoed
g9yVJS118vazeJeXvaov/T0JSsgJjDjd07lmCt1hIwRpcfvRR0Zt4xBd4BkqIG69
LrsUHqHXVJdh5RJxFOFSww3bxKJHm/bf0winsxGnK9uOLZRZHfm56MQIee4IIzta
6qH4YEs0R439LHOmM5fzK3CLPuw00KGLH9ajhYu0jD5o+vHiA1QO/w105HF0xxZa
fA0vwDyfF+Z282IWfaeprJKmrBlySTAVGbZK9e9rjvAcxDblLVmzSeL7tjLYX2ue
vR6IXBxNMBW8/nbaRhgrVOb/w+fOkZLKRa768kg4xJmY0Kstxhd4O7UYPxMH6bKI
/Li5HMUgxDxVNxYAu+wum/hYNDy8aV8wdklaZqPcLyGy+4Cdh3sfOkHEqRz29ynm
XpUcaHx9txXpNJp7W9dUeUd2XCff5jz/S+Nb4OzfhahRfpHB/yZLWcvRfouZdt8C
BgaqTW5cW4/7NlvUbXHwbWc2zq0MpnMh25NRW8XmKU9UG2z5tmSA1s93qh9tXcqV
vef98s5I+wko3DJsstUMKhyQKBYaygstRE5+YAVSBBdEhTVPZXa1ii37/ChwFwBw
2lBvKSk5wD5Tauky+BIkfv5+i3S526ycoSea3+5NcViJ9hWupLly3gVtfU3MKnVE
ulaawX8IqzTeah9yROl0r9jmbgqZ9XQ3EHnaTaswSZBo9DjTzHa/NyfTnMFLyCvF
OfmU5yxMiUmM/rY5EYvZpWHYEG48pg4ndNy1NwKwIsSYgJwtEa9aC18grpUWnj0O
LrB2ELcg31AHlp70xSoMRWWHRvqXwbM+j2qR1kCHe7qkAEy+RuEWoLidVtex7VG5
ShF8H6+urIi4rXQ/aghMrI/ShNAm31AQzjrQxV4DWYqsBXnAnqXRKXABDhwkTZ0e
fkW1/QFl//625ly5a+FwURdVm8YSqXjADBfBdL+pycJtZSeYTNmH8B/b+CHSubdv
pr328UUBqBmVFlvGaiMF6BbNZ/tzIhmHO3edG9ViVoUHxMmrbrO8Vp00uMVuwReG
Uwnm8kITQStSLaIjNHpca6YZLusbMRlcIvdsOvdCVRTnpwqYZGk9oS0s4ninj2ke
qAxYahxkrtLxgALm9ZK304YrS69QlYyj5nimD2kDa3+xH2y8/eVVlhZbfdIfKDE6
VIrFPIRcHwStiLTZNVp0xO2+DTGWnWL5ygi75DIuGFkRk1dnl3/YodQTF8LWR9ZO
eB3o2377Ef6Cqx5TVfN6GJgCcv7ysDKU3Ui9qLIoq2ky27TcHIxB6I/1QqLi81bB
3C8Q0EV2vTEHGezsX/+tsYUE5y0g5rDqsDgkOKJpHPdnF6gNhYkRBsIYDdP0eWUt
ojlUiKeAQNdXcLuLB76K35Vx226LgzWrYG4freZ6aUQX5KkucG312lYUF6nUJXut
RPa7CNoeakaRXigeijlTHGshetBdZgbW6IXyzMFTKiOkEE9kDaxF7VQfZoipo3Un
7XHLqBqDEQh9Ef5aMYGwQJIKcR7oGO08m4Pkt8jX0hPeDUDuSgu3pIUHhAhbISAF
nJ4x358yuw7W1BxZxfTmOdjVMsczP++U+VGU5OQUfqEQaMkpAwBM3G9z8or/Hvof
y/mYAU+QPQl2WzIyWQai2zamSUidOn1jst5E9WiRC31iNGJOXc8OjlrtL+qPJEHW
J+A21kPe7l9oKKoAfEnbvjo+sjqvDSqMtDthKpM8+ldPz91oRi3mJtgpeb42MC7I
l384yzPxJ/p7kF0ZlMv9HReiyYPFLm+ggQ/hNRen6xlnKx1zE0cnDpNXYN2QI4je
gRKuS8e3cwQ8y7FQpeLYl0nT8vP3X4yKpsbAObf5l2MiyWHtQoAkfej/YoN7shJT
ighdSa3INo78CV9d4x59O4c8pBltUxLGwg4JlHHq2Vam9JFhmrrVwB+CxOfCMJAR
bTKQWb9b7IKbhQOMvS3FStYJSOiLsst+DwFVs0rgk63Rs2fB1LC8KOggdOoYmeMB
98sXJDkx8f8HOGWF3a2nbe814VPxRiLR4ncK3XT61VwwBTOgDtye+8gMbUmvF3LB
YALH8C6i1VPXgtAoE2yhK5xYdxYDuJyDXTd4L7pcWEzPkuA018fjPkI1AfMPdifn
kiAQRLX7H5cLlB515Cj1v7zVYm9w1qcH8EUpAiEAYHfknJpjIRq2CFdA7dorWJSi
fSpYHfGGQ2tdVs5SAhmfdq6JClOsxDYSIlp+g3NaJ0FWuafiIWM/aRWFnJY34bjQ
lRWlJBu+9XZ0ZRYeTDDbeL4sHFZI/qzMd4ZB0FgAd3HOS79ltPq7qrCbysGkzBEK
1BTEgfc9TVEKEijjWDs7EWGNyqISfm6lraENE1xp0vtTxyDkkT89rep1h0P019/e
I5kORZ5MD7lJbG2tJ2gn2LwzeTv2CtJGQYxF4NgcO2IPM8FGsVPqJLsR39oxM0AQ
Dz4buRCmfjDCaUVyIRCE0jg3FOKKHrDqj9FH2jfKPTrw/6wJYt/wiwkwvDTOfcpL
MMU27MiyUEdD/cX8HjTwg3Ekg/1xRu+SSWlK+skyso8N9/nVoSlKbnWfMKmnk+tv
b7g2I8aQnjLBOxDHC/VKaFz2lX6R6cdn8YUos4ruGNyGXLSwayTxKEC4qp3TRJd8
h7yHcEuH7WPRzKmaMwXpODZyxYIbTUIf1VAW6c16iIf7E/0oIfMLuOsu8trR0o23
v46luRsQMCEXYUeya+7Ris9osGSRQ8eEZa8RbhG8Sgmf9pEUFXUVJkFtL5JAqqsl
cpB8zf0LfIhfBmPvxAfTKaMp7NbM2n33X5aN7ASnWRWBc+Ov/VGCkChS+yp1YHkr
Qv3N4QGoO5aDdUA2O2fqrkoiP2SDfQW07fP7QBRjLrF468QQSU+TJ+14F09Uyp/Y
2sUlMeMg6t1Hl5SXAXhwowOBef9Cx0X/D3ouJqzcpMNpD/95KPruqk6Ch+Urt3M4
WFGoN2jrEmACQ2Orug8DEukMzaj2DEriz0y5Sa+Hw5zNS66+NY5WUSPreDd98UbA
jYtdx4ACe1SbjfWycUDsjPVfNXdUx8aKoBPTI9DNN9o11uAwuQOEOswyPHFlaut8
RGoGMHJWNOqtln441+GxLo+cUnVinaQTkvkyiLWjKpHgd7iC9/oJqJMj9fubxm+v
4kpvEkxFbcY6NOpnTwZTaE1Us2BXd4oP1+SJhwCl158K5ToQbIEGgTlZN+JF5zLh
k7NpiqNlrpyoQUk2NtitYBaKRWXg3l8Dxb58kxe7ha3ol314jTnqcYCu4Npz1X1M
QlBlSCffiCVtTAYLDch5LUmG2S1vVzQI7jMk0VSW7Rd+EhSCPIKi1QYSLwzyRbim
X0bphrNodbSTr2BswZ5E/ma7WtFqbbMPr0DSuPPEtoES4V+5Cn1xWx77CmI/HlhQ
4uqVugRK/U//3TId8kfnImENL2gV84hnjBz6jITj22m1ynSGgRwHNPpmxSykZwMw
ncZrIQSw/GWJITw4nAYC80m3rp2lzJipNys0LifymRY5DsFGCST1pp8nlUjIUi2e
e8Lb2MtYXk7a03r3PYpujWmwErG602iSgnG6ng8htdNPzGJPsMocKFHUxI/n5OHc
bx+AjIwac5PvxTIoMo0mQYO8gio1Yyp08nNABhnTRuznfck/QiX70qRouoS0m/df
xhjtncQmHUznIfoghS+oMFLACZhmvovtriZCUvOI5KrYtc0puka20DE2SuBqimAx
aAVr22XgBtYmitXe+hLuiveD/4o3fFO9Ieif2VFOSM4LdVxltoNF5kB/fyITUOB0
JE7Az5bCsE+He9on994tGIfV1H5Z+ic/OLM7r9ab83p/eKQ3fVdRt2ahHwz0yNLY
JndOivYCslmuaInjE7bKsyBmiFHW2GD2ByBDbXm2CqSCzN6o6Xf909UJmL9UNrN3
48W9yeDBjkPDbuqbJU74yPb/OfifuT5iSFCIipCUPkA8jAanpotzfSWP8egrkRoo
I5FHYaX/uvuD5F9Kpba1KqAeQJ8tGsj80FIrhHO+kLKKhu+Lae7TzW4yw2V2AiRd
5QA0JRNiZ4odcEbF/aW063HFg7KU8XUPCmipxY2PY1Qn7rzxRligxflSmz3fVq1+
xrCegZeAE6VOztQtIETkDmUQg1XwGOLJloyvsDpYPpdUi420eYvs5ImKcqmOC5J5
estzNq3KdCUH6V0nJfttk56SBrc9dW6/MIvUwkO/Dp/05AgxP53E4LzqxHQnOh68
blWgKZ2/jNI+sT33XBKX8LTO+fjciLPEk9iGpCv1Fibv3+WXsOyOX1hOaPpXSGiy
qWofZEN7nKaPnEINgD8u4vkfCW2+PopyG4INnL8SW9K7oXvIgAgin+VKU9l/5pVy
eKD0gV0JpqYOm8CPikAaczYtkQ5nvgRVF/oz55hc90elOHbm0y4fW28D2bJTVqKo
2ilccRJNBKuAmgPfFkHZuuxcdeye2/qLurerdXEs6YJvMYM3hNsetsSvFL15d0tE
o2yYF7E8utjSrU6YtFG3aUAJuRBTuc4Z5MdX/aQ2y1IZqpCItsegvWRkH8m7g50W
0MUFBIEHRvt6qCxW5tGpaFUHoVa3Y6o2wM2xCMal3EMurxH8IthhhCpIMDVnYwko
+2QMzSs7ijf8Ssd3R/lLbiRkj6ZiVZXu63eAwbD4FFN7Eun4Fa7mIzMT55tBxvCp
m6sy/2AL7JPlkQHo3Tq+IFra644niwbJs6Esu6guCtCDA2blDgCn4wIcADCauEfg
NBLwukZBukdBBT3wavCEEPuUyjVuyP0Iy/K+l+SkPQ1z/6KVQ4u0DJseAB42G/VN
TUGpA+uvqk3i6kMjYjUzp1wAgC7Qj7K19Hcv4JxgT5EOXHi2Klf/PBIF9WyOzWPs
irZiuf/5mnkaZPZdv5I0afHs8wR+DO3/4YwTe4snTrhVE3UTkEFlQbDLOHuoFvjF
odtzXMfK9MzZf5mqWWd0WjJC6aOiCL2v0M8C+mf00Ib04jLcU4vNlhDh2yyTPdEc
8d+oub1ZvIi3S/PJqhifBURlOaBbkLouqehnxw2zaM4dO+s9bVFeOYkiw6GwHZKH
I+VxW50qBkd0RXs7ruaB/5FLvnHfSrbSlJWdbEUqH+m0mZkv/NC1MjZUhVsEx4v8
W92Bm/6Ydqvf2yLo6P1oWCXBpyYO+eXvjabvxmYmwcofEXlJa9XFuaTQngqNESUK
mjAQLG9diGvrGNa063aNC+0nQlWaXSiykQkqJP+Am0P91USmIYk5TFF9ptteI1FN
uJBldlobyHxXFmQBgfiy9u1Wh7dk0k0+5EcCmPckJMF9t5TkUQlRBpGW6KubtT3x
oTKbsVzmeVREy201Bfu2niscAtpQeu2qOgtM8GH2OaUWOYsYL7C4EvWTYm+IJwgt
TrCHCHjcLRpbTDis6BwZ2ARXmSIDG9q1aMoKfhQMSf8ROxpocdJ3zvBOROkA7sgN
XChmgST1ZVuEvmm93VXvRaTGJcKB4vKTQZJfYZLukFwSMpMrCFxRwt93VhH+q4ms
dcVIEPVKgxrH+H4xshrxuIaVXvpotOEWvCKpIJD8yfzU5FRQHc/0xPJSlIP/d6PF
jZMYPjLe5Vi+zJwx0PAxWt/iHUXUBwrd43YV6uxqRB9LbvOGlXdZZWotxxgH3Yv2
586fcwp2IsDfwZpzL/Iqs7aFO6vV8PHDvhMX1/3NFUbmOMAs/sbXF+v3C8EI7SOl
og/hExBHv+hsr3PKNjURjwF1elX9c3f8BkbImdKR81mByzTXoEVY4K53/kCyYyuw
KsSi+o8Z6NZ19VQXOwmX8dT1LdIM3S5suuO74ow89Jb42j8kIkc3zuNS6NOxEKsf
yDjFCebM/i4XRJLhxc3NfsXchXMhCDcVe0QhlgqHvcmIaSqZpihvFy6odQ4BTB1K
RRaofVfRT+5iEpFpKx0ZhbTLGZOPG/ohAyCVsnFyxt/dUPlx2AKnRQjOtLuhBC0E
BQI4YqQyHIgwE3NSOII88JrkArX/kuBjF25xO/+sErNjrPZ74zYgeV2olL4i6Pik
rzfwVdV3M+emvddp/A2ERpk8fTqadrjqVUc3AMbwtJC8vgSN8+74fOyagmdIR445
ZlDP9iYl8EUyJNnLdTaTvPR36ePc+sBodlPE2HOrUfaSsUhJVfGgd0nrf+S3uHkG
si4o5Ug74dEJIvQy0NQthioPWgtrFVercUVZMC3STXsmJKJfrz+f5NXPRwBtbWSX
jyjfFQY6RamiWzrzXVTS1M+0d6yMV2cvKt+CdO9NoNqwHxWdqPfylgG3QYc5UfEW
1rwYTosdn3RYxldFEVywsku10v1rUIjyOHiV8am6B/6KtAZoNkoqS8Px+7Kgcjl/
9jvxpD2q6Qqj13wvW/R7Xs2gAV/HA3llCWX+Ke/JXI4y770kjOovid487Ew9ScYZ
V/8MCr2W8q9lvaHEOIzHqIhFWC9M8nGDF95FoHyIxPys0nnSaILYMs9w5x8WcmQR
fLIA93vDzOAuRTn/TYz4hb5P0V5aFOq+rixKcW3p72GCVAOSJM7E5/dn1Wocild7
SJEOcyY8Eo8VaYITIYnwfSdnVQsQFN9tKLHAJLpKrfoz+2Y7cP3J6M/Muftdlnje
euujMY7g1Sw2SIh+FsE8KtpY3+/AD3fC2DaOstIfwxPHzwCi5x9mhHsyemeb8BXQ
CYKFp4kRD8eij3//YXwHvJDBFlkwUPC6cQoXqQxsB3dJCFBRBjleB1DXlN+rgh7h
foPbE+HlJ2CJGGkDWD7YUKsp4WPdr6rzgGFFxiPHyZ42xBKf/1zjrst8ybJ79MyM
Mlr2OppX65csdKJbjziIrqGbroGIarzQyuFhYxgqJII1BiOzZgSJgrU+j4Kv3I6r
5mdR1r1IOFHkijcRCKqS3XKWNN5Az48DnH2IpTqtfI9xtpnKHIGxUothRCM35Pm2
jB3cgPR2US3s8p6Vf0fgxZzUo2B5yGcLekYMdTuKS+EqRGkBPipkoPhddRirWAID
5Acah6TYz6g1OdaMhS7nKo0Rhb9BnH5zxB9yRxg+Zaxw4daQQsp+D6U9fr/+FAPN
AVkPC8zurpJPU143iIHapin9pykdcXpVYoKlMkkSUGLSTiqk1qSxMfNR/rKhbn7O
dn0s33iW5gHlsBQE/CQBF/sxmAbajwsZJHKG9UfSddlzi6m5uxAFaf6unohwAvxM
u0JPs/LZmvK63dh0FyQpq/NocfL01OemLSYkg2ooYn3mEqAc8vef7d/FRZ+M3D/S
OwsW4tO9xEoC7fNWQ3C1xu/iF8lmmDgMaGMrWKunOzKPMmKdbUDaLCMXiuusiAAp
IjL25YhvcmOFmv9KoDReXWrL6QgoVDvZpPZcGnWKJFJUakPOEKJMAbOr3+LIyJFV
FJbOdrzxueBX1+2sy4OmUW/wZMJOEmdADRf6HU0romerFvCy2YN8c5P+3HfJRXSG
CVv3hVMaavboe2DGol7jKPZM3YnrLKToD4uo7Mqo2idr6+WZqDP7hENZrvrDfdyf
2xNVXAHw74UdN1PVrvT/6/kFAYrVIIf4ZeOiEgOz5grAA5HUDurX1t71JPCjB0IE
VOJWu9GZDg1OWuBEAEutja6ySuMQf+bhzI4Br3/VumadwjW9Duioo+QDfzNjRlne
FOn1iUt4247oHnLQD5B6hSqJV3wQzRelCS7onVY4s6Mm0ywMvHZGq4+0JXalppSX
bbwE4GV+OYLtqnAInTjKRX7lfZk0MruGLxmRmT6J7p/k64ZgEpbZoItAH8MhONHu
DfoNg6+2osCKQQ6p94GsXhE8wA9z9/bOp18ydb9CbmvTD+KgDu4jiWWngiS4Z34C
7UNDWbXPgtfkpvP1ZOuUAHEh5MLuyGtBsO6Qsk0s0fne26Bc+Q5Ss5AV89Uls16O
dpTHANAv3cC+n9Fg+FQ+Alyeg3SDjepjRM0OgNXRekfK53JmIyiKj/YR9J6ho468
pKbfgVGr7UcalMlQnQnuhdzqsOsdN3xPk+QHGKX8eW9mxJc/7FdSkysFKDNtfkyL
9/PD372K+7RMYL6TVVuwmi4fsqTf3BAIQ9NX3sbb95D3heZ46fwCKw/7/PmYqLhZ
E85F3Joz2QEpOwbt756bmNkn66vQoyDuz1W3RAqF/GZesVbhLEW6pvAPf3xp9E++
PrOCMOx743R+CGgINplsll8cUz2AhZsmQe5WeU2hWIyWstazrmb9knwuxiy4Jnnm
lEIVDpGIJCES6b6dg9yYAA+k46MK1uEdMkQlAY2QojlWS+BM4xzkV3bSBAJtp8pV
pyTsMmd7Mxr0iVl3ydzjOU3cKmrXM8xX97vkSA3LiLQcNWp2cTWAePmhc8YrBkAI
dxV2bKPUDfPyBirgKWN2Vq/sPR93w++NiWtacD1Y/oou6SkegW4zvyzZY6McBbDf
/lv1HGXAeEHFW0bgq2c3nEiOsKfCU7dVQrDNtA6V6rXPS8Um5lRjUGMGmJlnLUSh
TmgaAS7DkhIn/HRMLk7G7NODeV7YjJ/wnyHsiJ134D6eOTbgIDhhzm+10qlV2A7H
fv840uEVDjPHS7+lro9+UvuBlxl1W1K1XOSn99dCYJcNAfKKL1dQ4XBdHRTfnjpS
fanwcpjK1fxtS5qv9MJ6ANP1BciL/qeEKMq91X92FnSH7dk/EoVd4KSh5MAUscBh
Sr7WcpaIw3HhCPrDkv4VvDUjxtjd/Hltl+4FIigA5e2V4MnMlQ2LcU+eG/xS6lup
qfxCnR/FNLvhqnx27neACR3sXy4xx/bRz1qfd+noMo83OHfVF1aknIjEZZ1vyiai
P6ZjwJP55pBsSLhML6LJFgWhL5oHhi6e70fOcZGtkPFipboTQXESVYwoOpvF8dVh
vlATZ5BktQvsyEjt2YXHns22RJjQ5ewxGQMgsfGQeHf5nerG2JWH0CgDi/ZlpyjM
s/+trtkoAFO2K1a5mpOxmCSE4RAbSK/fpa6k6zf19MKb8HXBt7mHvIJY/Tlpm556
wE+Em2NbCQvsmHkKK9jTyHx/qIgR3DHY4naPoGFzU/rxPGHrz9ImL2iYNNUnaxyO
46qeuFV6mLViMfvaihxAY5ZyFH9Uf9ZvEjPIjYFgnWcD2ad7AMgiFzjfeKBr/uqL
aLZz+VASYnmFP8nxRQ5G1MB0SSEiWd9oU+Fdzc1HELBE+1jRXklJalYi8chXvJNV
w9ZeNE2QDxd0TU7nlPuGxAG9P8hshsQjYFzFLfOskOQ6YB+gFJSlAo0ZNmtCrMy/
iKg2CNzprc2k9Ot2qzQriK3JvKbJBLPMLcvzG1/VNKSzZLpHHFM1EsMH9+X7tzhr
dG250SwHF7WpuKM+N5iaguMNZD+JWivImUUGkM0oaBaejpylkqDZshdl9ijkLuCS
R1Yj/Hbgdb/AmcGRUHImZKD/1s1Zx037+9LsYS3ABbvxka9HiKg17m+Ss9hPVsgT
XWq+R9lD9XpqiFSZsFtgfasLxacIu3jl7GxEJZic3PfoNK1Hr40eP3PH7JjOvB75
HLH385T7VuZrpWJJGgGg6kWiBcRDNSwxCLdedieyuaK2VkWloaVhpk3UclhW8TJW
CJgsGWOa1rQdjjHVBZOT1VaB9zGOc1kTERDtQH8vQhopAE+oZSLcRUfKhWQGdJWN
mRhsRe3NzsxPsrSUZCQX77qEFQDYrZ6DdB4DWcaPFkh54ypHpKxabhpLfSvd4U40
AKWIT7CJGgmNH0mXD0+SPJevdcqh+F2YL8NXa68PwCvn/fHG8tn6YU2W6zDtkYGI
5qHu97YU/1hUXr0a3CSRuBWS+FixZJXXzgEnutlzC/iozmwg1bODFKvZYqCppyoR
wgzHQXhOzhH9+klAkaKXEVHTwEMWv28rkVceBgd2E79sNr3evHWXNZopzvvO8Fzj
ZwyMtAV9Yc5d1uiBnQgHNrohubPrlSVQF2Ab7dZA6Fr2y9UIrQ9xGcQ1vUe/D15/
BmL2fABFkzjMBQzp4PPN5nn6uc58o69iCZwZZnM3p9GdKXIkx+V+4sq3TBvBRNxR
cZdpcY2xM4v8oD2gz/fDhtDa/qjgV0o9lEHcu9zx4vcJc8db07yTrRs1hGQgt9M2
xJrkm7YwM343cRErsBK7uYz5XPeNyYKX7sh3j0GDrzgQq0I+VoJR6eESGFyfBBBU
RjPqFQ45O5oMOUJj2WpwzYzLRcdpONJYTF5sceEwHJSIqHyaDJY2CsVNrXM8s5t9
XcX1HY6GVHbVTemVlKqdPtV5+YTZcXr3Z4tzpYCwjQfBf7m2cbhoPJDW16YVoUdZ
cmGnuATdn++oDJ8hlg0EaY+sNvyIyRKrhb4eZkUmckzYuBi6cyDV/q9pnkmgDMl8
//bjSzMr90cEgEy3AgMAbUkhGcFMSgNxft8h/JwVsPS40hXKr6RpCs3waS5C63tN
WWdilflxVLVkR8M/l98+p6PcooVSiwuHjKJdz3/Ax23G36KRhecf59ouNfFF+DCk
zmkqdFHuBgQMT5csutxwShjn9GHHHRPowTeYD4GQ1zi9rdl5SEa67g6J0dEvlZV0
lmbee77hbuuCSQ88faqa0rA/ti/uF+pWjwKZYYsiE43MKm2TxVJK8rjNcP1ggDLC
qq3Rh92VA9bujfWDVquxNhmyIwV74W+R1V+YDselKwbCB+EEDY7/srWSz6RVqE2W
rTwu8qWkwZ/PoF03ZIx4lTeT2pZZUp9r1AMA0dGMaUAhdoZQot76COWd7RdbOSe7
PpyrGDAtyzjuo1FDz0r0/h9D6/Arpot9A+WPMnWYxkaJjInazcEgoK9B0iJI/Oce
kbdE/FMCd8q+/dnRQwQdLw39a4SJcr1axpHaFZCd/LwUu4UxnxDstB9gVVi7MnwM
fLyvIrq8kCprtRzDnyCaFaYYm0bn8ORTLUnv51zjUVplCCGKDr89BCaQx00gr00E
0VPftUhWTL3bkt9FEVz8RmA7KJpDqAiVwi4uQbNLUXw6LqJcEntxzz2YhGbjeX2t
CMPlnYW8mSQUilRYPwfwZqjlY1BafTrxH2bR6o5TiQFKzm+AcuuDtsRN96vaGhbH
SYFuqnnS8cI6y7vGH/UbjJ33ObfIsYRv5IDP4bxcektAD5zIdgPymJ5GSe+Bj7ry
RiY4DjfYMBAJF3WD2Ns2wdRsJODXseOd41QXSlEoH7nuyEDNJBngRBPnfWMKMkjE
CkUdJh1ks0v0Mbf/IMT4k11uBfzSew03xzNxi/UWywrnUVAcSxx94LSzi0TEuAnq
u5XKakl/0INjBXrzdMdIY4jOIzASSCIvFLiwdSz6tGD+e0AbLFYPFXhCdp9q/3VP
xXAiotyNvjGDPb8IFNZ2KXsLmVOM7T6A7esu6aXMxm7vxdX73x+95VNVlXHy9IUE
CwLrRnMcrRVFyXjwFUloqycd9kTMzYhzVgnP+7gC2SerhyPlPaeMFwxXILMGcgKm
zwK3voLLyjz17bPLTMzWQ6iMHS0LMcDK4+t4tbQXn2xRt3ArHJAwSPZRGo7bjoI0
QRsFGSZGB79EzbAasWCb9tBb5lmeh5OfW+zQ9b1jusR3iN7I+2B7WXLbCjqIlXPB
YIC4j07sWTILEyzPWrWbrw+qcGzPTJ9H/uJoAvJmEgmSlwSQ9uxAuQ6JcRXTdjsI
T2Oz5gP6bb6odxkRk/LBjWrwF/aw01jwNGF7EvNAR5XZ1cnmFqu3yL3fqwt4bSfe
wLoR1EE6nkj1JN+uKKrYw6mp+qlhUOrvCizG1UZelFAJDDpNP021eL6y9uMf2l2s
nGN1mjL8Q0aLexq3whuYhQpbXQfFqnCDsLVA5b+6jBNY5/BwADK5z60TtsuA6AXi
OKhqMTrJQcXXkEA53FYxXb/9ogErVAtty3Ks3t0R6IWriWz37e47VEyA+uJoV07F
aTLxbXfubtFOeM5QakbM+60lXPSISQbjYY+wIj2/f7O9elkf1FBo+EpMmu1gRbGc
FRqok7Z2iKQNMnkbTMulEaw0kVOr2ZjCwM1eczywVkonzKZUrHBlYOwgkm1HTBIS
Ac3Q/eOXJ/TLbOiYkk6dBSVQdNLwKjJwkAKsodov8BVfnZiXFY0wqUJEHmlgr9u2
EHxvHO28NTWlh5xHs7rW3TSpALVflZpmBqZNzjX2rAwmuqJs+5Oky8JtC8qx9thH
nAhniOp3rbAH3awAvc7atXE8LtjcHL+v1jNcIBeMBKuP65dX7HFJtb9kh+3LfsE+
oO9GF2lnXFgvKV+XQWw3mUfAuUnj0q3eNsAh6+/acYNWHyigWFBaaBOctheaJcu9
TvlkH/w12MyB6ciQ7aUQ/2OVemLzdzfMkliI71xetKmdiaLbB1AHFcaiG5H02fuU
wkFiNeTA5Ak7Aps/WBAt7qwVStAaZpn7PBQn1eoIzeU48ztSFKaP0Bky/+A9mwRv
dO8Q3ggX9b1PyE16Qc/K6X5X9ocj2lGEKU8oIk6Z6Y/YJM8gGakqxLXwDKhBLBCD
Nq7913bO1GrLEFEkrPvv1ZVAME/7K0w14Rsn3gsksCamQY2C/t+cr37WPMhvkncE
fcLzIzMllWvRICStW6Z1CmUeVqfwHY2VM8RMaRlgyLmRQ0Ar+OS1cNwJgVSamESo
vT1QKY3M3TJE50t/3GcGfK61o3JlbDuTjiYVCJIJjiHhjdI4EAt/13MJ+Nwhh7DG
0DsEZNRFbbEonrNL/hbN3eLD0Tnjug9CwqbTPTqfbRcI/fSlRQ7tvQVDadKS29e2
7PzVL5/Y4/i0DHjDf01LAM84N1NRNLI5Dqo1zds9AXdTx/ZHkFZLzh+ax0Q6aWVB
ApotK/UfbF6rcXPNJcDWrLigT+HXq8t0kVaXp6dye3TzLTv3XfgBT6M1HO9gsRpJ
mMimDGGRwbj4i+GLuJ9ylE8I/Pdwd0KCLJKLKAHQwoLB1vtfZ3+B5+FSmUIRx1vy
gaRalLUk2zNN7w/H5xPZqrO4kP9dz7ao1nTV9CC7fw0dK3ow5G0mAslkCS9WfVgF
J/DI5HF+P7eIJsIm34cFoHdMXIqJavUDlECnRYyAhTsnEdHrO8gxD/susntlnu+L
sF/Wj2dahuSATSZ7Kdp7fGRcWnhzjS7Dw2/6tnN2e4RWCysY9DXQ3SvshzNYD64f
w15+D7NkrwZ3IoGxZwae49AfVFoWo9OXblazDQ6u0i0oFuj2bk6tadcVzzuBEMbH
jhybAbMho54tgpo6VGjjdbOLAF2D3Hug2pMgX3yci+msI9qmHsZjbdH5gbgzWNa5
3XvDY2zjxr0CIIDs1nL7fdOmCDUQTHm/yaa40QIG1gbjZuV3O93YrbqWC98vZlNU
2TxqMkoMVuNs2VSFjxHm0fdjhxuum0nu1xuOjbrXEoQy/x8ajGnQEtRE6lWgdFsk
3e3kfTsqeEazjJaGNbE2lC1aAFSFrUnw5J1WMC5PBQnxNSV9VKU5YVI7RHYfQw0j
qqFIZTvSiixaeI2GZ1q3G2OOLluGtG0N2Z9cHNvxAboCh17Kh29Me+baKjyGTAHK
fWWEP/2zgSf8/tfd6V6mQ46L4G03GgNyCRAAfFHoEXky9G5b3NZM+vqVEFsTtrsP
5DFAKnt4t6pHr1UIn+Dfut5dtb/dqocCTQ1ZTfDxJCb8H6taVyxa3Gnvsj30Okjx
hRKg4rZQQ7XM8j0lPQcVMDszjUtjXtGCHQ0Vxle0gPoL2n18EPA06RIp0yew54RT
3Xes9ah+8yHs92HXAEJZZVrWtVjiv1cWyeOfWsQzw6ZC9OTS1uY0lULnVuWwWRXr
E+yrgJD0qDX8f2H6roZPWaUXsTGFkWoLQ1bGH5ZLjCp7UPa9gZMn+I95Mtrl4bAx
gSg+JaFHWE0H1GJ8IXiZKnSoNCz+1sqJ+XcxZhhGvlY5xp1guiaN1yx+fsdmjAdF
9cOqUmrmcN718uRePR9x8yOdyl7KnjbYO6a6JBwmhWJBccR91DgqneSZrCpKx4lC
PutDcZlsUXRIqeDBGBgHOZhjvg5XGq9s1X/sNSWh7J9Ssrs77M/lyrNTR9IBnTHi
PFfJ64DhGKSiDJGzkFaLfPmDvuTI/rDn/R9M7+c0jVVMqHgywkYmxhfRqzOMObq1
AaTuZ8kaDga2FsPe7pihcCi4cFhrM6UGKPoO326nKbgqQ7nX2YxcPNMX4w9xdqm1
TMgEafthE1cetKbcxNBp5hqmyYcTiWlZu5FemIusCZOZrGEJd2ME5NgJssi2eW1s
ABWckkwE7/XjVGSO2gp8mglD1jXxN96Cf/lslv3T4mAIyZdIyY61kxLyrzQrD87X
zowSe0dKJ58/ohKhsKI88VBurm48aHvoxYxPtHwZ7Z2Pw1CAZsVm2XfWLA6JeEkE
YSao4AdluDxmJpIeX3oncXR9oV0sASIle+SA0HxdO7yP77rD9ocMqKChaYCtkiJv
4FbMpXH7ne0stXyEFifTNrc/On1itKKSFaQbMDRWfkFspIvuD7pDla+YlFGYcCuq
59L4sXIaKKc02XGaLbD0A38RqnY9K0moG9yptTLL0PJxK84SSwQSIJcdZxP06tqu
NvW9ze7/9lRzvDM2mTjqgoRH1Q2871n8zaGFYpeAhB8LSoXhUQ5Ix4DncUhOjue2
KRHAwOi/jrOz1hqLA0JNDPoGNSb1XTsEDHBo3ZxdxzUoCkpepxVP9WGPcGAiuNQX
xHO9u3SQYHRYX+vBFrlFaG8YPTbgTE+yBH16Ym6Bl6mbShZqU+0nIUDuJAbvx3jz
qV5R0p+Y6wiStvYUjaacK31XvcAdoPmtekP7W2rDYvap/KtDOeHOf8CGaL4gDlj5
QcZ04+Cz2Ab80EsOP++LYz6r9iau4BGK8GQ5+qXj3uIvlP37T66kreGgO9+2gMtI
BWpYl0qD3gdET+HEyiYMnqVkwEUvrdabFa9vslWpDwOIk6vhq5GUxBvKtBHznNh0
mDYOSeSUkUEwW8R8aGpkPbVhn9uGnP27p5VSKKceD9gJEdKj6hLWRHgE5vvQRwHh
aqDWDwkouAHha8YF9nLF8b/i2yTKlKDV9IJF2nORJGQdLyCorso/r7LphDtzjB9V
jQNkNXKaq9HKgdKkRvT0VoJNuKq2uPl0gr/jn+S+T5K6dp2wzUnDVJq+Ubwbk/0Q
5w5qajsOp/KgQEpLvquVMrNskv2A4GslGZu2hvi4N5xCdvTfJGvycg3S/Z+aoCik
EsIi253zjTbMNknAYIXH286fGF+Wd6K3QYiRkfNELujXJWC//GsLUR7V7cuW01K3
ccnyT8nQDYxk3C6akecNoalhIODZqnFssmMG07K4fnYYNyv3N9js1SLXitteYD4I
FJ/QupoIx37jK9qlCxjPyq8e38qi/h6q+F4Q8AMT+IhFwwz0AxNpv/hUehjPhH7e
MoacDAQfqzlffMqbNinQU/Zzj2ivaEKVg4U1MRgRuoZ1h3IxKUfQbAw8f0MWahwY
993Fnd2zt/Q8vp0oamNHLJFz21sQx/z0KYl9myqix7S7Dam3qd3Jl/U4KaOAQYw0
rBGisFGfntqUo4Sbt22zd1jFSmW4XWGOc4iHOOoWwN+0/djrd2D1bjbT3AiF2NE0
XN4Za4VyeJ3AUzkUP5OlYLGSmRlDkVWe58xZX7I81gUhkmgia0vykDylVe8Ja0a9
NHrBxGuIUrCbitR5JzTDjvImwlv4i3yCQyTwwDU0UeSU6bpOjm1BncbW4JrFJOHN
DXR1Iz1eJv8lygRNy3cobrwZjGRq1EvbZq1YMr6dNBla2ixU74dfmpW9pQuGeSvA
6uVU5sfv/lOG1XPPvyT4+YcBMqrwD+x7cXkw/eVKyREMdVRpfgI45aWJUGm2QXvc
j3RM7dsmrm+e6jupQJIdOJF1i1/N8hcT43BV4nWnxxSO8O5ajKlSlPKNQPBVszJL
lmhCb8mSD5W3S1CFWX8vRnAxr5M8BqBeJuVbP0o+9F3dNCjLoXBDpC5FS3weLwPD
fzc2nwK3PMCcLXIJQ3g0bjIRJT4G5tLvfhwC8iJuD8j5HgvmIiI/m3jWfunEuBO8
zm0EEZ4VjQgXHrALSe1rRrJGgsuUSRodVZJR56X+tJHdrgNfnrmikTL9LvlDIcCp
GV99MePeYZNSN88jjI5BxZqsycbFbRmL+qCKF91yjqLKMlnmgAyEGTPpcqKJBagU
H4RUk2JYrDSIymJVDACL8tN0c1hAqg7SyWgSNDfewqNj/5aPfptictMnpf2dt8Dd
NJxVIRT4CzQo15kfAGkuN0EAfiEJculUnx5bGb1Bb9AhrD299kVG0nafXe2YE1a/
3qH6o7UwXGa/JuFVazhkmfvAPdmtihhh2E1/jb2AJvkiFPeLWt2jIAVTZiiz/UKY
l3Ri68C8JNIiQD+K2H4qXlnlx9fQCEwGg2dl7WQo2qoZOdS179UwaqJAPul/2lqd
Q6Fb6IASQQZQZL29Q/Gb3JOMtd/KN8i+0lMw/CCZpcJdjBLmo/6CWEEWkx7bBugc
+Z5oipoXtlCg7auu8vIQZiXEYk2dNzDxwD5TW4yl8ybtWhkARPfpzzulooZYmzaC
vkLl/N6vxnG+JFvf/SGKgrgtjpqApoGjT+ianaI18h5biZK00vfprxDOa3JM0BHE
CmEpUd81Nlq9Bn9eq6O8EX3+yCo++AC6QSc1z7j8XybEXWSXXvZ3lvGa6fBZssLe
GYsjVOS8iyc6uNDXm1QeC35f2tCM8UmWDZHSRZOv4jg246ZIj6GiHa41gE4acuMz
jFGgLYWdwKJq3DODOfsy6i8wvqejlQNaMm10fHScH1b/bHLLIv7NCDdGt6La9aSQ
ZwQnegL+GeI2VLIfB2/kyb1ZQV3PWMwYK1TXnLChW0Mkt//ZwEcxmN8n5qc5weZy
M/TKHu9H160mgXYx8Ch8QkQ0XlBYZY/BK/+6db16US4Slll4wliy3Ssp9euozTTl
dnlfeRGegulw9Bi8J1q6VYnKgC6hv8/Aq+BChQ4wLid2IH0p1TffOLL/vz4OvAsF
B4h9c3DbypG3iC4VzLyLmVA6gG06wXMqCbz9uMT7T/R2c76SMxiKrdEoLORUhwit
drZQ+Pp9A6kp1A7FBEnb/jYYQmIqiFIbmFdr+VBqdgb/QLqU9ldrj1Qf3HT6kX5N
F0I7cLkrLJYkWkxPB/VYCTRgCDdVKWKF2oyeBmsTvN+K2ZOpxSoLeAJpMi2V9Qcn
YIOBi1c49ORFR6fy0L8RXsqFui5KJfwZ+IX7QIVxDmmLdVhEl/6nVTXF6CIkEZcA
GEHRuFZRpsJF2UxWKxm+ICx3VN4/Jqx8iCvsLWzNX/ERl/Qr5zBASnkdEkrEI6rI
gsnXAiqg0k0I6tjfKvNFE3+l2bsxIDmToOH37T9+AIZ/zOLedBVOMEP4Ucu+p9F+
l16PYKniItUtA0yV+bhltJbzF3H11lx/HMSC8vDfJbUaliJMQS4eShCb7BZZteH9
oOza03GmU3kCmbWP4PY9jQXZU9Cis1i8FFrpwEco/ukzineLkfv4DyucGPyievCM
vn04lfdHI8m1b7boxo7QbqWS68ue5V47Weq9O3VVhclt5Ckokj7yv9bAtla1uhc3
+sQOhIPzr3vAEoD7YFvDRTZNMprMRGgmT4/AHVK5cYAzdDP6S4bH4qtpNKV/C6Z3
QDenCgtyRf+gqUx09BmTyTNsWwN8EnYAoGZvdjfdIPf8St+h1TJ/YZSP6iKvt5Hw
oOtIw0XeSLmqtOrkVcjP+fnUDKjIaeXPnAnGsGa4TjzvEFYBdYE1L0xcuIwvIfjS
LVKyPHixepMaD6adrXFPKAa8TIlGBy/eMpJOlTYOMPaJW9MqjVRzZJBFZhRicY8x
P9q8MbvGCR+0Xtg/swu3BlNM1Gvr3FGkpg4XYrvscGEIPcmdPwmrrald1JLUQ3os
Cz6Kx3Z/839fjIQZVI/2NSKJS/MLgrh3+eqZw8w6G1fE1AirmsvOfA5xmJFT3U0T
6qOxNy5vhWIFAyoG0oNJOMROhfxHwzDwNXiriV2QEQ8F0SGxGikf76+n4EcxYRAJ
h9uOV9vFLZDghUbqNtcwXeUsP45rD6Ged7XVXWpVZcWAgCp51Gt8fmGf9kqh4dci
rUdzgrKUfcVtNKXBrM16F8LaJRD+Q5eGADmgeYmFKcG8Zzga2PW7BvPcKWJqo+ST
YAdpCjPjtffAx/zgJ9de6x/UnsHUuKWppupvnaaQfuVTxINH0t9w2Ym9P/HPEcia
M/qwFhc7HtrCHHt7MsRcZ1BD2sQHk8R7WN3iRxr7mW+fhoFT2Rs5yXlYgccvDPIU
y4UjYSco3LeZV7mKEfmBWGnnFGVvof52Hd9DF4n29FSjH6FOA/KWOIHLkPF5QxBc
goWkHQ2TIIDdaR4CLe5pOAmI6iqedrOVIMc5/k/yZ4vbOy+IxjbiQXxwpvooFBvO
2PEA4Qo6hVktRRqMLa4Jl4TImqQKB0B2VxSfRt9ZfX/UpDTcJXvqRvddKtOoGh43
IErPsI1Dmctvvs9ciutxEPb8GNRAqSvuCot3tCnMDkzsyYATxN3rV2uLb3vYgyss
M9zIf5kB/+Qb3fGO3XN+6KlCDnaDgX29IhvIn6REzxyDDoeK3iOIYb9qoC05Y0lJ
baaRYkkFzdyTe8polrs6g0IIzexDNk0klNUIK9Jvhhk5QqksVZmFqOVu1RKz4Ve1
X9cWqcVlN4Kht3kd/pgjPbcGZbczuT2QVCB31fOkoXDhQeoYtvCPBA+WhAInrQ9o
NcwZryvaeO6DKN2NL4B2rRmQv/15z/hyNmI9kpihl5vvBlXtHIWehP8g2d+yEfSN
4ezueVqdEdAm9kOy8QS6CSD6+dnSZPHNl2J26CWuj+xFsuz8rrCuNhU1HlKLy7y9
t3QDUXmvP8y9EVEskmwxMfoYSR5Cn9WoSQMhawFs/6+JC56qilsYDVbNz/NGdYLo
sxglCDRZSiULAdm+J34QcxrPBKRrlvBzB71chri+ChsR7BZbhT9SJ4Z3OfgATm0M
vtJJXe+EKt3JFuVtHUYT5kgQHZjUDhOP4G7VOfmwBHsrlJGDGX+NuTs5sahGiLNd
9Y+E/WhesEMUhqKRT6odd1B4fvQhq/ejSZncmTSwmuwkab9WER23OO2jHNfQmN9h
nORMBixaana6jGjSQ6EUM44TVTluOuT5g58yjh+uHu6gnWeFLXJbfJto0zBTmdM0
2BClJhkGUFObwFrhb7j/+FRF2MNFE/T0MJDt+jdcUNYGF98SYqVy2fW5/NyD7rv8
FiBVH7Gk8U7E5jjMNqIX305+peEJsoRQHHNwbF292balVDmtaQDHNgAARLiDBd63
Lc7MIlUKi9y/ox+/cO52gr08Iu+BfqgDlPmRFtDQC4eEm65vVjX8oa8gljOoSIqe
Y0iCAazplgEbUoaW3tUWMuQouRzXlgyj/+Aguj7i+zBL954xAb22CkQal4RqQS1/
l4GqI3tTkAmEsiV4sWpjX/0a1/Hahptc7OB79l5/xcAXfWv0TuyxzdT8JQ6rzGHX
ufakZxLE5FJv4eMu+PvL50JlvueM9J+qc3CinjuObHsLHhMzBIHffRO/iwWsjqlp
ugM+g3iT9yETPgzqbn+R3bxZ74yePExoFUFYJqo7e1DP5J9f7+u51h7mbTGXdPcU
vkJLloKQkLKJuJROct+wAu33Yomir0VpISSHPlswx3kX2SnF9HptLqV85w+lv3G2
4pnOZKDshZO5Hv2xyxyxZGLYEZmZCN3Kt25gNFoh1+zLfZ6cdQ807afEbINK+eZ4
Ums/d5NL7vPsCkrDEgcquVeVwJEoaf19Afp5jYQrKniO9ldj6IqsI00Lsxou9yNd
UFgSlBICqtWFLRBownwd9/V6/m2uu6FRB5MzlWDcimu+uqTetNvVBiSUheUPZaGA
DiX7Hw1etgKxi0zsiJVhG7MYS+EMNEZK1R3fF87zYYm+v9FS95LJPjcyAILUeXnT
QQWzoGBvd+//dnKSaw2+M+5OjhnBPIsgrWk7mx2aCHKDAD9P1EH+xqwW55qUT76I
YuO4n2xS+jy/VAoGpLkkFlQl3aakpBMicVsC/DaFyewt21NPS3F61cWQ8+3OmZjD
vJw0j0L8hiKEgKDxTpoI6Wxz27te3XY2sOyM+G4FjB76Pl6oLb9J39dGt8I+KDUv
dF/28z3B2Uy0hra7WLtthqfvlH9BGeqnYivx0IvKyzS3WL7Poa1oNK7KZILOnOjP
SkaS8u8FiiYVOAyi5D5RF0xCgkMNLoMy7sFEMklmLtOPqlowInkjNX/U0tWOwSzG
jTCGUgc8zn1V63QZQwS7EVnY3Q77xzGn+keFretgTEuk81O6ELpaml43CLLMr41E
kIIu7T+Pb1KxD5xqeytUVadO0my57uAMvUIDMKWv//K/7zDNepFwSJ7vagsRDb1r
vfn4n//xG0iHlzg4l0rSrzvZ3DttqVjevXG/RD2LpPuthwlMzHBO5xLHlXjWLqSa
5ydV1Ca0BjWvc9uR0ldfRGyg4i2xVykltnqfc8NREPQSI+umH350Wy8g8DHvvs29
nSuhchgsFSxYy7UCN2ounRiSoNZnNcJUt5lnZiB55zmcUi4hI01oTE8FnT2Uoc65
OmvgvLB3772ooFrHQbZcqG+j0KJB/8MrsaFvJbUxfQ1V36t2X8UhHq4XgVyetll+
dmfFSu11a85LfCKYdp36KSYG6JKvEQ71wsTMXvs9Gn2J+1g8EpK1WRNbSMd/8VAZ
4GyRDBoU99Qw1kjS/Xx9rDEfshiusA+Cr0AC1qiZoBbkS3LO68+hWNEHhnnf94JS
3WvZRLryjDnQAYn4AjPrw7lq5bKmCm7EwFMRZcLn9wQ5w6fkyyY11G9kTqNfGMdI
KSW1qsee3l2HWSmxJ8ZfEExYvwBjL0apKsBzl/BikBonXYLmKu2LcSvLyrhetC+n
mtEYYy6OcCtcNlqktsOX+MjbBEYJnt44z6TVHHUeMyNek2fVPWIafJa3LmZM792s
Dacf97s5TKwctCgB6ljZMWtFHjNCWBwbgFc0CBykJ/oRVNpGlIPRJUm9DB7+lx2i
4kRkleYEs1SgQlAZDC+Pe6XCWMeS7odK+ub8PdpnPJ+K/N1imESbUv4F5PhM5IDd
RiW+b0KxlLt8qqHatoT8ZCONhyOmPYeXYLhOEZqiGaQbKNzILhbJKyRXb/llRRpD
iVR4Yqz6Hh2noPJw7FL93v4TrTmHWtMwDAgbE7YfkFoJdLGgRKgbNiShMndeh0Et
VDdheQBuzO9OVIT4xHkydnILK47Vnr4Q6nLLdbDCuao5Dr59qhIsE7I87o+yX1QD
Kdq8ZvO4YSvDjyRIYOETIAoE6k7kkpAYyKZyxHb6PHt+Et2TstfQQyRoJrNfeONP
Ei7pJ4ra14DQULnvG7gJMih4RqUu/dakYer08QFAHdNRSsuGy3LRpsdlR3P0QH6B
ffYZ/152FpCfSwtDF4cQHTcqkUcoLKfpCEITirVINlJwzEjSTeAo/Zfpm2vNq3My
+5IZLpEJ79mCwWBnQ5ScNhjc4n0SMi4bMU/QHjlVdVa1qk8BkSutCzyLJbM2cdKv
Z0Wog0gwGc6OvbhQYIy0HzWGRpzwMRxhzILxHimZrUtUlczNyTtvSyXpE/e68MQ3
GcyGWoXGDRLnyscLyUIDOkphjlQvqs8anSx2uMTf41LB4g+mIDysOdQVwiaUH+sV
uxBayAN1fMBsxZrVqCKIO1PGeR5cu+r7dJzsuZq2O7TofkR+FHHy3ENA8mJ3VF9y
D4P6MYkD/VawKeBclSpxYaR+dYa4pW1pWKf3ZR18LY73l2TEPrvQ1LLXeWmqp850
1kx0KSrEVBnbipvm4Q7MbJOZOLWd2n9ZuVl67z0FMJ5vFQj8hk2qLKyQLNcl4dq8
kT0vhr5459O46XTRCCPKiUCQbDOdHwL9Lx6si9vfH884Pl2yYjBCyN0Z4FjCXyp3
2CTbRhnb9UTS9KJGfnoy3G1N0I9klVeBFCFfGssswWm9wrLaQSVQhGXCWRt+EO15
d0OJ9u3L6ZkC+cNrXfcwi43llU3ZIG6rFwTufNh+DcH++HCJ8/ekAC4Un9an9LzN
tV3R8Um6Nq4jNwVRasVYOMtvGqO8Q0Kcs5s0p57CHInk42UQ8hmvDGv3D4I5kHwm
qi4KD9LNX+jcC4jaVkybnb5HoCSgr0W9Ar3eGDXPePdyPVIGOxd1HjzaGk3LWt5B
NNU/r65OmRwYvhJCPK2r3Ejfuy++L+w72OzfzwOiFG5/9XXEDl06mHa7Fth3dp+I
aR6L+w32fR3Czobgynf26l+RzyM01JIYzDKq0untvabBOXwM2Bjz7P9xLUoXLPT2
+b2u7THpMbbNBHl4hreDp2i63P5BIZ7NAan2QqLvbvHQDSJkuIf3qaBu1JRTLAo2
9MDeBcKzT0Y2a0G2IbMkdRlkofybapwzgJpiG5titEDoatW7xrUBtiQhXxYMNlcu
0SF9KlX4S7kN8gEVc8hKbx6tDjM1Ueb3nZr/gXa5ayYQU97Z4PatH53OndtbclKS
xVWLIYcpx4kEiK5PYQ8/0mr5vp5ZIqJNgcVfkFEEAkRItLXNR/b4R8K/AjWYannx
RLL7MFQ1lL70NJxB+zhACtf58coV3qB8SSQ59Q/S3On1uzM5M7ReZT1jwpEpf9EX
URXULO5n+sw8taoGVnEHGGnWTItijd71eWrgkqttOByA2i6k2Q3TBnSk/mtP29/A
Y4gG/Mf8H+ecO6i5oG3yi4v29PecB9uDboJIgRKXMAv6TgCAY9Pg2UEB9n9YZQnQ
kt94NQPp+MSMuyvYTNqGVhtqyTijfVrblGq82hG7xLjRBDproDymL/X/sY9g6iUu
4DN2pJBALMyRMrMx9S6IdSysevRLJczGIo7sO1BYF53i2WZwyUhdbnX4V0U2IsyF
d4M7Zj0Pwk7tdOcZkrPHrr9yS3V4kEDowM3y7ETOh1ieu2dv9EWn1zsFH7RDiXdh
/WsEkdjWIs0Pod1SYhruNOI6dSn40UEUtFyHJU2FKPqRcMvi4pEVPAzF13ZOzVlw
o156MaTAlQ3VslO/56DLRkN4zQnyjTOQC0ApjtpudhcYTOG3l4xopsCjetDg9jVR
kYxqZxFw4BT+SWKptuTnl8u50PmOu6dtBL4yuFDHy4Qe4xx+jXOLIB5eOtsKhq3K
7YZmgW49ggjge9nCmI9xooXUoJ3QTvcjvVC29YIqrsi8M7AUY1JnuYZz2ytWbXU2
RyUgMQLc86oZjYgyDzMZStzHUK9Jb34FcWSYugBHCCrsJyQSuQx/WWrAchijYYeK
MLTjKMzDt5zPFpA85HoQ4wllw0Hq0i9nssMgH5Hxx3BLNy5GCWbF8aNXhoHksIBV
z1Ly36pvz2StldVlrMecUOhrY6TXbx1SE19UbYmikQ2Bm3yMiRCzKSBgREswh/43
EAdg1VvlRadaiD8USTrLYH/ugeAsJNWfCJi7c4nlUUEJomQkKSPfbzJPet1k3vXt
yvD5hYMklaBiaFk929GRTvsXhL/Dg2m2DdAfLqj8W8W43lgHgZFRxpATHbk7tnm0
yWGHGB+PGp2zmHkl38BPHviGurHf5YWuCV8+aSiofaCT7XcZNMaMC/Iilf7Fwzg5
0iXR+Uv81ud5kjYfg434QfiPrdTxkiyBFFSTUVpNf5YyDupx93xeubiYQa2LeXNj
65pHgngpTJnfT1yy2po5wkOGE2vnE5Qtt0J2vBZls/Aa1viHyyXfm+jrGqHlNaLX
O/AqChBgv1i0stHXW3YL8IukJ5MHwY8/+qYqgncBRNScgpj2nVxtOGhBj0KZqzsj
/NBgv1FFB12jnxO5aQlt1G6tN2Wc3ME4bfouIdoKTn6yy+1hTj4e7QCgX0hlHSpa
hZ7dA/YC2z0MMtsVMzQXU+lYpqHJCV0Dqx0W8ido+4EKa44QBNuHX9Dgzav/7HUu
o2X0nlqh46SvMbnmoE85H8kYP3rV3ReQlgyVdpaZ3n7P6DFyUCv6Y2gEkA6s4FQo
fPYVrZaR6aYOAiAOZAuSjRuSkkevWXmbh/DsGyxEyHaxnetxg4bORwizIUMGX18y
O2+Sv7TvuFjs4wxrgkHsgGqt2SSkwHQMpNDQCbcVbwZDtQ5ZlxXthXcbnYhkY0sY
gJXPnyVejBesLJ5zDu9r/gccnuQDHYJ22IWWind8B41EpEjt7RxwZBXVOQDt+DV6
zSS3/5r5z8ahKdCOwl/0e+dn7f0VThiG2OvwYoH8MOEJEAwjM4ihAyj5YiF0nNFW
Ov4A4cpUeDVdMFAs4Nxn/HKQEDoA9tZSzK0fudx/KkJaWqJECw/jxZO5+UJ/Ehd9
Q6U67fwcE52CPWs6cC840H9rRtP28GlTIhUue1abKE/4HJ468W+qOF2IS97UOLn2
PWckR0N+kC6zDcv7yIvmilu3fB7C2xEN8kWjQGs14hDnxezE+ytwy03KsWTvrEJk
V9RoQKB5JwAXtrtb0wqYqZtYNVfjoCVPzIz7dyIkSKsDKG+7faVDMLrTy3n4rHxt
/2IsUhlBm6L54crX0V16wtC3fEM7A2zMLJd3qQJF2aV4GGkeu1kG0t2CoH1LL9ga
smM7hO1H+OGb5mP2HbFBAV4BzMxPkw1RfU1M6/bKIaaYIZkq02mEN7pzpQYhYkU1
s/e98rKt2+AnMq6KsL38EYfWHeFQfiEN0okcBj/7LcjWgJIzJ760XIQwZZhHDP00
pRaaot0tE4YS/BZPvzp+tcICFcwpUoaENOb9iam/cGfPTrhPIBURlrOgjVVMRfP3
eoeLM3xWio4Vi42Gb7bfgNY7X9xOgFQO9xUxqWAbpseGKUnbxNQx/jmWV8o+wE4S
Hitf/+kzv3NdSJyyjDYucObBnNx317Y6Xl/QxExFzynnMvSgym0eonE6loptagRE
gBJ4zKzhS7+miU54B/+P8zDx3hj2xubNJUeFZN0PdEqPT4bDu8P1XcZuIwUiIFra
+1Vqtwhtkvjed0YkFOfH4/KYuOM7tCo1L9PuCSwyEEJ5IHOWTg82X1GoEflMiKfP
MZXlitG44lGYg6edvH+WRVs/mmrRhCZk8zuJW+/md9KkMnQvknQuhkm1badcHt3l
iHNxtN1CydYscMZ0SOtstq0aex72xAKrKQfL3e5hBXUDONi5sMSWK2KNTfjs2Eo+
YCbJ8dBVcaTgVrNifx6+fKq9nKF9ORueN+Ly9fxTeKXnHbHPxEZ05z2V6WpA/h0B
qw/6oN/6v56zowkx3nFB5n+r3BLWBM316aXTwznMM6Mu9Zh0DUVyu/LaaHpmFHui
FNQB93ikpO1LiFUpRTI47efp907pzG9xP8/Xgv97PWAwRyfhD7ZFj09ovcPX0/Rs
mp1vaSGYobmSrTY159veXiDGim3GKQlHIgwQjHFoV/6HWJewW1g0bmhRJrKtxrl1
MWPcqx1lxkJpkbzyaRFEtZ36E1cvrySy2Lfp4zX3i0r75f2fnYrpyusu8fwoGFWc
QTMJCw9DPJhrrb9beJvg/idIOI+jokPl1MHKkutcDZHx+mxutJgFRVWY1iuq2cF7
YlpShVeoaNZ7+4UZCUkUoVsDP6ws08haFl6q5KzJcxYy8FQQoymrG5jYUSjE5ej6
U0Lv0YH/pmAFJvAjERfa2aFHMBPZCqJ1cNEyHiEpBSrybXmpSfldCSYc+mWoP5sF
GjVd8BVeRSritgvO5XOtbT5+FwUd5ISh4MGFpBqJj1gzKVr+swCRkmI5UhfRkQw7
3dBcw5sRhhbvj5gotm4cV6mvoYNNTvplgliXPnaDrtvIiJgrIbQsi70Kqii2QCrJ
WzgJVkNfAvxUhOoaYYlhGJRtd9z857ZtsM/JbVUMaUaB0X7YB7oLoGyUTyEHjrYJ
AU408fb5rXcZtY3wUoK8uVRf13ll9dlQyAi9xDSLFpIoyxNhjyxsnIKdr5h2rmcQ
Ud0MOi3dRod1JIG7s/jPWHDeUaZqHQmF5sohVEj+O/AdheKn+FbbMyGfbfX30mm8
FNRXrWvDbFCPqs40N95RnebbiPrIgFHaSZ8KXCesPSjFFju3bIkjhlx4iCWDRMYI
q1Fj1JnwMI4xANcJgLJwRMMMvAmxZz88VSQggY7uxx6MqIPEOLRrGz0gi4n8XwWJ
miJ8Pviup1Y5HzVs5FSE8RXhxKx7fHryzE5l8gb8i+yWHz2YdXjINJxABxjMYqey
RJi/NuB0lgXrdplKD3iQF/c3vb3YFHXgjVwwTrQjQ8BFXllOYz5PZGa/n2TSqcx3
xDNNWIfR8lPxTAx8wvwP1k6HXZgjlurGir8UO2u7sq6AVLmOUcWf3vGgW8KES3XV
QcUl7tVLjkKjlYTf4o6ndM6+v7Oz65F/epP0HbiI24WFkePKcCixTVrd8qKee1kA
Lp8KbWrVwSTQSLx1IBdAnN/MVot9Ka6FIKyHk5FakotdsVntm6p9DXNvAnJmm93T
XuWxc+37Q/rpRzTYnCUu2y19wg2kr2lyzjmTK3og7xKnB5G/emwCZJm1G4baihaZ
eUxZR7pJ9ZFZKTRI1+i1PSzTfQbUVef5/cIvTHLl8s+XSZEANX4lB8gel18mo2tA
Y2+nd5IuMdTPbyPXlBb39l1V43aMof2XNCHkr0DuXFh030nn74cYOWYzsZuekgjx
htcUbcRjuUL7Y5UFa/aoBYlxvOU1EKKoCa49YgAEkZKVk/gsUR/SclLy53wyqd0Q
8TN9g5+Y3XkCH5xqqeCg+b42Azcz3ElIHIOMgocC4uF3tmdtfZY0+t9Ncm3xDhO/
TdyDfeOKe0cPFH0TB9p0da8FPdJX9yJjXCEZZDqIALgGqiocPwdus8x3HKpkYlad
wql1HZ7oVZBmEJ4WOCmy3ibS994OVQYgZ31YpsXWFZjfZlYTmi4+xrag+G4CAh3F
vgKVf1mJlXtMgJuGLdT6DF95c0tYbuD3zjeZACmS5cAR93/PAVX8RlMj4xCL1uhb
c9zHNM1E0xc9KqRHbnQ/mDMwFgtQw/nqrvyPc3kCmjTRe0A7LyxdKHpZUU8lq+M9
bl+ZRMfQ3avDix1jkukRShiNe9SNlyqockz7QE1N9W3CQwzywby33Tq5DKvc2Nvm
ppD7eLDUp8WNDtqtGTCl0by1DVwpzVBQ+COns1ZAkkd2b5X37dhz9ci+L2mVNmgY
Q2ZX9su5+rIcepF1TMustqSy7sV1l+MRoPqVyHNz1BjNjK6ESRw+zqZlkCGxXa4U
VJtwuVCXuG/i966+g9RROzv7kgwEYbdRwsZzkVL/Vu5HlA6JbM6Q9iZCY918oVTQ
LxRpYbj9PXjsoj4Sg3omcCL+g84nqcitvhTDmIraoPRP5GFG1CNHhpv0VqdKUm53
SNZRvOjZj5EZx4LYVB9TAMh+DVlUB/LrNb8e3llnFDCVTdHebvQy9ceSxVevWgTy
i/NzcAbZptTbJpHb9JcimjBuhbRja48QzlYVnpIQ5d1j/LdQ1G8eVH6qoPjuf9tJ
BnoGWAY2QxgQgEx+ZCfERismePxHi6gcA/kOjlMlpETDuitEWIQwcObpaylWfkbA
5zwawkMsaKCi+icMP/BbAmZ78HkwsgEM2PHE779EspOgRT+4TPkQojXbjso2NxsR
ql6Reyy/OYjSPbPpz38kpcEeNNBW8+j+PDVjVZWdiHuCuFkzTJZrUbMADqkOkGmr
5iokABxjbg0205MHGE6RlLE1qQFrH22OYv4CCwTSOb7UqkneCVMunlBLxhACuKhv
sHhlEyoyrWyfOpNvhV8KUo+sg60O2xVtiwrgaTybHbGwqpeFWLjFNJFpA8R7M+9L
7i5bNDPXc2XuevgIDe6nnbjCFJucoVSSNUtjc51N9XodlX4CB/Jn23PbuUvSPwxv
Y7pE16uh/ocRXiV2H6sJJ+++ApPLjQSWgW2JyIq28yDLV3RAL0T95vqjtB/FyNdV
ZlwGvcebCtTr0qKYILTIVwEPq3voYzcrxfsb6XQtlF8jjCf4wTo6lXKky0qiTGGO
HR42Ya0iIgW27kqCkMczllPY1zGPOGENJG6gzoFyDHbNZE+Z4177YmdR8awZ6h1z
BjOGynkR/eH9wlHtn1WG1of5hCADmd2YfNFz6acVTxPVTTJoBrufOaucMVmIbRzf
7p5SeSFchLwekoZ9rwPN6ZY4JvLTKB20kxJlBUuHGLEVo7+9jMaEh/mzfuttiRIo
/e9EPwKwWxW9p4FTw6Sp+p76LiA9vjBBcKzB31YsqgVhlYmWOFDjkdeQ5X9unStH
kHb53Th+aDc045pGzmnq4KC7VWDKZaNXI8z0/yzxIPl2l6Svl+qGCg731URQUHUx
69tK1w5JJw6tr3iPxaEyaLYRJd1lMmEw15Mt+/2NWJGVOgRqmMFqc+/GsZeYTh0j
Ce1H1Vk5jz6jI9i3qCnVOLbaoEdA4LQkAH2xdei56IlwnM/a4gTrTiapO75clz5f
2h7s1DL7D2WciQ+hqF/gHp6tMQ6AETTMtyzsCe9ViwYeqMoIi6vgYFqqkoL+CumC
LT2cirBuVxdNSX69x9otUncCXJ9EBJjB3qaQHAWqloQxtku+V28B14OG5/TKutoh
y3klOIUSrxuCInE1+jhyTntG0rAlqRQ7SEfk/0ZHa97/1+V8c7fWazQdWU4ogUBf
Y5g3PiZWqlCtE0JA1t7xPSWd1G9882W61w3occpHGlFyZ0obwd3tzj7YDUs4DTXA
mQMIHD3QkN9UhRMnzkJvgCUeua10+rIzD1WknoXDDSBIc8jDTPx3MKexiUjvu1I4
AkHFcTf5CPB9BYp9LXEklAk3ziqJuW4rXvU6mZ0v/mMrQbkcI5SLEwt7tujoAOl3
dYiyAISirAho16HsVvcb6IKVTZHm/7cS6YYeLNPV6KjWX8bfTFsC8xdTeRY4odQV
3r4NifwXOS/6QqNhYoJRCLYUtDqpatbgSdBIW2tCxGC1WWQA8uJYggAxI/y3GRiW
AvDPAJDDjUunpmFcr7dFc8UZ1RDU41g3hkZBInafySh5/DIQS6PGowAmV8vS/jqc
1MKhoTfh0Cd9rHX2t7l+bAF5bxDYxEV/tXI0eI50PfegtfAzigmmN4+TAu4tl9pO
TcPw0ZoFBgjPOmjWzHwCL0FrGrjGd8T3xZe/gTpspbwF8hR1FA38v8KID/0bdgcy
5tyP9dygff8m4AVR5aKGo0gGijmH09qdMY5RlV5980CUiASirKvjC3R3wC/rp4Cm
+d+QaOLvljRU+z9xjgGO6t4flvgOZeywLTN0RzrzMIbnTngvU8peNohoixVq2QID
dy2PJq0or735RMFDppbLE/8jjYqSI3A3zFQnlqbQhSvdkvIcLyrKbGhfdAmZm3lT
1Ay/ZdvnaQYeiemqMvzGOYes6n9Yf11HEI4RR9cpyRPPo4uPtPdb3DsykkEoj0JJ
xkL85hReEqiFSA2HH3EQhmn+PxqCmSjM3z6HxSFAElnD/3H9qX2wqtkd3Rnhl/VQ
FsW7g2ADykZqwEQAjl+OScOql4XC15SjzjAIeFoAFtkU0d/qbsR0+vS72MB7thqp
uU74PkfM03ELYay53B6u50/vJ2XZJBoVQE4UZABCE938Eoj662zgsp2hkNXhSnUB
Vwws2lMIsBV4Pu69Bq3nlc8khn9AIpHoaTxW6NGj93LoUrioAFsYLpY0ED32hNcH
xf8ADC+YXJbuTyPmWylc+y95TaklONEQMXSQRDYRA/g973jl3+ebfNBT9mb2NXPc
aQGO7Kn+Mlw9w09ko7NGZoeD8jzV3X2dan3CTf/EWF/qSacQdfPSP6I5uHfuarmx
wzBYv+jm+iUxuPfRMSO9rThbcadBMKx+DCIBP+Qkzq3PPy/E1xTanLS26KPP4fZi
ZlLiYbdIrOzxX79Mi7+aqVEWquzsdl6J1nBa/MAVNx1ynW6OYeF/CsxGOwO/ZWrP
Cr1qVJytJYHp80r49B6VkIY3T6uJS/trnPSMEW1WHuyVtOOfIT5Qt65sjZN2Vn3p
0b97QSJVqNDbV9IoS6MuIOIW+Tx0g4m0XpWMsJs5MC01eclcXfxwFi+B7iuFOvd0
m/2z/ytmdtkmr3+A0pMd+3hocVtbACwV843ym9VhTOasjW9X32wBLPhq65NRGBvP
e1B1o7ZuTvV2D4xFlRkezaeoktvZ+X3nLJ49Qlix0X4eqeSCDOmEDPpxGoRHQ1mz
R+W7IdNAIFgCXLj1IjHQQx9l9vzx8/hdK/Ir+PqgCnEjjwf3rU1Kg/WE+tgjVLiF
fyMmg+xoNkbT8i9tUGlYLGDSBnQMQQuY7XmYDWo3cS+irl7vavlDl1Za5SdhIjhN
XlZV/QOJxn8x9zfllWQTj+LbPOySgT82zL1joPj84yOyCCgH037THyIW5OK3jmZH
bUt20KAdo5v8/thEpAA+RyCR4TNafrzLvdZKBajnZiG7sf4ocIqSt6hB8UYNvu9o
HrsbtshGTtSWZuR7CfDQgy8G+R6G0R6O6gpxWpxpyZOBzcboNXDoxCas9i5re9sl
fnl5PaKOdQ16W/bMTm8cZQeHout9PsgvbxgQDAB/1UDKquzktmT+6kplMRE/drVx
HZfJgmJP+piacoBCAeWW2ZlSlIjNZtczV4Wc+KiHH3CjCnx7Y2N2+cbhrkaH+PIM
h1XrC87UsdwvZgBlYHue22zkEbj1kAIBf7RzRjAjTSYLfvxHTKd3CvpEEs7BxQbc
hc6Sft2owsg+rC+JsbUsuZ8FUDwCrdYyAuQRdCbgTXHf9hglavFT6oSaY6V9cLQx
CShQKFeq/ecNpoDzpMqgu25idwX6UswD16SyA0dv7yRWLOkW8AzT1bLoqRa2ZLPg
0SstW3MdoinXQSj2nP62N3oeIko9D2lnmZNFA2t1wPAEsoh8wcHeMJR91rELEdtn
c63vbOU++KP9G2IlwDmq0BeuIE8YVkV9GyhqM5vS89UvXdHqITj4SrhAjP3bZTUw
TXnl+uRcb5aLwmT+pB9T58Ai684XJLcRpBYWW51RPxuxDEtfntkFxclH12f2GP+Q
p6b1rHcngMVu+VUkTz9xhyvo9bOowqjdKA+k9nkFDIHTQUng9sfyN+YOl7LLxWrF
i/jxkP37hC2kJ0TrGBXbTKMB17+VHwXOzlJoXXb7NLr7SkZ1fkGeCldOJqO6iZVd
VdP81I4ovPT/e3YP7BpJ/aTAlRlWhAmfaLRDRjXd98eSAwMZ629i/gIPcZDZaTQ4
tQo876p4ZYykEL6RAUiNL67ckLxWMUM2pTxn/fcSL9LAuBxtplzZSQTIStLRhXPc
ik5Nl/bmkKWLKx2p+uHx/bpEi0hkMEoGMA+obHXjlQRt7hYZ0LYD8k3AAg6lAkF0
N/E6OSrxnBcdpSo+v8LMnDqbpCY3ONJhulwqKKbxlzbOX16D2c/8AV9PoyP3C+DK
M68yRuZPBc4G7RDfr3xE6JFXRiWSAQ8HsIXFAhApyxqL4iSgh2YEgFn0Dbs534r1
leWGCix4jmOuYLgXq2Hk/OiwQ/vU0T1emQuprMUKMKMaj0veDHYUdtYF4YjWKxvc
k8a2bswuV+uk28lXZGzD15GKfV2BcoLfgCqr/ytNjDZab6ZIjQacY5LxJASLYOM6
S1dLLGHYaU9nRHn4f1TproBkxtIbKftyQsZuLfxD89LfciVfDEMW/0uPPw4VWAvC
dDm7BMlhODM0sEK5wRHPY8waJEdbq4YAQsOP9f3B56dlf9h/8nVBNMiH9qBGvJ7m
d+vfL7vmeZ3L5xVlIqSnEaIVSA3jWBYsh2Qoc/lw3dVjTCagJRSl9wS8fjv2C1C+
NkxXUCcNXimxNrcrGdEdqMnT2IwVNBaLcofHoLQcXEqVeUtKezukqIKGVOQJOFdT
9c/xO5U6S4g+x3/sa3b+oaLvArURN8Lf7Eh/tGpnwiiDSJIHnEZrUyCNtaiNdjB3
JTMxebZ/d0Yllpt4lPtjf0gIUJNzwNZQ3uMHMpERF2nKFfz3vf8+IpV2VtCwEfcQ
9zuZ49PhOuDwkKzZaDphMlQSmoQeq89qmuewWnnTQC0tpMpiumjZgZy75jom1Mks
vgSgJZJ/DF4lvHkluM5oXKs48oATfwtpJaqybbsbJzDqz//iJSsv9OCbROIR+cSS
zH/PXb8XHvkyFqZ5B4xXSmanTOlSDxVztnbJJSDcUIhh8wH+7UwIzO/AwcuOxyae
nKygYJcXIBwksLdoAUZsEXPDFTvFVwZ2b9qJ8515xVpQuzW+u7u4HEKAx7Er1Btb
lc/YMflUE2jplTRJP1HrF9Rh3YRVbJ7foFGsNTyFmA7PHfPRVjwRLukvRctFPSLs
tT2acYdFDNrTqSMVpkHISu9sgmOlvrDGSo/0SpKMeu5C1G8IahimQvUIrHUSuJy9
bELNhpofOOztHCZsA9C2Ox5/5mAd873oitBRWHZhbhQ+EqrQBS8zhbkbX7FYMxhx
z+77b035fqEFBzHPiGT68QrnDtM54gXmsqoNxMzLCgZP+kn5xrGojapDM8LfC3//
e1EYm4cE7tJEAnwqaYGIkBNcqYrIvHF4U40Q+M5mgZDs3kNWZoS/ONUWuBG86ZqK
pF/3XSUF0QRvEbOIBQ1jNK6fFsBBwyCYWa8KFTb5dhFk09VEoRBist5k1V7Hopm6
ALQhAtbryxEnKywl+V9kIIzAFDwmXvtrMqSPSz3+KmGCcJJpSDPaoBnuBReMBLlz
oSE24UBjcyxRQCVJQZpksDMt8D48Wt4ZyZ/6bd/mWGQZYrv3k2wytF8s/cKHsO2q
nrkW4NXz01JgFzhBsqqN+CCV387xgULPClrDeCQWB8L6f9LpStTZ0QT6qwPGHygE
1DW7H2nm+Tui3V3f6h/2DRbNdhPJSDjNjxOHo7mutZBdOMhBMeHQA2EE4JYF6bbs
gZOcjC63njbSVK+vG1/x2rlTGyzSXK6FXBF0pdO1x1EmvQ7/4dF/MR5pjze/mnW+
7SPBZpi4caH9GT0jZc4tGmNHjrWuRX/eA8KxbLoVDh5pgxi4SOvNetGaZV+OcAaN
ZSu5URzTm4cNhtVYbAH72YG9bxA15G7zZZnktsP/UqNTWSrv7ah3QlBsrHo7ndz2
znR5FnTMNYNT8KJNroknQbNFQxyXXie1pkHYbDtieChqsN/iyktT6y5aKYQsRoCO
oDzUwVeDi8lnXIW2pkcJS5KimXVH2suD76JIOJ84ULcRFQAC6shig3NM5V7vg1Mj
3JB0+6eXEdiR7uN7+aql7/8R4kf093hemWoQrVjMhvuMJiqg4JRCaZJV/snVMa+8
o3eGkE6wEvdsTdPo2gY71qZx5grn4rV31pIhlLpyxi6TnuGweIeWYYI+ECkJyFLQ
Q6ZGK0djpyWlvRcFqxNlop0TdFNPZ9ezu8hmz5IEocXV25/wN0I89flgMJwcRYzz
6tQ12FBDInFy2ECX1L0TkH9Pe090QpxESZRKuzUKUxrttdGyb1erlkoAYsEdErJF
A6Y11VCT6Y/6QJIKvJUTLaYmNOO+PcZUJMX4j7Sd6gPUfnLSWq5gsXL5j4XpDP2Z
tEy/Ki7QVnx6f7xChAE3KqqAOFU2ZjEC957kRsC+4M4Yr0KqmkeJrJIEr0HaYOeF
8dTcf3jrFdYDs77lVkp50zUQ0ywRuwuy+4JlHwsoPhfpccVm19amb6a2276b58fY
Wvl5ggwXzCXdkySxyZEBdxlpL5fy/lkKgC64/vLJhCTHp2hY8eJQN1kYCKNH3Ybs
I7PiZ2GqrYi7b8TqWKuh1LA+ePmvzniB9RlXtj0GRoxhasCvrMXdapyHVxt6EZBl
/T+FLGE6HyzNUrLScA5JCjnxdwrlI0bj5Mx7wP7B1qi3gCkrC2fBcqw0Pl+jfVRw
JCkjI1FflK4aEdIvqj6tFnTX/7BOT9M/TD74piMx7p5KjKDIMCiy3UkC3UCooL/9
aFSvqXEEo77IViI3fGAywheef8lbCuWt4AgX69G1L4bNLOLsjhwM/5kIVScxcJOj
W9IkWXCgmo/W+H4IiqitRqxUD/uwxMOn4tB+8dpXVtplBLoTaqHEeEWwtg7XyABa
bTb1b+MjcvXlGOvwTie/t9w+PazSBk1zzXcDgTvZeZCf3SNPdoNgyDy3qBtEZoSK
SsyCA9Sg43rYr/gddWFmUD/FQebEI8Xw5ICfeLEtN8vKTAO7rux8x93dkpH0mtyT
5zL5GZLkrVMYckVBUgCzA2ceoHiGTSNrRQ1DchAI2gdm7P6fTBO+WQXxU36btM24
Es1hhQb7mQZmqdeSDRPQIdnx94+SVeTyTHSzspV3iTKHR+/tIpZ2LyGaW7EFuXKA
VM/u999I64uNZzNtR7HPM7tuCV8GpTz7mW09SBxwd16NVFfmuCu2lrdSEU1Q+1qW
dbOctMi9NO0roxB0AKSyKX47m2IkelMMsBykew4z34zae9YQ7LFVEn05aAE5jSS5
ttp0qWmLNZ8abOhYQ26U/MpM8VZgUk4ptsYqpoQCEFSivAFqQe/99gtWGItt0be1
iu/5c/2UxjwB+3xuOq6oel0zSRK/HhnKgvADzF1A5WZl9xWeE201vM5++CFJoPbi
lLPXDA/R1HAeOLQvVW5FaeDz1g31z4mvylehRIeXMzwF7qvFwr+tebpQuT94/p71
duBtWOs7t2X2VgdAKam/eGk8DITzlLUZQNp062KKwe6l1XHHHGt0zipzE41bhc70
WtOJClIOWFfUa7E/vgD48esNPX0MBW6z+h4ZoAMvviFsBgmTLqT1zH6uvv3UOygu
Ju/hnRJ8yEaquthiKY0kZD56yWGs5mJJMeBy8O4t0nS7nBCL9oakOFY0JRE4mdR9
44VcJE/Ik4NAGy2NuK7FQhtnFichugbk4NR2DBw+X2vY1sO77GlQK1bNOvF0ep5i
lrkZjXjdVqXw+XjrtUZXlp0UyXjvy/0u6ydNZjl/C0VymmilOuIIkNxXRcdzspc6
L6ExWVLPYTrPffR93u94bhqSpdDNSFm9BOrSJntas8t7jyDjEEpORjzZELpgm8SY
QkLnrhmUnHiVe6cbsaAgPS3n0nmj/Bw5VuGGARXNv5J5o9SmQdVJV+zafkR87oU9
4nvxCbo9Kr7deoUT1x5AQ9lCcxvkdn/2mARL2Tf4bYUcme3SOhLpeKfRS8JJgKvV
SBXXirRGMEBnF0R5Q5ei0X/ugigPW99qZb4lnv7/FvkkZ8QiZMvrWp5XewvOzN4I
LDKtOmObkXfTRv9yRQGyurtUHUklTcLt5pmkH9XIM0MnN0ZvqmSjWmDqbanuKHZM
04Vi+FFC1rx5QjTDK1ntdEWKB7prhRQ0yP51i4j+ICEyNFdBDm8S97/Vfe46iiCy
vPRdg6zaFzxwIJFUIAEdq8ZF7kF5vXlrre0b6F6nyZyaFCllDlHrWya3/0As9nTn
Yz7Yq23jG+KmV7nXF9J3PH4e8C4wO45OfhjkNNcWNTvucEruYwFIJc15Recea/2f
OKOFMR71t0W8pM+s1etycU4dBPNIPCWgfM8idklyhMNDiz3XFZ5/FMc1rdNGXYrA
BH0m1iC99TKgKL22+C3nS7g8zP+akQGWlBqJ1tO9ajRKw8SXxk1jD+/T0LbrVCFm
KfSMj1xEEft6RuC1AZb7G1INCVR+wmvfgzsfhqKVeWNbS+flHdhDBdObCPrDSzX/
BFXkUbe4eLB7d5cBVhNnPlBp3ieeVSw9ABrs4QqcqYXbBq99+lGrncEE7vlMhueT
kiVzPPqTkUqLfm4bPcEy7RIhBjGI7Bd/gnnrAZY1z0ISX300avskaLqEMzzE3vWK
9YoNEMJZj7TbYfgT86MiHBE+HZBw4Z4p1yiyBq2hwkL7X/DZ4ODnWJl3GOVvjlgy
2lj8eG9+UHgldMIf7ND4D0iB0L0BZNYZafxtagKI2r4IhZQfpxviXSJ1B7YcAthe
HuIktUURMWjgy0sb2By9jIqzQWzkJQE4PzJP8K7qH0lsuHpqUIa2zOyWQe/8DyGq
jhog/ep1vYKk8Ma9LvtGHYRWnN/hA0sp+Ev3taSCeqLsTNW7tw0eM9NGuzrNsP8G
js5CAhKQTWyiyGZMfh+e4sebPIBsMsssn/QYPO0NWqV0leSVbaX7xFkj+nVgnMr1
6gsa+rvPgaVBxXqhbjd1y5WSTn8xtbpG6LhXHoiVMqRSoTqqphZD1FXz5eiG2zZ5
QyhU74jqRWIV0mprtocGlO8L6B4H6T+IEetOmn7PET87EwG3w9R1hG2ZAja6khPN
qUvl2Nim4StlLckDRnXsGRv4SzDwAoe69fV8f4y+cqc5eFEkX26XeuW6ZLT5FRdk
7ifgJd0IKKm//JyEtu8d1SFKPt3AWyXI6CEyZ6nLN2SDr42ZDghYaixyr7OIzHTY
JS13pL3+28wtw9SIoI4azY7xWXrrpmIvfi7R1N1AYhPNs012ud6yroxHHblog42c
3yVPqbGWhjwrrx3H0BhTJJ1Z4WaTSET6WM3wbwAm82gARlJWegl9EzI0pjtv0ttX
BfZbDIPiD3cCI9Qe7gDJXfsFX9ACX5xUfYetC+X+pxP0coY1FVTNpDxgVC+pOAWi
+UNHF/BgO50Q3OpEd8hypPncaIi/vzauRWOO3wH3x9M3LoVQhnv666RDcCp+Oddb
8Q8TyB371O9zCab47aKieSRW361gjLJeLif3g1RoS5WqmGCO9+jMupRrq5M1cTVO
erieSLqGCPvYy7z14DC8oeIZEmR/iGvJjNNoBExOlRCLPAqUPnM9n90i4GYLfFs0
F33kYVtet9lWtgJ0hLr2XLNHjcfUV74Yk23zhzs3UiuH4FwtQeAv6R6EVGAoW0By
YICR7ahxsL75PTwQ6WH61JlMRNZEiJLU1y8KKHxUN2uMh6hsjA/yy0NbVZcj3ECp
yPypRjDQt31wSuXjJ8j47HBr0PrRkLiT3w9jikb+tqtFsM85zn/6KjOvlh2HTxOc
rz5dy6DBuUidIgBzeRNcLTeL7F6JeRu1Td2OAtyXyPGfUBhwQ5wXMglJyVIcSQ73
SGwAmHvq/D/jGi3CrC4+5Bh+rkX8pf4xz+4OfkncDfRAQU//G/+mRkHz83hzRXLV
XT7ATgr+9TK+0Ue2X5ayZPDIEa3rhPg0RZzgayqJAgGSY9QOGVWzQV1DQFei4L5p
64vo7N29zONxkPCED70HkubozfniZaM/gwOnSTfaOrRqdhNIrEK2qaj633aHO8Oc
f5jSCfQjf4L3FfBOQpuJbbED8f43fiKCi1QwSrL3+VldKEFOItuIe6q83fMGZT7z
Yptcy8mosEmQ4q4UjqJjjnwssEGbzQPRc5zJHKmVyVVE6/kh4E6V0vw5OMOxQf2V
5cgsDHSApAe8JxhyGuLU8a0TtCKn4yO+AJBVLPr1cIl1v9n7KR3TIC9fqKcWYkU9
rFI22Tt1Si8/VKPPGxzypEG+S55DurqdJVrfLQ3EJ6P1w6Ar1FxnScxUldVE0UiP
O0WEx5/sbse0fy3K2cC9YC+6mmrjw4cQ+WQXRDmh2ykt4fyS/Bs2y9qOZRQTjD9I
9r64wrPYF0VazVwfOA+tIwcovdnf9RfClOLA6FMqWafu64w1A5xBYFOXB40HejUw
teSBMm9wjc8ThXRgrMsCxheIDjQ6ztU4+sBDfqoQ0/vf4UQmOARFyBKWIRLllXlN
FICWkyFsIsslO/WGG5DsaSuQzlSp+YVRp8eE2oMTuWNksd4d7l0+PLg/o0FzXEY9
qsPrO/DtcNUJSIpD5GyUJeDxkylcxSolHSfZYSf4Kz0jhkrc8rWM/H0tS32GS+IB
GHW1FleA5GZtHB4gZkIrdm3RRax72+jX+gFQ3Nu51FIm0UZeFqnmVV3UTa0ZNEJw
+4HwlS5lrf0UunCMg2FR0jQrEteg8NROgEs2YE13id3LVXtMPVn21AKhKLQL/pwA
wEmJymMsqb68sp1RnhF1w89igyp+UzoV+avCwKJFvb3lljNloSdxlXXBMo/7I5Ks
VwX5QKicjthpJKyWphwzTNbhhGqhu0dfDbsS2TG+gkyG6jQpImyhjZimiae4q/9b
125auBxVNHQNmnKpyDpTMGlqnfk30euR3lAeKwd+z9591qW+JLSig2Ka393hHQe6
z7Rwojb+7HSgwaMX8c+XK9/SoK29xt1MZmyfJmknhB1/eUkCpmtcbQENIbcgcU19
ejuKqz/LKBHoeBmtziPbvjAYPGKqoN7V4tPoUjDghzDehoGGmUSDVuFniPnE2vkT
enPrtsaWXw7ZzTPLVzJBdg==
`protect end_protected