`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 2848 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/9huKRhRMtvnNqb3Z+UU7TahEoHV+T8U3P3ufru7l1O
3DlgtZzb9QxCbOjthp9+wDkjygH0eUfDrEl1ovhZG61oZWMUaqCow03TrYa8PU64
JX1jw60LuqFp08q2yJylSNFIOsyFrGk/3EsyJHyWqNk7Ru0eLhTpJshK49k75B1H
/QWolK0NCpylHDJ9tvJs4glf3iXxbx25OasuOvCRklEflrViWbbkG4+oAdgsJeOE
+12UdXCgMDRdfjvDYtO2g+lUM5yEzKDFmWZsxLMKZpchGOl/Y/dY4/hYZtISsrnb
/a7tUfN2JTj3bBejmnbp5M9Oc/lCD4LbKQNQu39RtsgSKfpcqCXwbLkGJe8Wu4Ad
wsebacyGJOAd5NJ38BzojnmiYhbDlwdxGXOItc9/OqfbjhIwqtQdGP68WWfIIL53
TKlbgsEVu+S0YouPkZQvj6VMqSnI700uIPWeMIey0jv8f7o+KxApeyJ6Is8T8XWV
QW9vbPE2NdEsn+tRgMRCka9sdYAWqjssWkAyj6Cc4s72hWvb39ySxsJQGgs2gldj
jb5YmthSBnc3vGte5l/C9thlLIc4uYpDGS6lP8JSeRDJuH5AQU9l/R6d6/YhT4MY
3ImFPCY1lVcyGexepro343gSkG1m1ydH0/6KSPDgycSFN3ge10MIlMFb5HLg8e3t
MI/4+lDLLVv3NH5yrUPHc8gBqvsAscrtWdDnPfx7enMyQaTw2tROqY5JmfP3zzrQ
BJtSSNffm4VzQ1tHISNhxTZuvHWsl29nO6JrwEIL/dpIDmMDeSdJvA6E0ZX4HZ7y
NQYw7rjDev8kUCnSzt7Dwy84oLJT0oDNfTwvs/kD7EFT7dVDY6seEa5yUvf6ii9b
faWn0EpBPU1E9TXyvf9k+/LL9MwCWkxygVtZWHvReeZVF4KGYUbaMeohoOvhFXVr
P27H1iUVqSEyqK3DSlaCFoQ1MWLw9UDVIiL1YFxCMxxsiXklS+lHhlKhSCNPH1fU
yMcE0xFBCS8K7U44nHYreqLIA/CinhOtvyWJzl8kxfISXozNLNvvm07DOTN3xZHU
bWlAd49l6viqd8k5Ng9V6HTI4I+GgFFAaLTK0QCuHQkqh/r1Uwiv3vIHmHocgE62
2cyYl36Li3f176ntvn26OSmlUgoZju7lFT1ACN/QhAKeGrjhn7dcPpYdUC+jQrS2
hc/HLVKqhAawE3zeIiGRBPRD6Y09nQkSP6ETYlkbZt9IPJ+UoNMKcE0d6PmSoxO0
rO7+s1s4TLMnWQMHWFmfTyrl1tcOJMD8vWNIlfa7WDZSJSdMVBsSIWItURjGF/tL
9T2WegkZQIisSxypBz2WSjR/zQLjoYGjJLHMtOjVk9pa+hG1SE3s35CkG9JUG1tY
3GT8yURcHPT0GxevwfQNbufq7OUH88j8/hwR8khbRL7DWGzP19CJQeHTG+gaVpa7
ahUNsraKl/fYnguqANG0rL7yxPSXNt/ulTJVnDKX7VUHJwXav+q4zTU89GQ4LkLk
r+Uzi7zG3m9eYaxi9MDbF1DPMDZoW9tk3dDYow4KCgwZeZnazK3JNTbhZHBJRCX+
Kzs/YUCFDZsScvh3LmRY+BR7QdMKdV+j6Odlwh0nVfNSqYUw8clA1/4gwDvFv0c1
84pyk0qmCtHT3oDC6KyOiJOcSwHPn7Cvz1m5wEsbIOPznx9SR8mxbYwyBe6Fiwpn
FwGCFUq3vmbQvdu7d63OK3liBCPNTQz0KBVnf+JrtIkRtmKFFiJCNIyicqIefUrY
kbOvm+RUWlqw8/uoXWgEmGQhHSq5bXDQ94DQq9tkrS+vjrc4ygUUYrwMFJ66LqHd
/KBjpatTIhrYCOZqupoDinxoTUUW9uj4KntkaOrjlNeHIpRZYc6ZDoORn1ckvBcs
qzZjc2G60wYBgQcpaEcqDoOjoS92JERR5UlrquklkFMHO5VYsO2VGh2mwfnWPGkc
+2J+e1WnPghXiJL+wbddISWXDvNYNDXyS65BvKxUDLBgtEMicKu7Mmjd8/mK2xNN
v0F0DlFCyFp4v0op22TSi2OrCNPYc/dWu6QPgNMABE6rMgB1njzWwuees/sgi6Lp
kVIiVGEx3mxUQhZobRYgQzsJ1cnaUJrFeeYcMCjq2yImvsLVbi65F/YGGtAAlf7e
ps668tH/8r15hQnyUSoMGcUUgMiJZvsxWnozDqp+Afn3F4vTNsT9N1JqvB8o+ReV
ac3Txqxy+tK+/QMubOhIJfH0zsjyZ7rjhirOguHu0PehKCzN96TpH3pGvozFE8Vu
5OLPMNqBZYy5ojysZncurgM9T873x61nb8gxuo5Pc9ZYkHB/Yo0hWf9zNAt6NReT
ENIODmoCknqwClRBWRKDZ5PWxma51S5JUj6kBDGMZbTESu92rX9Zrh1qMZP2S9E6
bZy8CTKEP+f8+firDovh0tOgOpACHdcspxnH134z7zB5C7nN88Dyof6v8Lj0Hmmi
chaR++2negtKiK2UmnFf5B+KHYq4NcsvZKqCMkDrO3WJedZKZ+dl/ZiREyPuAtq0
Xk1vMkNY4FMjj7VoRBKfCKWWbztbOzHH49KM12uRZDYtj62BjLakJvmiw5UDe7jS
nxhi1+xjxX/TdZZwxDCK9lO7gM7HBoz+rDey62ADfXCSXREDv5xTCRDoCerYOgEM
zHDCB7j7zi36+BZFITcY8D6wf9OMJrlqw2Lyq0Ba3S+tr6dYwmNSBRj2ZedosiAQ
1LvXTeZxyFmGiTsNFzoRGKtBnwf7HciqzsoeeXC5gKJrJBERjIyrgBN02sGp6kXR
Mmo0MMaN1FdV5ZXJwluDtHsJiUw96xtUWNp0qW/jPv2qmA/W2TlQhli4of5mFty0
gamdEMTA14UykCmzyHLw3+4IjqVNquvqLJgstSF/IFPzzau1M6+1naKiqc4U1tP4
fh/9IE/JB+f4Hs8yMjtrUGLgN4xISBl8tcnV/xVyoN6q0Ma+9UFnyZR+vDjT6R5O
V4Y6vEjXy5l7JzOwl//lls7YFQFwY8vdpDlbp2Tal4G7VFN6VqG6fzHIyvkQOPYr
dPaMpYfd2SaBFt41F59gYg/RJOzJ3Uu/pdyB4d4JSSYYEFYnpXVi6cb4hijWDdO1
V2yqyHXRW4UrV1gEHXN8mWvkWd+1sWkvmMAV/KsqJqid9fns6Vr8PF3pcnwnNM5K
a3g+Z4p9GNotYKvWvJr5yNK+tjDk9SEZrNVXaYG689mnQb/FKKlvLb2jn8Wg/YIY
tUQG/kl/gF/yNupdbVFxjzkP65wAFRuzpyWt7LffDOgodUz6q1JDyK0KlH3ypSZb
IEl38OjzQbWxWQHKFLIx2+76PxGbIfljCkmIFdfc4EHS0EPcUZNlzU1l2u4FwA1g
iKwwmH9r8kYoophd/qXowSfPvmwj8+mcENBz90jfJ2dFqHnm7h9aqaFXL4T9ENrI
qAoWsyUWwGbBAjhYJzNhBLmV1ZdBma3ybYDBeoRXHejgu3ZpXbcJquWft7VoR0lQ
dLE7KKUm7jZh/+8W2bDRPa16uSNnKawmv5wTY3pyOHpARMEzKtPi0lynBOaeWba/
Ns1G8zyMUBU86cKWztLuwuvOSed2kUVLUjPyTiuYD3038ME479gSWJpKSYJJ74Ne
vpRaKOFRa6aFz6cNIzY3bIwjbANRnavfw/WkXjB4xEatPEI3hmPhS7bCBA1XpF6S
gmcJ6e0EcFBVYh5mtH5HYs305SIBAlWyUZFpZ+I3f31WjtRt3LAnxHgZlxpvcarE
DZrF+K9ewylhOngC8MWtyg==
`protect end_protected