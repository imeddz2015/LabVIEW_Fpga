`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 12304 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/9huKRhRMtvnNqb3Z+UU7TahEoHV+T8U3P3ufru7l1O
3DlgtZzb9QxCbOjthp9+wDkjygH0eUfDrEl1ovhZG6295zs5EtXcjf/jST1PNYcx
jBG/2nvj7AdhHk8/pmIsyXZ4Pn65H0aHZbyRGZPg2wDaPnqoqf02ZEaNyAHaWe7T
RxDONzn0u8DAISXkUf3hS/NiqaK4052fUX8w0PYl1OpGV5zusbezu6Kg3gTeaZHK
mJs1/XxwPgb4N+RrrZUgI38poDnsynV/wkA1RiJ0fQ37LPQU32CmNX8mRVRNEFdS
+x75BmwVyrduMR4X5fQjunGMDH+iwgV3UomQYCKRzqehkmbintOZR/gPR5pgGGvk
cB3UN98LaJ9pRLfLlglcC51W+4XPJykIQr8I4OZaAX109zzlyMbtwXP9A8WMU4vX
n3ovR4h9FphESfnozfyGM8uu12LslPHhpw4tXti8td83qyptJFgOvshECra3Vyk6
HOyM+eoU89XKVhLTkOLHP036TZUZJm+P6/fdefYBK4BFZD22H4IR4fNQVFsLpJxQ
yxUP9Q3R5fYdJXi2p6V9gQhbQrnYP2h+tZKnv/50TOKS7qq7pDZ7SSRG+1WrOLeE
6LkqZgTiBDSwvtN4hgErPuKNtzsxSVZ/rKvhrSvmzBIVhcDZj7OkAcTWOoNnP//n
+B7ndl9uj/L7p/lsZoY+G35mAg+pX/FCAU8tApxvV1qUu4F9ITz9Xe6j1WiPyaqX
F5ACNBbLRvI3gUZ75BC0HUEF7jn/KRvwVb7I6spy9jtMh98EU7FNx2s00lN3kLHv
85mCrwEk9io05fBgMtODZ9FI8oXP3SGi/Puj5dxjn9uHY4PpFpaCXy9qGWwoqvSx
gc92RHja0/UDK+f2KWyAbgpBY5MLUK/hPhXC36WqU6rzF1r0Egogdr+47Pbz59jM
h5iiz/J72QlHxkgciSa+XdVnHCSZR+YY8/MBjsHI+7DFP3rVb7wMG44dkORoDTGZ
CaQqDWumlpcNWrJlOwkdWa75wRiCUiiFZ3uz8O+kaHd8S6NaGuY0ypC9oiyIiShy
ayXUzdGAN1stKiuFhtxDlDAep9zCp2p1wefHfXrF5oDO29nIARnreXM1JyeUlTLZ
rvrvNoVQ79/rvFrBzIuR+XZntnPRxJX15VC5t6bfG2X0qEdUmx/MIi1CmjlwPqmu
OWU+mUZ9LaeA8KRjAHDzVzkJksOHoU7Anq36VPvka/wRtq/GQdAMo1aMuKzNpifr
YVdy/jotIhwZZs4SETs5FnVRfn8vi4LgXQz3HqdZvZ6t7DB9P/2/yD2uN7+XDxDj
E+/DNyX0tUE/5pwBhuQLnHL/2K8kiFCWk7ZGA3pbbCZdbzVglh+XqxKq2TtQZcJp
SO9x5xw0h4nM5Pk+QfskcSIi/l3x4+nmlrYwPcjMih7LX78i5gd+cp6+qgsHVzok
SMqbHU/oTc9PYc9Sbd+3qpzSnjeMBRf6LcUJH0ClsVyhxOz8O12OG4NuZKMmdj3z
2+h/e7nRKP41rdyd5mOm1X6fRveX3eaA1BtkkE+KyaF3Xf617FQZDu6f5HZglvqd
rNk5a4c64DI9TsE/1tN5iBmh3pnXaMBIxmyKw46mZTqgweGCIw3irzcVRafry7st
yT2hpuYMx4ZquQ5or+INmL+tLhQNsbf+Zr/DoL/X11nFcAKLVkEt2En2yFzWTp7L
Ny2QPaAUe+Zdx+rIqWUX3iosqTHAuwGnXmRPR3oQd3PafnKSjeKVqnznJPqMnMej
FqizHw8pbyMUCoqUEsJ5yYGR9PstAAjkc+3iBcLNIiM9aKC7e96hWhsEuNWxKN/h
S+MbrVVTdMQ+2pzKiuTqQ79X0hGgl9XySOCgtIM3UF9N13e5uXBH7vGO064WII14
2IjGzhpmspINQRd3yh+IhNzFXBWENf5Zl64DNJJ6zibkdlXQ2oj55Iyji8MnDQEb
0yLeUzS0GFEGBV8R3m0TWWhZkAJ37eqQ+C+n1FG8xEJQPoKHY2d06bLdnhUJ7Kk8
/QLc/UriXoC2XgjR4XxL9cpKFe9L4SDL+M+VoOJaESY4Y0J0KI05sUB7DBTGQj9F
V6Yq7ChvOqm/AVBkvC1x+Yc6s5yOaKyAwrF6TY//o+GFjcKNZVyIqkSt1n89IHD2
I10OTN/IqAWer9ZDKFPorxQ2dw3TPAXujr7gzF6mRiRIENz7Q0c5kkXpB+GbJkoY
YbfeQY/h99OMY4X2BWjRyX+4xWuSX/dupkbO+HBbI1gBNEUDCEJ7wAusreX31X/+
wsNKnFBQkmNiY08Bqh75A04+LMnNeXXP9mO/SdhIagNZxodDTYQ1ECRf+VcUcgCs
N0YQTqy7DUHYw6xx1gfTkUux45R8fcibnd+u9ZbGEB65z6/NRXoOSIeaF1tsjnVf
Sg7MslWZl7rlZvEGlqJ1AUJe4A9p4M/JgcENM6SQfipgX9ExI9N8iUWrCfLx4aeH
Y7AqLS1uGnM4SAK7IF2I1iiJoFfs6+ps42R5DLk6pQQOGm0v1sznPqZQ2MJvvsCn
CCHfA0gmHauz3Tst5n1sMYah8G+/jWvgb99oO1Y0BB2borB60ObPgaYTKrCZ0GgF
8Tqb4SHmksj36xLAyNWOLd4+urmoUzDhdWnon24zC87tFTYd81SDool4/fCFVYvF
p41IzGT2t2xTSn9YphxWCPFugK/SgRwzR799Rlh4FU0tqLPXZY4cgIkMD0Dq+KX5
0JsZsDe1v34zLGXHFsGV+GM9GyZmGCFnGNfMT021SITwof1Dv8ULyx4JizcFSUBM
zpjMNZm2bIfVTdmSPMfO/a1BdVQOT8nMhyoQFue67TGWJ7LvEooUxcgwH4OgWV3r
84c2a80bSTnNV+BrfroYPRheNUN4Iy8o3akcCCbu8fBdLgL8Ve4nyEmCY+Vyr/IO
qMbAR3fpMTfPU/JyWkuwmAqIqujydzQto9HEQe7Mh7lbh1cGnDzYqhiTZm+Tk1DN
3+GjHN+dXiF0hWEwav2YYCe3lti4REYVgbGnPA+SjGlpTYBHNdQalbNIELx44E6f
Y54rsHej3wIZa7bI+HHjAOY4sUfQRybByyrO+sr1iz+fhXjmlUZgoLdcXlW1wlE2
n+4kSbojQRtkhk69pH+vkrYaHy6JM+tSMtWuwZeXI1WknmIrsZO6MwIi+VXnOJ9c
kJNIKduasofr9sG7pp86ctQNfaEcEw7UQsE2CS9NPSdQ54XtZCw4SZstUlCa11Bm
QA2C1pmuuOzKsubDWOa3ecfk/V3xyZNuBULJTReh1HRJdtR/+60jaRlaYrDpTDe5
qR5UtXLOMswMFncsQsG5eMlpk4jnFofdxy7+b6ZOPUwrVOprr8diNgmUvHG1esMe
+GjDsEZpVWloT6ZQ9VYJSZGaBaObNMWEsNwO9Z/Io3FXcctqVXcZTESCRPLkz5Ma
JCnPcQDd+MWP90DfupHURYpa7mZVsIXaYoQmMY1aZq3+jdTGEYFCxqK8P2t9ZjQG
ZlKkf6RydXqWdYT2KB86nbi04YJNC5zIc4yXCLnXuD+Zah1mNTVUbc6NnWd+TADn
kg0vRg011/r7/EhAVgDIISArrU2M6Jskjzidmvc/18D0yyC5FOeBiccxaNZG8f2O
s2AIEtzXNfortXRjK+yUbhdNE8Iy8s1JroR0+BbZ2L1i7EVGanpjiyyJtNpeGmGg
PdnxwWafOgT+UILHIdMkmtG8R8W1ufVC59/JqBrYv4ybArIl6XxfcAgTMHMz1ZUe
DwfunJ60dN6pze5EI5SY/7gi9oX3DHYNvFZ2UOZImg8VQX1DtB8y1tDOBOMmO6mg
rMHn3askMjvC9RJWdlTTB/yg3hxZ/imP71/7R93iWaMAQ5fVEWN7V4cezLFu86mN
68R5NMLD5auBhnr3oLHvNK1rdQ2ovEAvQINQitXH6sg6z7jhekneb5ZwKei72z+M
M/74kZLBQaCoa0hMpx0hLOmojU35twxCD9CGAodeRm7WDuH2UMirpzZT6/7LF0l/
lNrI3DheMzL38tUBmSeZ2u96yCMCE+ELgqlE8PT2atJBBOEM7Vrx4JENuvOBVJ6t
vQxG0tmr8XNLWOUkO8lT0hJzdlCqcYFroHqaQPJ5DRsbyb92Q6WxaL2Y4WizVRRl
YcvWeCmsbqKxuIOR/9SAg7xNBPBfPKcSN5w5A9oZcoSI5cLmXyUToMgGxfifFgBw
Xmnochc2TfcqsiWxgCGZZxo9aaZQX+OQfA7NExUQ4K6fMpY0+BwhIlPSw9rhWvDH
ZJXt9LQkLLtt07yKs+tPnBAJDsZszMCywYSnB8YnLx+lxYmau42IXYo87hG5oeqF
0w7wnNIpaNBhf79aOR792R3oL4t3zd5/80ZOJGzo+GvN9zWFBizc8L581N2Az5gs
NvzAPXqsE+o92sDD+oT/L2DnfMmtiC3uX19bAsPpERGXAcfp1Ntw4oIk2xljdxTg
KTLwb2R+D982b0Riu1EcJ/0JZTs8ELobTlueoy7KpOuUxV+UR9eepKAjwd5UVe5Y
dt4ZWtS2d/UV5nYFtlqrjPhGg74Mkie1eDDUF0H58SK/UdFlzaEaYPILMbTIEXLO
Od5/VlPuKXUtuHHyiLArtVZNrJIV/vL2InA51ItBCMqGaOuAbDGo9jIZgRMBtXlt
iuSjp9LzWdNPIEonQKJMslg/ElB8dT1OON7BfL3GNLFQ+7qc8SKDCFlGx43Ph0Dh
3wZ7rQKcJUU6Q5IEtV42ZXFm+9bgcZymfl5ifNIkeOAk+YrxG4qwVlMnBQrjc8gD
eakqo0mEv9e6hsc3cv1qGdMfCeYSLN2gvTzOaS3mmyPUDvOb9FFeu1MR62NeNvLe
F7tS418lk+RO1DP+mLvVnxVh4qO06kBFeHO4x5pC8KRsqYSYtoO8gW+afRG3tSJS
4EQJ1dBMXjGqz0rEs2BiqYj/ctBZI8RXvm5crYHhKb4P/STvrAwPUXlh8G6O1ngI
uX7sBscipw6WTjgA+ps+uVKe77dMKRCN3zIGc276C8DATAf0bV27GPtFR635tsJ8
zsYCmBVNx01of0BueiwivZoX0bTdhUZhTuPKgVpxtVLGYk+V4Slkh0sIAgdULVsR
m2+CtQF1GRfqNywMjVFXtITE+15xSi+qlu2DJll372w4I2J6bvZV/6dqzpbK+cQY
VSvHmcycK391oM3u5n7c0nFvsq3GWiswPchI7Xsf0Ax6ynEDpKoy9L4ZqLZ3tlDh
6LD7lq1Ph3KM3JLU9vQTHMqGcPZ2oaq+W3dvYllPyhxLd/CRVatf1YcFnPIGoJpH
0w8pr7v0qKoMmmxWk+VoJRAaQreLjmJiXIoft6+31XtaukoqXVazHEkdI2RpnYik
LAdr4bspdUa5Vkj1uFwqQ4gc2J9+zIwRWsXFY+8wKppG9B3QVPSR5OJNAwpcpzSw
kzzkSVBIn2HbybGyKpuEjTWxi6ilANwXp3BqNSQmb8kiIZebN77lRiacghaZdjPX
Mj6rN+s5znEwurKxUWoDWSOnARzXg6TGI9eM9vYDHyAv3GXRQp37LNVml3wTId7l
xYSmUR4k9ZiJR//njpeAeezm9RYH0fh5KXqDMTda943nQm6d0Jyf2+AETlFIU3Iu
jVbOxI0BCeoZII5m+y3uN/TN0D1r7DOE+EXw36GvPTiViF8cNjIw5w62qVVWGy1/
JNsnMSXj+4flYJbnzC0RrtyTwONBy5mEorTf9ML9AZb1Tfbrcejqi38ivEZABk1B
93RMHhuc9CAv8Ki3GyEmGPhfYuU9DZDTFs6bf4xUdijlpoH5gMFff0vNpkUWJXSa
LmVglxx+ZJu2zi1iV2ElUjInfk3Zzha9hBq19TKyXNQd/c6Hrc9YutsdTie83qPf
w6H9vE2DoxpaTauA+w3d++uSMLPyG1bcM2C+s829+Ra6hvEo14PG0AZkv1wvlPIA
hDsjDIjMFqz8zQYvqlkNtPUt7yDtRVKTqRTjRjTXwQzO3pRYL1xK9N25b5EvVUOx
wYOhrnTysEFUEPOc0JYTeqMrFWHmE5fLHABeAYttIs3NPHEsAYYQHoBYUO8tGcmH
dUEesy50PEV0jWd2in+REFaFxuITvfdBIlnTBEgWgjcvFp2ABTngDJZ+LJHizl25
i2ohKfJTsn8OySpAJbrkkiLTnY7nIeuDtri3uXkgJEdIZgm6ECPDNZquHWT3Ofbo
CEv8VlJv9B73/bfWL3aybpXAqJ3k7VzkRXW8IjVKs+TzIVGoFimh4OPyWjTEYbIB
INoyj5Rp+21IQgUJS0VQxgWp8tUYdwRhi4r8E/ZLPnX+G2vvRS1ryAeq3vNSu2JV
xjnrklUJ2kpf812Fv7P8ddfHUNF6ImDMcHt19J1QdDJs9pV9QFlO1pRVUTt3huuY
7PlcKdXBbPrpUCABEfVqnLin2DAXnevpWdoxIxuEj/GNuO+LC60sLcZ1YkEze/ZA
hR+Y3Iui023DGfiKLrUhNgOEPHuvLd1u5jHdnkV/0KOE5ZtFWuQ9xPCkd7yl5FoW
blbB/t0GMklAo6QcxxzoTwtPt+4nYW5P1I5fFcazzzmTPcFrWaiXssQ41WJXaf8c
Gkn6uAVfpujlnNC2oYBIB+jlMaVXQIYHWPQym97yvh5rFbZp7+pR9jRXqtkYTIPF
aiD55KhTZRDqxOVRVF379IwWU05vJQ3WCRBELcCE7ltkX5wkeLJXX884zAA8Fmrp
McSTeLrN8V7B42obkqrbd2nGWQSThcTCtT/RkTnFXntKyBRSNEgu3hhVHKFG+N+B
xpvvVMbea9+ujdi7N0Ja5smKSZ4mS6NHNQkQfL4LvhNHc4EQBDHWRpS0DwFQ15AT
SyTGo4qa9p1LcYjk48g5zEZgPPnEjlsfXWIfDF2Krv0etwt5vFiYzapCBi+si3ny
BoGLM0UHQVVa6w58aTNK6bAV9OmKIZnI8ME0KwRCSV4NSuM0EE/1lDA8mo4H8+hI
FOAfH5dcfkyVRCLH162SPIIUuuc7gyJ2Iq2x8lKKytesmCQsrdnk9X0uDE9u63an
mZD8Wj7kaAGfOHDX+oiMPJ09Pt0ydmQjoljD9Z/LROj7g9I4XAtswpggj2t0EBSv
WYMvvIr7+hpYo+t0chX+Ky52ftIG8eT0eNrPC8eV3SBKhAUNsYFDBL1nWk0NC3xj
eIGHQsfsqc7Rkw4ucFZQQXj7HsIVW+31+vznDM7ENt2ipnl82Zv95y6Mvb97QF33
upLLQ+dSMrmtwlrAOt9lAV7P+JyFTHQ74sT7x13jV9tkQ/sgsYQwE8NhurVWjr4x
aRrMDqclW8jT0JdisCyZkWtipOOyjIp5UsH0uVFGAKIs1vfCkLS/6o5ZsIzvC64H
nQSWACpT9sB4EHku/guQlmsH5H23ZTUxEQA8TnyU3teJiBspJkgIqJ/LLEl/qM38
MDaO/ucAoqOqPYJ1iBhXTL0MhepwtZNXwHsTDEa8EL5djqISCkTi93JyKNzTX0tC
8ClMiL+iPcywCNtIXmY1hfijiJ9xJZaHx0R6ISrki3XJ1FSCdK5l6ZVzO/T1k3HK
SBosuvvJTuz4Lo5zhHzFtzk+qdUIUCqfagY6z4QxKCCkjrt21VCygrtJf5S+s4G7
ygqYaS6KpotIMJS1WLTQxybEb7z2pne/2Vey8+hdGRuVOBelNRbQPrrQwuPgKaIC
O4f3maMw2a44p1cnB61ymSkcpmNqSd4uvBGXR+IrMBCF1FhaiVziqyONAE1GadCQ
RWDEWuliPbo5a8CxxJ3vibfn9doj6U4nJ0W0TXso5lZxPzX7CZwqP2SRVw/Py9ty
fxkZj+cX6ZmbDaxknS1pzj75S/VSELoBYky66yDkgzeYx/WUfmTS1rpG1O0tI4gX
+pYIntohr+8IAXt+yVxDoSFocjpJ39Si1J6s53KywZiy7OA/LgLYnYAVTstoWLwh
r3EIczS75EzyYuoR14NM4fIBC7GHFXitfuPHEGtkatyCt2AplKIRop2irsllxYYD
tmQj3aFhgVE25dhLp/0cKsf3YL4gJBucJ/+bSYBxtt4jrkj+VNwFv2NDmHTlJAZN
mvH0S5gng8FhJ69zqu96c+5fonlcC13xUD766a+kieRQLGLneAXv32Oaj0S/rFDe
WwJByJq3EdZX+ivt5KvfJR4jV/lGy4V87pbUUZEdYiTazhsSm92N7Ko37ya44TF2
3byRtuo6o/W5lT8aaQF0aGhtMp1FeKjiGyDBpISDpNk24JUIc0Ll5w4BvwJ6zOac
Nmjy33OmsGEgcbINIlc6PkejAeEI8Vzrcg33kcJ07OuzqeqXYLPPub3vGkyte7Qh
+XigaC8jWmx1nhwXa4Il0FSyAVYkB8tE8X/8JsxjKlyVZ5YVBJztCT1UsjUfxEfK
+7bad8xbwDREifaTCy4rTjGc9K99/v2wBXiUrMP+/HS/98cH4yJIc043dn+9DMvb
gufGfKVlaaExkVVwx2YpOJgjG9Fc5JG57EWC+DqV8cD57qxDxWEXqh65UQEO/DWu
4RIkkCEGKpWDdCrMS0TSyEv0GJT8S38f+d/bobn5SgLykAfVItiA8krfPPJXl+yv
GnwIntp7ogVTnXZkVsX04tdiOAX67RJzP2q6S52saBt+og0vce1ppwJPsrKAVdAM
2fSrYyg7y5PIoliUPGkjxFs0j6a369FpTvev/IVs4ZgtkHzLqNqcWEMzwF1AoBHP
I2XYCb4DTttWYHTv6+u5KjwBSMZSwVIjh97d5vyA42gM5PwFgkONe2xebfWp9mr+
hfLK5uIVS6hNGl26xXlASlckhuZ+eIp1qjhHZkkTyRYG+WFB+MRcPdE9JR0KU8+0
BYc5yIsr2m6RlG2FvSqJJxB1nZovrZVg04KUBhYPsQrWYp08WUfz2KUEig1QkNRJ
o5Llgh126u1y6TKgaP2bx5bhzo+qqjgaG7hfOpPN1wkLl2Ni5rQWZQdzMx2NygEE
2lusq5uH7qSii5hZL+aI1Mlk5rFy9XfI3/XNdR/mH0PgIsifPlnS3ua0VGMdrWrh
upQrSIV6u9eSXywRVpjNZIBP+q93HPveci/m0P/Np6rVM54VYv94woO8gXxjpYX7
Kg+eycyOFZH4GTpmnu6/Q2UBbSrj8y6LQsUjdPtxyjozahciVedyQqiHw3vjPSt7
6GnlPn/c4yh/NEuDX3oP+Af+tPqxYExtoORUr6xQ9M/MkW8BCbsmBkVdGwkZThdb
ss1AdgSFVfUOiX1HKfF2iTIZQ8lONGEVb3GDJNjmCQHE8rjbJq9jc2CpsWURCXOj
TP9mnkLq9DgC9EL4A+qYIAnMGaiUaG2k3FxgdX2V/hKk9EGxU7MudsXU4uVlBto4
C38Gc8mC+mBKIiQCxVxa6yDvRQV6sdBk0tcPc/S6KN5f66clTaUxV9T9iobNpaBA
XgHPNyEG/oxQXpirpxAu9FeDqv7sgm1scTeHfOBrfdmuVWuTYWcgs3j67cD9rnZv
S/Fqhp6E0fbwv1QT3tEqpE+dnIVECzdgoAudI/Q7wikGGBKQzw1wTuBeAbkfX8Y7
FSEXTpbrKAntfm43RV6c9GSVavHamvI2WSgIHWySjyEQeLVpf8HPamZvtgpDHoNq
RbdejyS5B1WYiuJDf0AFMl53X0SZp1hRxct1tcu83Q416yLN+x2dTzsvo6UGDKQo
YcOO18LrhVD43xoMOQm8TSiNXHyzpQB4iEgW2w9moMN3T/kqEVRn7pGJcD65bODx
HNTU7VvklLVphXMcnlR0g0iMDLmF3+m7sz+N76ehdqs9U2kQgXowG7RrU42lcf5y
tiM6SM5hgr9xlBShW9esj2vs+MJF9nNVM9UpYrLJANXiwmPZanDs+b4f1J+gWkb1
m3ynC0HPVfwAT//cTTRsPZfJDA1PU3f2/nAdwykS1BBB8h2dhcqXo5BkWnVyuYlE
ofjP+KicnXHAR5LI4EjcHYIXkvE16JL7CKwRbFHPFlXFrzq+E+yjNg1g1g2UjjoW
WNMjBLfzvYzIjWBIfIU+CgvXMof2erGi5SRVjziJLnEzGkbyZeiNJyrVAfK0kzxT
ATnPB9jwZvtutJ3CIt1I9oLcWNtSmMXg3i1FDCPc4ef0RQ5/XEgUTjvoga4yMfuF
rHyvfvjn0xedFzSPYX8MSA4RvXnH2x1PgonOE5R87A78cwO7y0Q1j7SU/Ks8IpmB
NhWMfFMYtWg5MXQQ/aI8ZrJlpfpUn+UezI2pN3ld8PSX/EbbXKcv17ngUjw3iCRO
ZQBf1P6ubK/48gfy4EhI4+O3Lrh3ZZrrnXT8jqKw4ZoqKRWCTeigKVNWQlNjPuGj
Om3HDmgm0Qy4Ab2vfS4kJ4hzJEnieK3TQxSwXvfHbpb953s0sogWn8gwx4wwInNW
FzXvKp5YCU/DpdZ/8Klaz6fv4BlhQaxb6SngkLLtd9t0pbtvA9YWUQZOGFuak2gS
H5Frkepn21DgQDNkNDc4NhfMQHy7J7hEGO+4Zhg0vABfw+3yb9/OiqHD42K/oGk1
JWI2oxJ0XVcvj/Mg8U9NlAwYJY6iRuR6YdWxncezlzlCf+wue+GX8SMBkPNXjSbo
p2S4T4/XVSEqKoh7bUIkY4ygG1TpKOwyuMQ5VhaMJuNSoOLrAGcSSvzPkAl+f+Bl
VhX4iXCPDVuLVne8mVSaT4DZmUWnJcPjVYVrRTHJ3SK8KXQwgcD0v/NhbwG+Q0tz
Poc10lxaKcHJ0dpHqJRWRUNbg69Dh08+W9tNcezUB5hvNuAypDxK4jia0JlrCeDY
xKpEyblR+fcuj8tfTL/dHfB1kORXJlcQB8UK//pV6eRlgo125Mfht22wExejmuHa
2in10XlFzmtEUxRsSyiD3zsOJBpVu8QCHrTDk40fZTOa10O7czEw1snkMhshVUWy
RH7oKA6nnvBzak1LDqvSUHpeS2Id/vSZ20y4GLsd4Wd2028E7Qq/H1PaJVfikm5N
QFRfPjsnMp5j/mfz9TWj07ysHSk5LBNEGKxH0njD/X4fMGcH6YokD/uS/adJRKbO
NC6ApZNsf5SBjU8lhYs/U6c0wcJu9dEsXLu5AYCQJB4u2vev//sMTSgc0zzEEOuN
z28ioWo45IAyJWkuhgXUVryVdxSrrMsRsEbBBEmXmI4YcPkRQDD0PzbZwzhrnh5O
4O5PX+m9woB7RWywFTzPTNwiuegm/giVyZ7Ln8AT+GHvDVq8KA+3gwtCGnswDOIt
mcca7rCcDRJnw8reu/Pfp324nRY3bSwpF/HE/EwBe1OrSxKZcPfT2lLduGUAExWF
ETFmcjK8pZKa4p7vFbT3p+l5tojB5iFGGa9pJTd3sj6QtzABGNTL77MObxoC2QfR
JyO7QA1UQqhPS6G9u+zNzBuhViZFYsI2JnueK34Fq8AMSVrKychD/759O5k8zTyL
Zc4kojuz4qFFneaSkpmHJDgAnYw9P42YlwDHPix3xP3W5NxFEThpjw7NAPxwrrwY
MnorZHGSSqwmctDnomIh3BBAQEqc041yZR9QutjxLq/1Dl0/7/9haraQiaKRN3ts
ZY5yY8Mt/jL45suo6rN6jfIptgsi6ZfF/uL7J7oS9h/PPnhoMuJbjffi+2jxrKG+
IDDXo48alSCDGLZZ17z6eJ7VN2Edu1DaT9lAzCepiPfYKh/gwnOhEu+nmcKBqbWl
CsHSj8rIoX9AxWPM4yBEoDg5CQoLKdaLYqtNNuF9CWIocjTKvXmwZY91if+yueR5
7UfjdVmns9vddedy8dhgLeH9m68/lM2kei42i6SPWrWNtS91yFEuL4Wuqxxe8W5Q
lf4GrIjXq03eST7T4dmyD6Cveo8cSgFbYLBy6Vkdn4Pwov5qVjSGdlDswGgJV6LL
kQS1nrhOnmstZ01DhG0QH27ythAGmZitSMolCDG2r+CvB6GPRXxjKsfy7o/zx5oX
6JEic6EtkJZv6BS4edJMvxafyNlCjdqU6stSgMMuXMS8qw2AGOpMDX+hI8fJq6g2
HKd7MIL+h71l83Dlt5CeTHLl2LpbndrjIafwtoIDsN7I9rkoe8shN+4lInlTA26S
bqHPSHm40z5nk0CX7lWTOfmT81cgXhdx8UfG7C+Hq1VyzKoJNqyvK5JkEPpuW23c
IKiJv2hqzGTbQ6p47gY9r1JFbiOoAu3K30tmPBOt4ON/Cw3GU17PMQuHYYiCS3eE
vEkQXMRCVP16DP8NZcxDve204UjeU9U4M2k03eMnfW6CIl2wfclM2p8HckhcpDFI
brpv22XpdDdjsULRe5miLjlqX2LWlzdn4pL1UVo84xIQXMVmgeMTiJPkuO3O4WI6
sKYb7Ya4mEVvl6/NyMmfa1n417A/U2dCe5Srv+2oH/VNnD/jbJ/CAaEUDvIh3LF4
5HZY9ExvuqIchvZfYUlrIEQmMh2sUzP5iZZC2He8kbLi7Dcw/UqcEdqOQNyJENy5
/cwm99xr5nw9FHcPgFOs2gU9E14+8VU4CWyCA4BdnEeN5GNEDFecsRINIxCzbGVq
r2txIPhPXTwYtTmAQyjlHqBJf+s4qQH5IjCKyACjTaHTqc1igwQ3viSz5KxMGIJ6
AARgeHLcXA743HJHuykPCZ4NLj9+BqptznFTnIUQCccPPxplIbCOP2u1m2ThNBoq
ICll9I+2OxU0AGd4OcdMxy7nyZYEwhISH5BLP5o+8876vHi9Bc7GNIEah/xvGWaQ
iK9BxThhgD1zdrInVYJ/P7NqxiDfuxnOca4LGpYiEuW0w4o/F/3bNvR8DSK20SbM
bK/Fa3a6RA+MVqw40ITYNJnisoVfjg2jb3DBz7YImoBGkNLA2zLBUAAASO19zelZ
CqrQqxyqwNxAkXR+Pf5vz4GO87jR7dD6tuieq6FxYZAguHCPwzKZevnTJes8R1ze
xyEq1kPMkqGDKAw6IbfzWk5hy9TZuHOM87+K2osDRJ0wHSq4vcFCMZQCbjcTRz3h
Pw7bJrohCulEnuxDaR99+NDStiYUjbqkPpiAMHOQTlfunBEqFF5hetN1o8nzQzK1
thIYT4zGcBwFpcUHgw/J8DRNAeUxd8J2CbEIEpco+lRi6agJtDCWLznfIHsYc3fX
8/OOlsvp9J2Iidn/clA7uCzqPzk1zPFq2CoyKyPi0pj7AYnqmCIM6x5MsxVU5plW
G/QiqFE4olCtq5b+f/j/3GOOYwsRQ33n0586SjqoIvhVHAW4Q1Nzk9IRTda8G1DQ
DSpnoTk1ylZI2gICzFgQ4o3e5fuoocU0Sd+W8HHNqhsnJvu1iTTDZ7M+8I+VAH/k
YDJNhPtjCsuhV2SIDsXyXlkxoHtL8/2qWsRJg1IRZtY3Syc9SJImGvT6enXGiFKc
/lOQZPvT9wlq+YEz1mCl3fe2lF8AKKzxRlWwUDDvi9g5TEkvkEcrcN7WZ+n5aJ35
dCpM0sNvMjaXtB3cw7jfFJcNrPzAbbs19u5tzXyloNJ4xIvTZR4HGaHccSCYViEr
LtHgbve/jr4y96g14ZGU8v/q3YTLjn0BVZzRU6QiWEAcweGJ7nk+Ndz/O4Q2HQOe
kwBFSHMnt9uBtB5C/itGtBkoZEYUy1Lrsy6S7aEt3N0zeSj48ssoc4ATE8gTiGGw
0mVWOgbStZsMSOqfVEy2+TADPkJSI51/PYZeG/QYD6d3jjDnqN1Z6djtI9mundrG
hkMCbr7S87wDnOvh5o3Z3oTORLvwAtXRAdFMjYvRJA+bElLtDu/+E00edJ2qtXMn
Zm2cuSorlTP/Y9OaIruSjL51JIDIZPe0PDOAaAj6ss9wLKfvayneYP7gf333k/TW
tP+f41sBUYyKHTteYC7jLLWki2HCcQ5V+N0AH/iqKbPHzQSjh0EgLv/gNAT1Y77Y
KX2cQZUoFUIlRNpcw8okpiUYtocVAMcUFRKNsMQLIWzstUoSzXJsLfxnGwA/VRbJ
EAZjuljVeBTFGiVP55eBkBE31clBgPPKrsyqNEkOOkW4iTOJgWC0OY/PKN8yuBcU
Tt8ygo/9lhsARDdFzhgq1XytYQMQcCAwsg5wIowqjd6bLqJmcVv4Wx9i2dCnp2IT
Kj/c6MJmFwncVZWsS+fFedlhcxBAQF3EpaPEJCoe5BXq7dEmq8Wt/Tzv+LsxZQoy
udZSY53YAg//74rpHgzdrOOyGPcfeYq5cnKkjjGcH3hjG8rvbMmkWwFqKZzwSlQf
KtfRTHP//hpjeLOtt3uL/9W7tGkyfSK99EG1ijBOfbfMxA9lYoC1dIMrF6+WGWf5
3ivC8Us56XC0Y3lRnDyexRe6HKGDXbiuLkQEaeouTG5w4j4dmpcz5vdf9HNjDm8k
kiw7KhQZmzeOblSSkWv5R/Df/+FhgZy+HdXZCPu+7t00VOC6PtP9GPrfA9rwY+GY
DN9XEaiTEMLhm1Arc3WpxWit7jgGCTMHhBQc/HGAMwdOs0o/eIVcKhRAZFvn92UZ
VU0jQrffY481vz1sexHAoVsPZ/9tcEpc/Uae03yVjSg+UQgvorfmZrob1nAuJfN7
FXXMVEm8x0NRvAi+7aFA7kLlCQb7qJUHlUf2GIXOt/Ojzi+hz0iwfaxhTUi932ZO
ir6l8tJX5/yvbMUovQ9ihxA0x4qfJEge92v7VIh6WL7qXjnIOgLmTv95jB0wkPgh
aj3xTB21snoeOH2y6BeY9eWGfMhA8Ht4Opz8rnG/7YkA0qAl/C++dPDVKGCOYd/A
Kv8KAU4CyOlQajDgkdYORSy/eVaNTaC3JVs1FsRCdQ/VohVuLrpH6EDuuWgkagOj
c0uu43M+iZCholzU1mTNFf4asyAthcYHUVLGtzV95NRzwj/OoCVDHhXjwHyTfT+a
BjK2kabeI/t0rp2jVGH9kNce5AxaCwgo7buSTHVprRN+aelAtHj1Fk0r19Rdpe3p
jVlOLqAhwpdceqsYBXFfGOL/dW8PDLYvxjiCW+WAwQY6RMjIdrpR4HQjO6+VBGe6
lzB8lRid+t14lhU37h2RMSC1a6iv7qeehEOCq88TxXTubk74ZHl+ZEsLCwJux7+l
CPCGqTLvmmTSxVwG2m7VM5dGa5QQwUYDtmfQorxORb2QChPVtq4g4z2R/Ex0k1Qs
UzzuMfLomqJcPOwarB1R5AnebfBuIUng8aF0sj1Quj8rPWs7EZSYKl6rNrqqGDwA
gMkJFSta8y7q+7oDUU8RKFbaHOoXjZFnECn1/eyg+hapYqAAGfIA9EtNAZJ6hDxC
Oehnm+dqJETPgc6xc/9RlY2IqYUPrpILBgaeyahMi4uG7lUgxE/rBa6cPQGXSyQB
xX5/4ji3AYmrAJRVVDrIZ/PYYSqmmri5niWivqLLqSpScwOY4IX1U/Sz8Z51KZCg
mtnvvhZ1wuokDY1+ypYFpJfXNW2/GhgawdGhkwY3GJZU/MZ8U+dbVgTb8/OuIaIs
v98UBedRcJfbhp4lnudwvuKtR8HavQCzCyFgGHehF48hPlrzhmjHSb7YSX8oCB0n
lCEvnaOZ9RB4kH8SaCpLbzaD6BIbYT6BqqwCayrX+nh3IPpvic8iaShD7QRMT/T7
xn7RnmcPCh6JaogaAm8QXFUkbaWjEQ+vJ605evKKBYdda8AiRn7bNrdLz5zGKp5c
gYpc5l8yjuOSRG2oh4dmsQfKEJKTs3yDU3SqQ9JxZeaFlNVrPNay7vFUAyr3imnx
j16E5PiBWTpFEDemnDs3WXsAbwIfMBdygDAFvUzEGPNX9tRhKL4UeBRhoaOLITQX
yqWPUFELOQbTYpP9jzGxOARkjCE9EAq6Ky3iNvrHoUjrLj+QL79HMladXsnhe8uw
nR8OuJyfYx8F1rkf3Ef2ft4UuIW4nMNTtKCXcIaqYmB1tv/a//44iDmCUuO3mwMo
bmSU0uzQAsgHCyvfmsR/6buY+eD2LkfO2kW/KAw1Pob4PRkTG1bjQcgJ2agMVTEL
MulqzbqnGtu9dCCz29Jpal+8xRHuYqX3Ud+57nfpv+7m62BqcMYZgo/SjyA2FAUI
H/S3p1Xj06jzGnrMHR07vDNKW4iUHXtHoIsW0pfdIGX2rNuFBk6cpjUz2/k1/RyW
qBWVd4hUx+gFgrkPlhiug+lGoMVwQnTTcVTGW2cSg4mBqCoCPrEyvpYYdQWSLZSD
rBNbLftk4LWc0Hyng+ymXJixvp/O0ZIUUZ+1dPPZI4CxX3QEUMO9BpqT7EOWJnIc
YXzzYla8orwuTNzP9nBH1oRXEwzINSCRrwBM3dh+0ezYk+CfxwIP5IKfCwDDaJod
pGjaS/XBpAwpj9UWQ9IlEMjJxKV4ck3sqIxRVKB6koIHetYMAgRtlQ0dOIDL0GMH
R7jnFuJXHu6JN6JNizSj6mNeTAD/UYEnmbVaqEt55aKUmnLiBKIkwN+F/fbKEgmD
LBvqbAZUbOsq+AFI1768Ye+zX3hcAFynRugt6XrngQaS8Ry+snk0vFVuT1W3AeYl
NgruQY+bdADCC0xc51dlpQ==
`protect end_protected