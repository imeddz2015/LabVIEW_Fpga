`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 16512 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/9huKRhRMtvnNqb3Z+UU7TahEoHV+T8U3P3ufru7l1O
3DlgtZzb9QxCbOjthp9+wDkjygH0eUfDrEl1ovhZG62feDui6BbypB9cxVtcPU2P
ikbyy7xDFtUiJL3dyyG1Ebj40RaEPwOrkR0iFptjEvqXFwmWmNw1Apef0nQ8MwcA
dVDrAGQzArFtTGqtbNudbJQWBlG2fsJfKMaUS5chBzHDp7HVNa19u5Y4aizdvDfb
S+bp9gGn3uN7q7jcfH0csN7LPYvJH5lE/Wn5DCyG51Dezl6UMompxgdGIHQLWys1
+nHHyr8mmILPub4QZwgTIenCgdFtKYDeOFazdZdwV+HM02Af5gCemcxMN4mDpYFF
F9X8R66xH0PmIIXDj5/lnrfE9u9R82Ynz/8yYagmuULCbC28jf5e3DmUXmi/jKFR
9XXT5ssdzqWvXGgrY15b8Gvvu3drIXNHpFfTRp2Yq4Uei1PSaCdZobw4vZnvgz8M
O7wsjR1jNRbBKTwewiNgQO8o1kq4PlRgZ+kT5Ui7CdbBlNqlzPu08ys+rKIImtno
M0VVZwNpO/aDtjsVhhrnX95b4twFmC3ztYUrghlIk0u3aMyNxABbgAY6w34pN5j0
JoLotkl7zHxsszG7BGkxSA1vYDNttDkhaTYvwZTxUM1H8RrH1qxhs5ENjUJER9P4
nPqpN98r1z5o8osaiJ9rlNauRim9L0LneYZiuBEFdV5wRvKDvjHj4JCbNNtnPb4O
M9NoWxBDwDbPqTN80u9d/vWTaoY0VHOQpCJJfl2y+5jKs/7MYNJ7QU7S7mwZK48x
MtGQcffUDeP7+ofjtZamag9RLGjuNalvmAYNBtLsmpMW+kgDVGlqbBQuUDN7fte0
MGz9YsXBahPQnIyt8W4uc+UUC3IY8ha7zxBcZ2jHXzNTg/STyjW7i0ncxVuIZ9p4
ydNCkholZJX5I8akh1k7j9OzVmO/7NlXGxuGJcQusi6QRhV4Uxkil0e5t194Z9ZJ
VyUwqPDPPR/HLslRiVxCNU9h7a3w5LCFnSoI5JbxfZE9UJvT4cTAQibKG3E7Crj8
gjP0WeHTKefmPWT7HfgnqdMTIOcSkRpByrZLr4VRb+rph5hJU3+0Dr4oeCjSwzJ6
DOBQ/AO7vEx16qQECAE4pD12WgPIn81xJgGL/VDwSYikfNvJNAmbUm4mfyM51ev5
vjpYkcFqbWhq8dR55Ls11wnX42bqY0DaawT+yP3Pim5XWUnIQaP/PJ8/YinDVuiH
WGzESMuzKLPCJR6UQ8dMOFssvY2UZFogLj5AYfm49YEkVPwi7gjoEHZYD/brF9yh
6iklBHvmuchNlfWTsHsDmaEW5e9Y1gaPQw6NdiKEXXs1Dl9rTCBQEf3nXBiAbrPW
iqRGCpteLk2BIyLtwfDZut/WsBKyAGoED6oJdTfD38ukgwfGGRI6XMjL+75UtqL8
eccT8p3VnVElqR0YFXwhislFbktCS2D9CUkDCMAn43M2002mm0FuAXawiE0JGw/u
teyG4taURPZboUn18wb7BhxlLfJOAPMPymKZ4uzlYVjoCP61LUb55UucVwOzyJj9
GZYKu/aGyq5wunwbknnxbdAVgNUBYHJcyWYx3zvyyb+p4J5kSvVo51hc47n3/lb8
y5kAneTn28Y0b05iYBPzNfUcHNuvi5M887fK4R7OmrxfKXXYwxHzVSCVE8ajmS0C
kovUa2YtdDEzEbh3SvRj4pIUNqMifsXX4LQVnOG+ZfuLG04AdHQBm1Fw5OTq0cMd
y0qVZIWrQEqFif67+VRrPqxtY8+5MwG43H018u3l4ASyu7VY9NQtaszkBHQ6z+/m
dAvr0yd0294NI5gp9uAhMY90RmGo8EagnPvQ7uoXewkv0/J4vgwuIfR2OCgNaAfC
M6id+YivZl41MR2RhAWOCaJgGKqz9Budmgqmt1y+QA+ErhmnGSzd/NxsStDXuCLN
qcKh23faVbQG+RTm0QIyoR5vP8LPhzBJo3R34kKu7tuzeu+CkohWgglAZTrqtKvi
G7ywwlfr0B7u0jVRKORVGPJDN+/Lcz3veDsLl3Z5tVfaR1vwo2urJ9r6lTWezMj9
yB5Tb1/0qhuL4WpKk71TPb8P16D8JPF1EEzDYCdWxA8xT14NhI53Q52fRVIhOGqt
6X79U5FPyU9z+lOjguJlNlZ3biJtyrbaCTZ5vAuaNPNzalJIJjae9jaRRFoVfvjz
4gP9O6buZa5rkt4Olk2IllX7nQWWYXOszh34OvV0b3aFfTtB3KVKrOzIqOQiXQN+
U7KQRCqk4+huA57Izb1jpJAavwhw4FN01x8b2C7oofvsX8atM9QgndF2OYXhGO4W
x5FeF8foTl2wk/JE6ktqMQ2Io+4Xh375cUPpASNxp/3/e5KJJOwv8vobyZdgh9cf
6QtHKqxDCHhzXbxh5ALM4RWH1VybbXTEMacqR/Yvczx10uem70X8bsXvhYj2PXqt
CKg6t5y0sDNzcmhHp8BW3GVgtakp3xsn8G9ITGH4Xbssa0zbQUJOQ3y1sE21LsMN
hZVILLaUF47jLJVXAxoIQplhvRt1N4XT56F7q/AXwQy883EpgIiilctUWc2LQ5uT
O5xxFRgmPDtydVIlgBQYoSbFNv5qZyp0LH6SmAJxqiNH+iRmNxqdSE+wynCFZDEV
UC3CpISgEDrZKbiEqC9XIxX1TdHCBE487kdLfT5TKxX5a1I8DeZUXRZj73Zn/DA9
TnEqpXCjZBroFlMxszUsNhh2yh1b8AwCzzizBbb5qwi2FcgV8j2vkMd9GbG2ZDQ3
yL0vgyGTVM2kS9fOiNIy5+qcXZArmutmwDBkGFrZ4PyTZzx2m62gA9eUMlNPFwgG
AQ22mBb1ygSUwm0KOQAECl/gUxcLRHkaJIC1/ZU/MBO0+BOiipKe+KXTvefrKyB3
7ha14Yeeb04IvgL+40Dgry/FOd7mmzJveMeIIIvJGQiGid1aI/NkMSSv+Muq+vGu
pLrobNc99ePdY0PegQc54jipDmCRXpBcZ7Z5AgPgOmGDxmFoK27d4MSFa6M3PMXb
B9TK6oQNMHV9+WrMcISnPGlMpdjLb4/KOv3R8sGpXQLDGutDOJfYY8+tcLhq23S7
1ouWgVHUMMCjKWUwXRxW9Vd9ui7mPRzqZ5uy44FXVgf0xKIwmjCFWwvXyHHuUMIf
ohPNCgZ6zWg5HL/939lEMmiLO2VEgIMdgbzhiYzwydWYfhD8Np/LY+mxqBUCq90U
inxjvoTKCeanNaxF0CUcuoFjDkaEyP4OzTgl3P/M3zFy/dNS+Ip6zvvNyIly57XX
5CTT8gGS/YuB4MLid4tVHzjrcCz2FubGc844Pnq/pQA/J6KE2I7ajsMZ76ym34hO
wZHIvxmVbjs+wKyZnFalpKZR+dNR+ouECjjEIIuXFHtdkzIUo2p6q6SVz681amCM
YoLRbyHTTbvoxqqnIbO/GHBPleD+m3bxiEs7+lBgPikobeOPSHLTM3hA3yshY9n2
d+2WBsA4nrDpAGpcyw885QmbkQNIedq2/BIp1hnBWDjIR0MtM73jJlhkbFb5a9AZ
dv9XhinhvPDZTYjqZAJGdk8Gg//uaY5OQ3MSMxXax+ge0NMqyky9TdZ+KaFr1r0M
sAsgshaSTvDreALUTmczhIsVoJlxRnWbheG3jCyiRrFWlx2p7zk6J59AXWxXIU6D
wzFNTa/TZ3xcUl/KN0fxtP5xyAjykRf3Uv4OPPyKZIpt2KDyM+PdesU76CL6VVXT
dJPhFtamgto0ofsAfLfeC68vnqE0VNmlHqiDg+iVV0SmE2iq1OIiCrCWYq4/J6km
Tf9+Nou0JSunRWfXRu3VCR+a//XULYDsMSv9vCoLscQpvoxP4HUF6HbYkuWHDmKL
6P2CV/X6VPmDcacY0MdHnvjjBEx4xzb1l0Y1O7sC5ZlvT6u8A7LiZaThpkroDKIv
f0ZTD5BFyPxxDv9uaK1sQMrQqpbCwwJJL/VCrfhe1XJe4WSM9ziWmA4Eo7eokQ54
eFnNqulvn2ZAnJl8S82RXj4j99vwM8eIa3bR1sENWwxzoHdLrqdueSqEPZPYHgr5
yAiXSK3Hi8wdNg2KkYZmJSwRUmKynkWkTgWlXZtPC/n3R12DaG2YwLNM0UJrZHC8
plqa77ckS40wmb+MxmMi35URPF9n4Z8A47kwWgQfISAQvje2CNcPpjh0F9Kiq7nZ
NvInZpFPNULuRQ/Yns13mzHL5zX958WYoY/PANxvKGJAFQcIHztCypFrbaqmtfU/
Q6mHQZXPmfmbpb0fpLhunyvpKZeHi0UhFM3lVqu4eGBMHUDLEwgCG0eOawubUmjb
Ue8dkrkvoafIUvqTRhZbW2yagBpGchDLPTWNng1G1707kunqBF3cz2FXc3zQV9hh
9+HxpP1+yUfykDRATSO8ek9OzXOaScR00nEZcP920d5Zmq+q/tlXjjInQbe+a4xX
fNsFCqOP6crG8g+dY79nFndfA+MowjHuxAfI2DfVZxeBhAe3S6ditmE4Jb5a81V8
ZSIgNpFmoHu1S2c1Ga5AMzElNiUiUXFzCWF7txMv5ZlRo88ILU8jvaxky5e2hhNK
xDJ1L3mlLFhAl4fkm2H5hxwWtC0rAxEQlnub2XDsH73y18FFEBeXpa1NaCflZ7dK
aSfbmUfr6Kc0i6mzFZzHGI/Bq8nqav2RacU+/d8NbNKGHFnnKbgI2/6ddv++ChzB
qGbCtH52ErVzebDN05MJMBMliDV9Ijeef/zzMntNJV2otJ1gkLRvJHBKrjEFunXu
ILZPYoIc35WfJYS5s68PqZW9GPO7hHnu+1V5IflEEYI8HHkodRV+PrTqc0B5Fa2I
Vp0ErLdTh4xJCxQEBnPygW152cOWhJv6C6uVkf5WB7K85cTkBKzIZzYiXF5Wnpr7
Ob9yY3CEq1g7B4txXmxidiM/1aJlaFZmlyFI0vVzKmxPi9yo6a9wR9hwsA/eO0iB
9EX2VcGJ59MtiinzwNQhLk7dhKH/etYcQURCv0H453Ceyy4p1CLWxu7tqUm9SIaq
ZHgQj2L26aF6/RY9WLaAKt5gK0OJEkogwcm/3sOFMPfmCMkAIuK6PpvihzvQ+909
XKMCY0wANhvF4vg41+j1pOQqdEcePzgbj8NK86jJu5lBD2X5TkFP1rWTOh8CMcsr
SyC+NP/nFfedgNUDa/loyEk8OiPYDfnak6l30KLFxS2a84cEZ9/Jf6c81fApLGKl
kKU0/eV9FVdJJBdNSgVxj7muxOx7RU5gRCgHVTsTkc7W8XAUowyx18SPuQjWBtRi
9la5zyVVUNcVWZh/8kHFkNTA9+j0ZtXEu+fDt+GHId580iPRcid+t2/E5fPbIbrd
chS9YFmi7vsce0Re8N5bcXB05lx6dba1raKbiFcEVdf2g76xFIVHW4CCWujoxMbu
TI71OMzvInvHeST9Yf95hL5QJ1fgOtuVqhw4FnY+H5wjm6N1b1lvlpUoK/PxxTJ0
iXppuZOxGmTVQR0gjLbuxkWSdln//qyLML/Wotv4oDbOZG7rSqqtk1wCTfj4f+KZ
JFfV8T3GghScYYBX6Z3OXlMXbLTtaGe97eGQauU3kdH461tg/+6j9m6f044sG/qM
yWz7aVm/4rlqbOq/AnholDyq8b0Ha/chV0BlbHqQ6TnJh5K4420DekXAuaP6DhQp
Zv/abVlXEmLRTHYxTtLKQ0FYhdpqAkxQIC1MgY7TvNcXKocnn85tNhqPiWV0/IQZ
UAZ5iuSA6AbYzi2F8gMm5TYHOL1xAnHH8N7YpoQMJgWVB1Uhp+KCYiIE9OALtjNm
H2N9XIFdyZrVM1yboKfLILC+Mz41YHjUX/59jCQ61HzSf8vJupkVhXW4XmzuElY+
fPoW1JwHkwIKlIncy7p9HURI+VuDSiZFM0Ltb14MqtR58uvwE0kkI2RimMa9Y2gj
GLjh5UUpPtN5CrRcBAEKPNDPXdoM1hA9euv1DwAY/8vXfKtqRahDVZB0MGSeU/Bg
PvDsBy+89ZcyMEusu0fR/KLvzmKfQIJO8HQKIfRXhHBGMxTLOI/k5JGc5J4zaLib
tNOVgNwJxGRKW9GozdT9/oAZqEqot3YahI3lJaOALzpxFSFVcVaoeNMMnGA44/bJ
hNxRCDJP9NkDnUOVZ0s2CtFzY2wrd2PowCQCEOXZSJrJgA8tG4OnbJIyibYKqKgw
FbYvzWtSCBtdqCRSKHgNaXyikxz/8z1iBhve/gmpxr0o0vf9WSD7xS5jj+VJHj2z
LB49g1nPuFfpTv4x5MxWsNyYk2N3y/0MJ88aOgZ7fkYlzxumBLiw5LT1J9lAkuMA
yBszXPIpr3vAx19zy0PhVjb6bh1oFNDTqoFHVgsRqXcme91fjPQ7aGrJUcmSf65T
3cs/7i2G2l+lGXrCQnRPQ7N73nw1GVdBvMwOB7mDcXpSR/MDwMSo87DSvTf2Ttqa
CBMclARg0XQLg/096jn+k2ppF0t2CQyo20fSZW4Y0Hfv/6jnUGCvMfDfWrpDmZI6
MkWL82zjykMPMWYTg/0m58KEuPg7nMC0Ci1KBIeLXolSzSLT56pdrjRlj4NrAHzZ
9YPjb/IYxCzb2C06y02MxL35MeKf4xiI0WqDIuBec5yD3lYrBHNkb4cRnTEqsS+k
Zcar+S5OJzSwURDud4DWeQfruvB2NKL0ckqoLUmUx+lOt/flralMt8HwZpe9mK+V
bsAA/KUamfPGvDwTE7SD4u0g+0Qb5mnEW9HGjvi6K5/aUHRgA8FJBA2js/wtwyr3
ZuRhNiBO6B2lpJRWQMSbMIXz/KsQXfbA2vM+pnrN3V070mt14zLFbWSysMyI7w19
Y5sftjUG1ZsvYSgNIYXQw77a5WQ8/XXKXRQkQJRJOL8FzjoZs/P8KEyJKKGRfJAK
TPf8a+/S3njOX9KiN43MpBhisn5+V/8BsL07fiyzwvXuv7L7TWUWRSRxKcPax72v
j2SThQItP9xv/yS4I28E7WQPFd4XYRcBrmUxvymrCjoLIuu8YT0zNkrvkVLOGEYu
D8MxsynA9kC6xQYGVkJu6stZUpEwVidoaCxRtJf/KtDvb2xtWVGs1ShW7+luu3Vn
HiYGjK3f/mnvd345IzXKj4ewbncRb6+Oz+zgfAY2gOXPL0FjYIkJIzV879xgPXwm
4MzaSeaJjWfK9AWIdLIR0nuo6Fk2xU63sfNJk+LjuiqFxSkiojaZldW5I9brIbFI
Si5Wzhmq4PaxJFIKxcjWAcMDRM4/uHw7KVNx18QsNIR+SzEkWj5YQvInLsNr8Xxq
IrYWnIQuqQmTysH56tyQkShS3UBPlrjK3f062oHPJ+E0dqdzSOR10KyWc4GkdQjX
3ZMOKE68WN/mlqGxCulnyBrgPY7O6K//nJVq/UcZMRfjCsDuUYoKx/EnuOqVJtsr
Z7jW9sAwqb/590RRM6eIZy25SVL4+NPJ4al66EZuFmnMlASqdPe1YpCTt3/OX4RT
TsrPjlGsyW4qLHdA+6cakslwPhYQGguKVpS/agpZvr9ZSfD3XrBCMx37rbnuluE3
dV8yxPaWGdvLCCDsF3f91/L3Z9oGP2RyoKVD23ouC7pgqJpaP+4C9aWBHnVIGIF9
UrFpzNj09hTszJJdYdp26nhTPfGn5WVvkjiz190IFCxfDCToOOtt0uFZ8X3Vf6Sy
MbU1f1S3e1VpgF0rmN9LRvkV1h0icJ5aMQ+LBWlPKDfcWDxA/irtTFBKfouhQfy+
+9SZqAoARbcg/vlLcs+LAC5CFGIoEgm8i/H5LyN/Ml7G4ocVmwHJ1fxR6DvQiRqg
BWHSrqu4CCKSxsgZtVyXuSY3fadidl36fmnO6h/15LdGfuX5wsNcvsZOG2dquSu+
AydhvPMVFb7m1+ZtjQfXwPMpAyxhbB56+vf6219wtmerzIl02EJXIkc0nKjNnO1v
1F0T53LNsHbuYhqEwpUNnNim40FveGhKgOec3egFgSYxtk2adFKw3JoJXqYXTtAh
G+dD0ZdghebwhY3KPogAEcNNrTp3zh4p0zCe9G0PuYGlEKacC6eC2jmt+eTyDH6W
/qwk2T6zQvyNHL6bPde3ty1C8OmgNtwiL4R1rSVfjsMprP3vE3qJW/awtT8OXutm
9kXKh1ZzfOYdnfdv3leCmsZOmuRGJi+92L19AaphFVt5qdSYBOsD+pE9VdJYQoNT
oAxpKX55mNMKfftMwqTEzCtpwHozx+UNILpq/aNdWj3b5vLLpgJz//6gErl3NrXh
lJ3/QAzIpnRItSxGFg75JyGC30op5Pk2l21C+a0MscanTOVyCqLQPsfB9uYZYgkz
GIW4P6w+Cby1SiCQ4WvDDq9YBb2O4EGFL3GKCLAmkQHcTkpdTAdTZIgy0YuVVU4g
Q6DuwyyG/LDdeEW+4U1Z5zeJcTOaj30PbCq2FL9uzNC9pVFg+9VQViE+PFc8gqWl
FtUJL+m4chCkxY9EXZvw2zR+YBkrmHs05R1lklWN8hjaBj8OIC0VhJfXu3uL4rEx
+/vs4F9J1V1tbI9BgtP0EIkzW0XljifB9nreRPBmIkr0RmszjgXU1dfHIH8Oewij
2I/uuVtK2x9NtLZUjEz50h3HpnPQASYNWIKtchKltpM8N/g4h7XELydQpf/5LwP3
nSAMdA1BVRE+6LXvzBpzsjgJFfqpLvcbheO3WlH3r8yJt12trEuGhYCJxQ75ZzBU
jHKCzSNyJ6mADbDYxE0OF5ML6C7/PBMZgj+/1j49ODyoF0gbZ6fvi5Lu6Ezq0XcR
ALPXkIvKXwZwx1oe/J9dZKCZzD9cmqfINo94IssrqLTVYMfZX+oHtTRqrNHdJ5Vz
a2cq1Fy0nVqL4ZCaXA8nFuCpErRGIOdEJtvXGR5fOooGKLRFpssL8OQNHuf79ibu
cQIyDN6qAlxRY2zB9OFhu9kSRn26OFrVRoIQMz7LdmR26ySi5gZr+OWfE6jpL+xg
X56vvnljiiTgs24gzO4etCnFQckWJ/AHPNlD0bwI4uo0i1UOgPOeO3vhmndoQoEQ
p9FoB7eEbnOLvEderxlzRv8YP7IE5SPlWEwcxIUBIWfo1+oQlie1l12gH36cFW+x
VHVJdD/WeYR57VMFW9NoSl3a8khEip1RZNtR36ivaKP+7/J7XkZsHwAzhdaed8MX
pw7hs+T+z4sBGvTgixK2LyGRmfZ1oCvKgWgUUfNCP/0XUEhM+MkrbsuRga812m0N
BNbVVw+DeArwzr6+E0RKPrUVifRIIJKHlP9smLgdhXN4QTbDlRBnV7Vl5vEPCrra
wESBSuwULm08hHQtBBvUNt4vbB73V+r6NVZBnSgF0WWgnS6D9jrqACS2OI+LXhzO
oojk51PV/9698p+8sTpv72lA0V9U5RdESt9fzn9KlczS+892NAVqXx5fHaCt7CHi
ZHrkshoRJLBi0E15Vo7yZ2tdrGFLG3mgJb/Xlu9QBAxI3mOVothkSgFPvgvTB1km
QqXGL4IasxLV5e2IqVqnlO3otfxPI7Uqdjr8BNJiuxfrHiJa0Cv5LRsuGsxCPf4d
4u0M0s0RycTuVDws0VpHPkasIa8iws0xm5hVlC/CW0a52Lb/Om2mNwwLb6ya0i0b
yIoymT/yq1wep6uVgvec9Ov8BgIlf+8tMWlmQMfdSFNAsg+MWuqwBuUNVPga5KxC
qe8hB04sktIa+q+RGFLDP+t2CtNIRasYe/FLL2AE/iMWVaNTjyKad+fwQG0xJPof
zOsqF+zxs7qedYb8g5iIwvjfN45HXfc50rJpCTbJW73OsZpeFwlJrMwsM8rWVex3
P1Lkx9s2Xn1SsQ1EpH/c8bYBeBF/RdEtBk4U3RZajkdOKruUwUbgJVMIFIAsgDwc
W8GyeVKDZKqKUt6fkpM9/zCLulOAmSdmZesiDl9E9syFASBe7SINRq03xWY93PBv
wZCTS2pnoWZiGa7piubsviYDWRlatUISPk71rQHwM+Rn3Fq2Z9IYiDb04agc8+Ns
CP1lKxV4Fu+Byss+4J2jzXi673fGY76RTAO0zQqHPuaPhK/PHxk2929uZWUoWtkU
STlK1WBLXhZ3ktEAGzHiAnEDGbyYY1VFMlNpQrVkEBqdoXOCPHbimMrtjvaw1n5D
T5P50BsGWZSHH/YbQAefC+pPXpIQOux4efo3Of/sWvh0fyreYahaekmDQVWqFG0n
6oLJyjkWNIrPsPWs6YiRUQ062xgyD1oIk4fsmMPgR5wnpUM7I8v6YhRaRaui46tE
ibLLrh+omTV5DrjZwaegD/hHaPhWMLeuQRA6VKAavq07KODJdU+rOAwXNB/qHz0C
hw+gVmSSOkDG9NO6QMNxBoeuqfL5wKAZRZB152KRqNqVNwpMrU/ABrvlV2ztVwmX
mehU829tM6GQHVzxcmbzxSUwyg2OTU/VnZ/CAk9RpNpmJLWV9VnuToYjXMhgGapg
uyFtp52L2OHq2LLa6cEeMWsnqYbatQ+wzzGi862gdLLZvrUXCHaZiOsdLKeiiLHb
4PqGbatfNAS+uUTc49EP0udt4WlG28DeWnMOeevrq7cQCMCh4eEmWjykEA6I2WKf
x+2zRo8fU992/u5M17dvmeerAx2w09hvPfEnLibbRm7KewpsiS6HfGVOgICyNOBC
j6qw01P0lQGivALP65QeqReg+XgY0BwYpPCKlLt/+PgROIJOC5vIK5nKfIQDMi9i
aiSx9DV8f+el45HqioRb5HV5er2uBU2NTQJZPyzxLhK3CGnqMyFfmQJ34XaiYEJG
2S6+lSvM1cvq0yiSA3K6Bvdg2zCJexvJcr+wR8/C3u6OaND3yH2hZ3tJoHrlrQWu
r3QgqTiDrPrzfpit1texxVKmo5FnnOtFDMFBFwJytSlL9X4ekGIs+9qT6AZ8aP8Y
7SxIHKt3UV+MXAzIhDf3gYdf9NcHYd+SRagktU1DXHZvi2c9NGMNU0pYjw9+AfIE
coo+NPNbXLEVulJAh50zziJ2MTXv5eMexZR0zvcb2E7OA8H811eo/kiOO/rm2Mt3
q3kAPqmIrgT/ISIwSejOVRNEQhbqPwj1gE1hDm5WlGUtUmO989sHNOsVzu2RqP2e
lXat9tjgmJez4jp7KOYLcqT6jRl6G5R8P5DvSvLqVlRgPSk69COTXONZ+68J5ttQ
JvpJh1083pneni4monqlP6VN7JIRqGqCw+5KvcbndaWplMcm6vgFONm4J5igRdvp
H0iY2X80El9FDioCpx15AkbqiR7PP56blgFfGKI7EtFiqcqQmjp+h7ZXNfBxdHFx
9RePmflIlJT1/xmB1BPhGuDehgTTC4Ha/g4IS1vXrFrApi5Yr6iM3YMuW2GPXkna
YepHBbV+zo8YefOuavFKdypvsXhu2SMtiS9PAjeWq9oAVvmpTawuFi8+LNgf4OuC
veB93Fv4F3Y3YKic6ZL42o0v+erkg+aZgO441dgN5MQFoh1aREvREprHHEqXsio5
ceukPvO1KkgHTN6pK8zL2jbKtt1L5CA/9jPwqpdX3MmTtqcYg2tgH2RJG8s2mAGl
dFMSX1BcIDmK62NKfaX03ET/U1+HvbGDUvdcc0DQXQScm9a7+kJPo63wkjYAgg9U
+jdXtlwwclOXMrkPsxjWNfpHHKjWqNs03o686Mcd1IPT85kGPoeEIRRymcQ2UkLK
YoYS0NGwW0Lz9aDNbqBKKnQ8EfIgR4Z5MYVY6swKyYbBOR9K53vGIOha1CPCmaln
7LRR+S5aB0WfTPOZNLWkRaXDl3iljYEN2D9co/w2RcxkwcGkU4Ax/iGqFEkewQ6w
AP16HibEihDoLhN2HvINkScXRycs0xn1TJt1H2Dqmy5YUw/gINc5Eaqzooc1sW5O
2NiuQTnT7pzsag3oOudjMvaQbvEm0xuHI4Z7ZLtVTEWzXkm80hPic/SSZwg3gBrg
Zki8ffAfecKlGEuV0GSbH7KDbYxNlY7yxvqWxuu2GBpDHjKxr6aAvQPQjrFPh7Nf
fQRoP8LOdYN7CSAIAP66z6vLPr0XhwdBGnW8fFDXz3kSRj1/15hIZ2wHb0ENqZ2s
yHpXPRHQRcA3rJbgoSo44fmdb22tiGBHg8rQTIg/g6N9XwMsvKLBQ0709g0cv5WJ
yI/iSYF1p3b6DsqhUwy72K+iU9qmUS3VsR/2YfouxyHevlFNIzu81fYaaQiZ7ArT
FOISgIvzMNKYYTPq5CitP2U+Jhen4kXLq+hQ1RN9/V/dfyOMraYFnNfzBydiwn9M
9y2OdJ4LmOFcsa4VMIcPycE+LpFuPJWCwFqy2MZzQ/chNqMn1i86Noz99MckVxK5
PJ7ugRSPe8KR9bRSCqAuRI6mrrnjNy8J4oABEkrkzpSgLsZNduV/VbD8uEhIS/J8
h+So0uRWIZN0OareJWyLqKj/P5e/KFDiyfM9fIRy1x2YsxXAk+N/gvpHITbyBp5k
XAno8jpaK+0oqA8pS+7B9h6o9s5nk4lPUVx5cALccF+9ZJxDkOgjSl+MpBjw0bIm
zFf/itlI6m4hzayNuh6mneGiXTJR4+vw+4eAXHQTnpsiV8c1DYT17Z2TFRJkHdaN
g5mawlrSwWFYuGduU/Gz2eEeM2Fj2Q9D/ulSkUT/bFpENQ7fTByc9T/uS+LZIF5l
AQrUQsxpLvqcCqvR2IHr4SIW7QO+KfZbVxBvN4j9x8zuDc8mNFmutpMTveU2xtVR
nLvD2N8m6ZGGbfHJExw+iTLXihD+BfoAgwLeLpb2xW5aP9duBpzWJkS9DhZMUffD
ISxS6lw1JaYXzF16V8E2OyiHJVGpOgvfGpTv+sJjehw8PiXMtbRmx3bHtvhJCsoD
4mpW/91WkAHvBstNFu6knnXgwZpPQKX5JKOWsOzqOlHXNAGIUl17gcK9Ng1DFjk2
6Bgf19Ggut40xDVn2fR674gpLh8FnFhY4Hk2umgnkasdSUtm8l9BWUdd0XhUfklP
zAupZYyvf5DGVH8abBaKLLvb5rfgG4xGZnl0J4n3Q9Xbger3Uhc2kQz5WTdIuy2d
LpgOSFyUX104Rv2k46kQzZxufQFM0zo9+hT9+yvI4rzIbKQjarxpGaV2ufBS0kux
t6W+BP/pezb5JTG1TDNwLU+8c5qapiYEw/d7pS77BrkFpowv+CLdUVlBOITdmBqS
QJHrFHqAzAuMzBZ3OQTmmCSgutRYMqVQ1gVfIS2epPEPgEAf1ElycafLWlFchfh3
F5WwXGwQ7bC+PA3BJIVklLN7N3etImv549TQo1TcOL1N+M317rX2N9NU+OaL7W8b
yvf30GFOiJVHleSF8M4F85VaSU/cd6+kY16Vug8ALB5oZwNTUod1AlgUXiIhi/RU
HPL5/QoJVRuREkUHlQIb5GVSAT5kHWMMJlQKHM6eHxLVF7ADsdsP5TpcWvaB9wSn
BPqXcnIP01swy7IZg03lGmQ6nndVPOUCfrLezg7eJp2VAQkTjAmbVERR0AY1Zbi5
F6ej2u9M0uhphttrHQ3nRRtqYpjhek2b4rVyBTZ6/VEthZL79FKiLV4U5hcKbGpo
mxqIpt8W3X2vKSR6NUmTbz7mYs8bLyol5tBsojD+0gdX93AygaewZyMopQOCsym1
K2spkj6Mev+ZK1iTTYMtPiqFtsrc/SJgGDGrvcbNEbp7li64wtixLNpxvN+OyYrH
upOxE+uEt2v9E+QBe5bnALB4iXlg6xxsY8Mqnn1D4tHh8QNRafMl8iQjndArOq/R
gxftgdwuj15wuBU/p7EWYgpsnGJ4Brj6p0a50BMZUhF7hVKQitAcI9frgwvOfePR
nz9bnpzkMC9nWqMPUOsx42S2Vp5FSVWZCOA40M0J4FhWhW0Ix7Bb7cr6mUzWK/S2
FTPQHupnLd6iswCh5HjF5puuhWFq0HrGMTm4DEEYnueSP5KBMIGqGB6w0kG3JYEr
uv6wZPgetos6WmZUX60S0uXpyWMY96dTLx+eK9QqlBSWSpBQN4HYHueJrFG9htIk
mvLCWGNJqoMHG96jGHNtJVp0VWNoVo28EK4APFCzVlKV/d5O7HtHvAUEwc+YsJD5
KbVRE1qd4hb7s69tO28OcnvkIr1KDFnrvfyrWLe5mqroeLgQ9tb8/eu0jQOATPJz
hGpbz/hulCr+H3SdjXkEpG2XzrbJWo/l6HddVf6ys05rXIVegHCqaGyBu9NZL7Or
w0E4C5d4K36bLl/L3EHTs/+EfO41LzJYOYPSC2e7DZmKrrwQb9jH3LjaI4kBeMBh
IvaFXAqeOPaSCtpflh5N1SLWJpZV1lE7BIzSGR0nNRStE5IbyXPvMUZVBVICiUFS
bxPIJVykxMu3BrYFHc0lqQPY0ZoUw7ivUD4jJ3fPn7XUddtFYO4BvD1ThAozfCZK
HynRcSdzvd4Q2CPx/0uqvMVzlhrABxBZusrIZaV18VNxP2AOBCQkp/axAsyGKAgo
FbvgdSJY4o4NzsJ21jRxt93nR4xN4g8wP3xv/Y9afbL5AiHP4f6+4XuzFlfBQ8xT
oG6NevEPlPdumgZo2toY+vcHV2AzAyCYCpHZMRKcQVTeu2sZXXBp7UwrKGJIUPp3
hUtfwty8lxu3eIHcdcc4vNKh8ofI7AAezLlirLsdVXS54Uf8BAV8N1sqT3KNqpy+
9IzZXNSn6eWBljXn9enZ5ewMNNkITAy/LQ7fpa+cwSEbw5Pvs2wuUzzwA6fkOjPs
F2R47WP/yc9VwlyTLqjMRseKlnOO2eXOF0i4pZiYdM96G2sSxpJ/abLnymVzPFj2
hEYSDi6xmwvpr4wzAp5WXa+dP9YM4moxZJweWgX6cWJe+0PZrAkR73U1rIbzZUFu
geroO2GcNF35bcuuUqBfEmZzMKsVV+leSblFFkY4k+q4Gr587o8sjEDi46ydWQX2
D1CsXVycJ7LmsyaNCDC+zSEQjEt0yp5BaijOKrrxgObDExEr3rQwJjt7FGdnJX2H
1GZUQgT2456k1Ui1B3w6tPpkr/QenFny8v9dlhfCN1RFrenuayECU21BxDVU5hWs
2JG8pvIf0VIODUVoqLWKLXjr9PrXL0vCjDzT/WRy+Pml9HHd2lLEhwTJG/VV5rEW
a6P6BCcTpVy5PKlecL4pgjFqP/myoUEIXELJPIQ55LXG88rNRcOu3+XxAT57KpJC
M+6rjJ7n49tSdK9dhwacMZ1ppEjTarHcgZ/0RtRFvGvOiQnkhN/vPvOea8XPElsd
o09uJmrr4FIuEiwZckUoaEIHOH5s/Zy4//AqEQdeK1S19CH73H3Slb+kGBgnMwBH
78gqRs0SwxEwrFF24S7xmP8vjSxpCS9997YB4q/L5Qb1UF/x80OQljAcpQjaujbL
6UyNbS757oB+Msmo9pLAhCVWddci9HKwbM4AjtAkGq1hIZt3X8qaes/GQHM/WBW0
Yl5qBnfCkiYZX6kuw2ccyIe786KXtstl9Xbuqtae+FdE7NfVHViFdxmaIkMWsYnW
hDdtxAQrKdafVFeOsJF50W3vD6ILpnTITxl5pKnE40QF8WXjyqOwGEwIOLIF8lHR
8XQnJnKxGyIlmBM24SDozCnUkKpYO4YolEcQUgwXikPsVrb26Lr6bN7xT42MK+Ot
z6cr10Z1cs3piHCLs7T+W0wBMo8skCoo/i64V0zW2EzKUeYi8RlpeBpfp8ietc6M
rypaoZxDoKkglEgvuhT1tKqOxQTkV30SKVKIxC44eSE5yhjcfTLVilbn3MjtpNTR
ETq5zpTIryVZ7llATzAxDWyzrGKN9uI1+IHX/qruf/3VOvnSSOgkV9obYfoF8xdk
xKaAlNCbzMf4ML/3xzdJDCpmB+gj6nMcRAm9fPSTNIEW7ExFPppKXY1cetGGKdBI
lePjAxKBwBGdZshH934ANrDxKg68W0PBl2tOURgTT1Eph6x+z8xzs0E5z4U9h+z0
1UjwQB2JGISq4TEh+vxboO+ICwrckeJOY+Yfjs6xm4jpBuPdHq1YtTf6LygzSaSw
u47M6ITgLg+sjqEdw8aCYtJgCdzZYZ5e5PX8WUeqkVOLcIhc4pA0tg7bimVvbWJf
e6q6vi8MSD5UlJpi+hyfPnG/lY5kWHLHI0LEaS1N9MN96QmoNUw3XK90HIAS8WmY
Q8p7bbyd+gSJhm2VjmnOw4vMJby9kmlzGP0FYkMVBjKlfYvaWqyPH/Gaqpaop70y
lvdCxWnfiD6eIEbZcyAA/aSdrMJcd/OrPfyLt4Vn6GvLXfCz910O2XCmZiqB8S5H
mxUvyjharN0DK+/AxRD9oIEZ0FQrEsyxaFJg73IRnyW/PaIO9pF0mjicfjNr1eu2
2CDGluwHOzuXQxHfRWccKjB5byZZy6pF5eJN3uD4XTS50uhAsHfecaVQ2exhegLI
Hjumkkzm6vZpG0A7KXlkPvKddpvVB3sV2Gv7+lxoRJi3y7p7r4b6K4RkcykrTdbW
V77MgiDTgZTdMlqH9K2yalW25NkHI3gNiPEGnr2E/9KxZyVvaKkDPSqhARkrld56
6/POfdwxJa0/NJJgKJOlk4oGWeu6gKxWsZgBwCz0dbeeVUTdgTjGvx3ZnBcIsrdL
d+QYQGsy+6DISSBmhxHZj2nVIh2YupMln7Huq8yTPN/JjWMDwSYUgu341EOmq3tS
WZ/HKAVHeqOgpgYJcOVovh+7fBHGvlRkRgk9eHGDsLldtpU0OigfvfCL79EX99GP
R3ueRNcLQmLKk4myoQ/a8WUG375FXsBXgIdZs4+7OoW4yiOEqer1g4ljY80/3TUD
IGhHqYdd4Vz30Vv5gwNfCHBcKqKnIqBgzty4LqZxenCigj6fpmv53GWGo3igKK7I
MSyhsNJ/5wW7210zOYjvn0ScUhs7Fk+t1vpOPgWu0R618BD8HPlXJMhj/obs/rsc
3UTvcoZfPZBAGEyoA5j+1J8+QXITjh26rftNXezyfahZB8mqb36Lm+cDJwKgII3x
LbRfwdVHBpHrm7uOgpsYl/CgM73zI0TlyefyOUuBLPzkRQ/xR+QgZ0N4SM4VNlPq
ibPgpV6w2Tw1p24qYaY4o2LgFz1WLUusHJh0t40lCS2RgnIDzkIdDJCZs+WSICBk
Pa4ZKXF6SAt9fOchjXAERlK7bcycvHKGknd29/8wuQ2DR1Qw+AaB8A8H60HQDhgA
CeL0YLbKQSu95tVDooq9BZXmOxEay8zm4u/RtqD76Q95QwjKMIPt1LrquX2Wwey7
vqI8UiHGn3CKfkENUzgKpTs/M2kTvmgDnNbeJMlvpr1TCeK9LP0gUrmvlSfTzo1z
quVBI/EpzESuo22nH54QAaNIU0nFirC6bDu1Lfc/XuuuEos77FOhD62x5XjvndrT
BEwinBcshUluPLfvbD2Y/SdeXklQUf0hIM15ZtOpsOowakPcMSY8/ne3j5ZZUCQW
VIBP/MDVYetfB3zYwgXOGID6or+2aq5X9pI9npDAqRYsBI2IJSucJ+uDw4uP7mo8
F75wG7R5z0OFo4D91VNhaSNrlG4j+P/7hHaphwFVFWSUTMiGqhKOojiatp9r+OA6
wwWbvDp4MvccLbhnSzIvk1KocLftaotSjxFTFgC4INxk5nWo6WDy6Pj+QmFRwEWe
GSerUk92SGmM2k4ZBRHt8oX8O9Po/5aB1JgrvgxxVns9kUNVxNtUD6sgH1W9zFwF
CWGh9MmEOapI4abmABs/ga7EI9CPFyfMtFkbO4lbQwGkkFpEekktvtiBej+OYZXA
q/Aiv1+zztV1CZMg33R58LugFkk06iFNbUNHHVK0SierAS88MkID+ulFUplB8Nj4
63b8AGq6QomV+zQR6XB3NlG9LvLvsca8sAaSqd971shtwzyuWq0nNJPQpS7JgND6
Z3Gu/iOx2NJg41XiwsJsiBt+BkCJZjEL6NMdGrBWPxYKE1/LUC+Ky8RfVrGIMzYx
uxbGMJLl+uVP0T7HQq4vpXgQ9zoXfxMyDTYQN9ErPRj77KiAOgQEF5Kf67/eO92F
nP4dgYhUn9JzG7tk/O/D6slsuv3pX0usEPYHBFMjJrld4co2C3fIGHR1TxV5QMxS
H3YuXMzE0bD5fjBjLPImS9goyuDYAN1O6JCnFSc5pdMar5YtTURiCUAw7xj21T+P
FTq9R0udAEmvowQyyzYffSJw9WXb+Sxkn36rpDJpy9n+CK06Fye9TrfOtueXsASL
TartfLfqDSfxxnKSdL0EsHp1JDvkkagIrdXWoEH/tveKzm+rYrJ+1Gb3zszGpb8z
0WT5zB/IPCrOA2uxS++j8hCg6WyorXnAueShft/4b2RjMI5GaId7POXdUPvmWtN6
0i2ztAeZQiHjROQt6wRskZtlZs7C4GugVb+iGjxVnhrzZKQbsahtrbRwgmCIgnSZ
u7GZfQjqaa5oxuZBH67aV3rrNvdr1L6bTLPzF8WjcNK8ojffw49SzWeqL9Z6fKHG
ApLjULlg+xO7lWkkyCZn/X6beoQFhP6JeVxhCAlfd6nx4KdlvLz9GZVk628P0Q+C
zZ6h9YxR+SQuSTGNNqNJ2g5ryzM8q4bApKqod4y4lQYQ/KAoTcBrpc1heJLeXzVP
k5O9bMIh8G6eAEhC1FsrPy35nqJ9D27TjqL2zxTwc3G/e/C5CLSF06pBMP/glCcX
6d+j0TVwllQPXChmdljHkVKLYFlTrBddzT7/dPHHpm+aoJN8wsSIhmcQ1iQh1U2e
QcMNjt9Kl79YlodpAqshYDfe9L4+HuNK9D/D5/cKPjxAW3Jl/INeQTLa/5zr24ry
BWsz1CjS7+OWXPhrfENDFpNygQIMMeJf1+4gIRSMYVaMoKoO0vqTMQbxStIRixhW
7Ds5oTG7Ivwgh1s0N2d1Oaq03Yk64EvpGJqvIm2LIuue1Wmb0C37uGznvAI/7Uui
dq1pgMVVjwmCRmGDOpyfwPYxCmjighGnodMosCapGytIM8oAAzhrmHl6c4WtP647
bq+tSGLeZ8agLM3enhj2qBe6Myp8ngapPDXhqLWkkMBMun26Igf7U/AxFCa/nKj8
Nh81uQ13ABz9mlkyVAdnW45pFvq8iW897MWhtqsZ3neGPLSrlP0cbowV7wX9NpdR
FxUdxiQQ80ACO2WJTqo0V3BKNmrvevnvPXab8zmHXIlJUgP2So7gdEzynDKfkC+Z
8i4fJr9rmgNcE6ij39bMyc4Vz9UBnpmRQ76/JG7KZaCuZUPhSL0YqOLfjQEE8j6G
Xp6JNqqlOyKawjuvihwzKm59l5l4oH7v8VVSM5zHiOVizyhM5q+nEIEijEWKn+f7
woRoOXndxdYaCtBS7Eq68HRREGft58wQfl1ejPI5pTEp/GHgc36ZkX5N/Liv6WlA
xeeLal9o4XIxEL0J2ntn+gcTKcIogMUqLfJ6C5CebKjQUhhM21GhVHNIEncnMpDj
BnmBRZMnL34dhsmRgZR5jmIkBGeJ9ogxXlYWueND0acYCRuFY5CdM5Msn79dSN2q
qBKxBLkbIBNOuWOvo0vPIjYlRu2ZM/MGEnjnhTWlmRontjgih6aq1GGUz/Y9pOO1
Cv0cXtFRCPcT2kWW41nEYXoI7erjp93TkMr4irEuNNkswPbj+SOY2+nYYEAA033h
Bxzpi6c/MmVdNKtmRM9Bz4BBUqu8yHMl0le6Ezszd+kDfMY98WddtWETeOXbF2Zu
dxrJp4PCKvhQnTNSH4BoyHEzG/RGpk1A/i/awI79w/qz60Wy1lk3oi1oZ02M9Pj/
Ym59Dj3y0Y9qI8RGeRX+fPzPg3peNxUlnPgWIrjXuY2B3IlBtptG+InHNsDlWcYs
hYMBVjuFw3+phd3NaKOVVLUYwBSBgeWAeintLfbaRO+BAeAOXsuucs2QQsXerXMu
ZifVGL5VM7RSRKuDHC+K0iD+JdnajczS/vd8/SR2m8SdD8Sx4Sifzi0iLTGmUBsy
7FdqS3xxAtUrGtrTCSwANY9CeqR/KPJI/KHFJ/q3LKq3Bb2AtPhFrZrfbCPURwrq
drS3esm7UBvXC8J6opB0gW3xehBb2es+aonhpoa9T8xUMZNPvAsZEPaea46yzn+P
pLLycr0TiesWkk+1pd18dSnNytIllEas4j9klHBztG5SbUCnDl/ThHNAOqq+DSwS
3fNabTeUkgf+DvkQ8pimAurwbtHEJDynd21AhuT3WarNkg0H4hUWRk2Kiaxc2iMq
bGk6aMar5XwIOKNH03/XpvgLQp6Cea0i0UxeMBYKmqrs91Alz9KhQm4EQ0Hk+GUI
GuRDkg/Ousw4A3iGjwWsuEflnOf33srcGSXRfN9AZLI4Um2qy4qpIFLG+dpjh/Ir
L6sj57Szx3fID0nN/FhUDJo9Ipa8ONb49WJ8L43b1iB8YQ5BnpegA+B7rncy/NSZ
/2At5FXfXe34w3u0ugNwReddZPpn8+N/AZapyRH9szimB/+ZiYR5xycjpqi+AAf/
Z6iZqdfoU9AAgK+kWeAQ0RuwuqZKcQDm7Q82VIyN1qSyrR0CwW9QNFCuxXJPWeIG
j3ZMNtWynuUonSCxubvqe1k6wxstQkwfjJth3R96EioSfqXIbHGh1PcmmiVFA1RC
yYx7cygWx2yWOOGOGJQuCzJw1YW47fPmR0AMcaRO+KHsvSCRqjQip5AUaCzsflMC
P+tIfEbVV+un4xE/ohCBmMMxsWqftR3h9peUD1JS6pyhZQqgABcYOzGSVYMdQB/1
dStBMQz0R7+dZG9agkgBmvHj0+tbcAz+eMBbKssC/KLTqmJyEtAApLiV4YGDKYuX
hPw8WYC0BHIUok4rMju3ylVnYc1QvCGYdCf5853FyxY29JoCCvd93xzZwiSN9XRe
gIpYlKFywzUb6yV1OS79ZlgJamklprT5eLP+NhcNmd8NI0sJpigvnTsiY2DOJtSe
Svtsp627EX41Rm1HOQ6jrRBVInE/ow50pWCN8faho+Ek1CO66JkDRnvUGK0uNtfV
j7b26OqFeGbEMEkraNFNK17nQgpGkxH7irBwTlt0IDkXbXvZWtrH0S6tgqCfnYjp
2rL8v2QeKDwzmHLQvAU4xjiC+Oo6837yy1Sgo7D0IOULaM9qWIOjp3vt90Wds4qT
4LxLuauXQIigWhiLgB6GGfDZJ8zFWo8xKIvk2wZTKmkJRSRSnZ1ODfCiSNxYmSvW
8AlpSJRYLw8fWDmfRdGESCksS6nibiQP1+4QSNkQOq8m6DAtLnMOXFim1nN36uO8
U7VTVsZDpu4ZGUbkkmC8BDm0o/3bO8RdxJTdVsVo3u5nXWRjvhcr8It52IvdcWW+
3hOHkGnt+KjOnRDpTlNVHXHTefQgfY49FZKAVsFDDz1XYT7u60kL1Wh6yB+veD2R
hkMVt9jM/UM1tbHew97PSLqetUgFiU4PydhIgNot8EDIcEBXbkuTWE3Zt4UXy+4S
OOh/BZbBYaKH9MCxSyBKHd+gIftoV6c/xNJHmgZVtNVJ0KkQnLUkNBWbEfHvlxj1
O+vIHkLi3uvEO3LNYgJcpZugYPYjYqdO1d3M02qaApELmPomEYUoR/DSotyzsceY
PcF64LohGoKvzESliMbxpkYU94TAUs7EugUo/ISbG54OX4HFgo/NQ1S7YC0miEtr
yKnUXQJSjKE7PA4bQJOSgXvRbkrJYvdvphknBBaVGVPXdDFmSdKx9gETrjvk7nci
/fsdLfNe4LhzcoGeyj0oazeHxF1VS6TNR1bypuhNPQJayjF45xRVQwF2/KqgUL8g
m1XTCgKebXolTqQJbifFq3ZXNqMPkucy1RNrgVFvkfW4bBkwc/Xa+hcQ5duI+zu7
pojFQC5qQQlEOyFftES2m+q/kUgSKwjpPLiqDlWrPaUyO99fBRgnelQtRKRzFDZp
T7I4vKgbOvYwebY0XPCZvpgTcV6Emu++8L+K3wTJv0a3ty+uyzcAUQmHRMuxcwam
AcvI138WM6IJhBYaZmvKp0NIaXF0FL1EMyvBHOpIPLwL4etm+6hNcJyWTgToysCR
AiBPqgffzbA5TJc6kBWRFb/aybrbW60ihNPnPzEfbJytnLTGTNsoCzJo3tN9EA90
qgjzKSpb9Qy4tBmxyYMAHCJ5pg0HGTUaIlhzqyFsSY9MslJVfFz7yGR2C7Lzb5hS
`protect end_protected