`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 3520 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/9huKRhRMtvnNqb3Z+UU7TahEoHV+T8U3P3ufru7l1O
3DlgtZzb9QxCbOjthp9+wDkjygH0eUfDrEl1ovhZG63CAp6lUyb4ybxFL191PVWZ
rQPQUv8HQFZhYwkhjqrXZQIZqRBa1Od8az6Ij32LqSqyJDZP3HUWfqhFHKG+umDN
7wB5AUY3oh8VfqXoOP0H5HTIgJ6R+nJb+LewB6lCcxdGUZS+KQ3ryhBLORzgOkHM
YIk2dX5xlzinxYBmiHhVaoAOaT4J6LYa/FXeBwGEYESL5/gro92ZvfL4+RjTEl25
rRbHItZV36dHLo6xpuoA9W8hUBeoNvQ97dWcvtiyQ2+FUhqL1ZlhdK22UShCcZct
ONpF/Xt4w6pVx5hMvbRMt7iIFyYVKvDEZcGnuIi7q+y645ymX3UnucwQNZa4IKlM
1yNvF9nii4uVuFP4DwgNua+n0aiBlYwNrxNrU+zkpD69zAprGMzh7VEoa2/cC1+d
gGk+1SXgBySwrt7WyB8KoHdA/WO2EU32W5bsEPs0j0sVVPLOi2yHESqlQS7Q4y+f
aBlsm9/ibP3MnggPoK5mR+R+Sd0Yj3BIn4FVNMo46gL0b0xPwfAcEXwb97a7jrc6
oxaIBxudDIiDk2JrhGjLYRVenb2S5PaxBMY7ekajLVTXEzPIoxLFvqSHSQa3YXXV
XP0O9kAk5bJRqfmCYr/v5VTYQetatA0G6F8o5fmPuIepRa7MTVnjxVk5SmC6Lg88
scuJzFBNerrpuxNZQrzgLSfZfCuMxnA7Xwz0n+URGunZbgk+12MPzbAonece4rad
n92cQgqxnND8x/h1gBs4C0ea2d/qNlrz9DhKcUUi9TQICRoJhkqAXdVNvpUqxePD
WReR2sRO1ojQYBlXCZHSJRbi5QNkdO2r0xEGiXBYYHmuPoTH9oAOeHjvGk2EVtUx
LT6L7Wenk5KU84ob5+GrZT2V9HAba3zHzvp62bOZohGDDzrKQtct/uoRv8MhCws0
cuZA2R2jc/+SdntfYc5AtTZJA9sTTfPh5yONzD0dOPmY0bPC3Hci7jOZaD2/EK8k
4a1nFfoNgexTtJUYiWA8w3bZgmI0Mz2Ucdke24T1QlwhCLLi30CTmGs/aG2t09wq
XDQ20mg4hcOj6L9LQsI5jSvZnXQqJX+a4h6aYkLkO1E68Fm5cA2imb8xe9t311G4
UFVPBrq8FQ3gDeRt/DfBIrGPP0pTgFWudP8xqYFg+/Hm60BhZSn1ejPcXPdPA0bL
H1A7uHNOJQ/PdNj4yYQl3cErExN/Yo47UCDF2wX3LFTjXcz+951wNSP5UHKMNDUz
lhDtGXczyxuSqi/5QkSxcx7rcptsEFgsZk+mQbGZpT7K+EcOWVsBeKeNL8+9HJ90
E18iE4zb3qMQYM/lskENAJrQgVwylG/gdvZmEl32ryYUR/CKFZt+Q9M+M3Fj6Ya7
uMwSzkosgUbm7NNAWJy4b7vf+UahwWy5DL91NW8sV5jGYC6YZX66wiOTI6yAuKsG
I5bJLyiy5oWdOJTON7RIf8LMt2WkFcGwrq3QdN0Y42nV695kDIyHFNuItSgl0Fga
J5efZYnNFcIIjAU+8kOen3eDR9oIQ8ZBRl1J80Nr8EO6dz3scZW4+l+5iEFIPCGx
kzJsD6kYH7ZO6HLAf1ZcZlJd1dMS8icbwhIOtMAYcKuRyVNbb3TC3rXko6Nme+XH
92Srh7t0fFgdCBcqiD8Z609wrJMgG4IxcD2Q4bDQPtVaVJuBho+VSB5j7Fosz3Uu
FdBA1iL/Etcu9OqY4MVTpAJbgpAA3sHL/6CT/jHW/3gEhYzXWm+y6sOUV/GMyebe
Z+53noD2IFDsSM851hmkhee8jt442kWBvKsRoVesUjKbNlkFRLdt/tYYiLclfRbC
+h1tCBY/IuDVbAxep36WRnkiT92P9fk+yVQuKK282z2rS9baSBF+5LnUI6JbJe5J
l+SJot5/73vpFi+aPTfbY3km+EVZBuEdkL0Kw/2kC9GAS4pN2jqzWzUhBd15OLOD
XuRlMY/MhFEP8TUqkfXXwtZEWp25ySV1yQxKXEFhJikuSdHPG8jvmt9QRP6zteGw
2XCYBC++JtNsXtfSgjcCXdxesfDV9u3qfadzskFtJCJLMrf3ph4RyXDxLRgi67kT
pForYX0RLOvd+zneOSeENHVj4Bjace1KwfFBTXVYc9YSGniYA5O4IBgt4JlpxMEt
CEyl7cHCoyvhG+ePA/a9eJlBtGvHS5VOSUJ2JaOiK64GqVW9ywbpRbQC7BCu3nca
2AVnkpY2zS/fIZl8wVMxA9GKFVxUjCmMBpcf4g0zF17LcfcXxUNQ8rQd3bDKE2Dg
SQzw2bHgLeXmL8bDCKnBRzrtauGoPqZfqvYXZvGJ6Uj3KdzgnOo+aJ2psmuyMslQ
8UL3TCSBV+Eiwwz4KUUu7AdYH56pRMG77pKdeaZQ30Xav17G3xOsEkpG62BSIvqZ
fePQ102gBhFbO7l38jhsy4MxOFIC0gq/vPpFMuYWlQk5xlCN8GAP1jW/vqlW0Dub
K88KgWtSifNv2EKWO+7PWFgHuQU8m9myy1IS2rSvNmA1NPOJCj2Ycj/fyKRP3KJp
+ZwuEh8RT0Ti2+a5WgF0n3+o2vn+Be2OVKFry4NwNVgNJFZ3wQC5WXY374dKpd1m
k7a+sZxKRiWGZCXe2jCdezOb0hukyBnhypWOUMl6r83BeNHGxHoNyVhzdkdc6bk3
oVSRfl+pamClpqgVmhA8ErmAgpQqz5n3Nd2//dy/7nhbEXFBOWr/u8cgIGDq8YQi
5Zreb8i/brTi5fRP0FR4lZUvx/4rhuy479SN7su6mnf19un7InnXZT5QLhZxfTGL
6zUDMuPcPSFCzJmnMf7NvG0C3C9QOY9/GLt1hk+CPmx86PDjqLWU/8C9uOr3dSgb
FTua1OAz3wO3T1d8um+6K/jnryTnYFogGMj6GVbcGMsnMijHFb9q5U1xIMWzQKc1
KO25C9QE0J7W68T+MJzagKpq8Bpo8Ap/Qbzc71GDA5VID37t5qJYKNcsYTpolKok
C3yUoPVHeqMPps+IEaZ0Io7vUlFeN1rohW1+kviBFG9/Gvp7WWPbleIRg4UiGuho
wWGaS9x9x1SYJSFT4iGo3z5RaW/aI7SeXWdasukR2lz7tIv1mGkN9vTKoShxbcuE
1EY/oE/t28j04JDg3wn9PAP9SLhS8vINdD1+ZJ1cXZZ0u0pm5/Wd4hmfSP/ZoP0H
Ppj+cElh12SuTXzElptApscdFEtAPZyIe8FBZzsT5fxDxWzgU7VvC3Vh1zMj9CX3
6jIsY5GdTY9k0qQhKViig7p85hFf/jRUthbMb2cMG5ucUyuXswAZm/5PGU6Jr39a
BKsxCdDnG72ik1d7aYpnGaaAcyNM+tBnLmAqKD/B/GkvnfDSjbTALqWu5WPRhQhh
AZpOs8TaXyGepmMHNwULw3W0EMaBqmRqAGmnXnSjpBSFR5ycw68srjY8djJj9OO/
L2jKRyXe3DXrMDHZVlKf+sGkv1l3Cku1MD5U+tILgQ4ZeXKlHwJka1A0naOY/oqr
G2yzr/v9jB0kHZS7rPhGnmr+0KaRekjllHlZdB+5uP/4/ZOiByRjeXDLEhqpxwAE
/dKDBq5ZXIoEcFqwYJTRifSnZnZrZ5UboRbXYaP6tnDnz5s/1CZNkvpsndVlSxOU
z8ySQKihwoi58DHSVYRfqtJS/3R1O5HKy5V3jUvKWCAZ3cZ4k8R8QYTGL9xmKHdA
U39Voz5rP3pat/wzjSuSMU9akWot9V9WBq8IEMBQZn88wAM+OmG+R30RQonoCe0F
GZ5UEN/LE2o8IY7JOK3IhGSu2yTEA1imS0etV7Ea+h3aQ5GOBiG39+2Bbxq1+tka
N1wHa1di0v3Sbzu3rg6EOvMcdf3MBrKJJ2TFqwayGQgwId3KOyOlcL1mutwXu3lD
V8ZMp4rGLQ9SwDMJHUQsas7Fi6QVn+8pFvDcsVwdaQKAH+bvR5bMmyGY3hvpb1tj
gQhoxW7OTvSoTf9jiRC/lNW9MRzOrYgDOVtUT5ie3ukQ8jbscWS+xkMJjvjPxDjy
vimKMzsfNIFMCOSjS2l7sgYHnLmqlwOJQR5D9N/vDI1swALxmDGz51j6mbI0/uf3
oLV5dkZdP3CPkiGhyo2bVKpWDTXLynBTKVUZE+6jztrcUXbXlMll4CQDn6Gs0XwK
NUEAEL3LE/I7Bd5fbkEXOpHRvR5jfx7mqfN3NbMzOg6iXMV1QlL/iTcdNCXXM1m9
yjHuqOmqNVorG793zcqP28AFqKZbya8Lgscfbk8FcvcIrogEHMQ5ygt4GaktuR9X
+nfhrfnthjm+fpRkff9rcfPdudAQUq5rVc/xlJ0CbJHyvzG/CWeiDW7DtczdpP2H
O6gPpWAibzoGk7J52FbfTW3UXYh3f1u5MAlbqkTCvVhX176F4VA7ljJC2cb01LZI
MhWexLWxLAG1dHt4Mgbwvrsy9/099Nq4XWQP+jAMoV4FxaqU0eaWv0SC5h+Kqp+9
iHhWEw2NkiDrMi/jljR3fb/EUJAttJq27VgEhY+Wdwfl0stFYfhlT765/Nm60QDr
bg3uHGPL5JD90pTkmEt2vAQbUDNefpoO4/m3808rpC1A9WKqZuoJygGUwUNnj4No
PF9kcrMWvDlJE8VSEzmPzg==
`protect end_protected