`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 15248 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/9huKRhRMtvnNqb3Z+UU7TahEoHV+T8U3P3ufru7l1O
3DlgtZzb9QxCbOjthp9+wDkjygH0eUfDrEl1ovhZG60VqWQIAa5BuV1zqfIXAehW
Vsg8g+4iW/t1S4HyvzwSBHlm61TDO0cA/zPvXb9OqNkDamIAvnfwLGdHHlNCZWLd
xea5hVvXvUC+LS3EA6hrkukxawfpUpmPaoEHqZpa1ePLCRhD9RvfTNyraBqmeB7U
dshNLSD0cEICjTiU7uckSwCxFkldljkcVuWqLNX8+7DgyhxeHeAzIzQpwpoH33kY
F1SIiMxTCKskL5a1pxNT0rIYD/YRIQkbcKfnQo62ukEklKcVOVym2rOyr2oD2nrD
f+tNNISY8p90i8Qcmdq8uo7L/FNnikMhct6ciaHrB/QD7nf6e6DH4WW0yo9AHWEN
FgXpwI7y94VsX5jeLnneFggzlZriruuuieBXcDmsep/ZpobC9x9aD+/jRXWK9wHP
02nDf/M1tXAZx74qcrduZD3p//h6VS3/7jBww199zzCGZxoqbnzlr3jG3SjHBFz3
3iVLJ6LHNtvM1NKVOuV8LRDlXFJH8MRPs366oI6i41CB7DXLwyt4ALPGEgK4AosB
oxiUejRS/caCwRZ9S80aLqZrjVZUrHUn6rksUVAYZHuuz9iaLfZS+wg7q+dj0VCY
8AcXVsAwQ4ZSPCp2jM1+PMQriqExj1ZMJIeP9Cf83EdaRy6HvRhw75W5T/ebCIf5
3kRWSsh1yjmAS1Tex1MnaZxdrfVfI6XeDDo/2idotAQXkEYqJ7qetnWESZ0r3qkW
O5SoJXnc271BzQO5Ujx37W8GgpD/D7KgIXuLQiPFOLwDev60bVws3MV8RakdLjZx
Ur76KhbxKw+/UuTbT5Smd+DTqSla6qfoD9PUocb5NIzpidU9/vGveLVHnFvmDVLq
OHSYPsV4ys33rcdxOWZ+ngVsL+Eer9BeFtGXA9TLLdIJs9w0kY5RXBIQcscyO62W
SA2Qk7Izp1CG3nLpoTMBtN6HfeVK09KWmPZTS9rg5sI2HwHMgBPCG7H12LrJDE2B
QRKpqHS0jxgJqTdyHasXuE38ThVNrmCfcdzNmp6rQSahKDtrPMe+35VlOUg8ITpi
C6mrqTup6yi8TYVuKBl6nZB0KgebqBZF3LQOLsCV9h3pUsd4+84jokFlskl3Ase1
mObStUnJTm6Zo4UqS2/VSvesj8KMba2d28H+xK6wvK9dzXqWOt/xM8gllJKbocNN
HOLHxe77+7zljoQhKkLLyfvl3wv/L+VHM6LFEhMX+WiMj9Q0y4Y/p29a2tLvyt1R
OhF/9LaBP8TxhXLcZuTUo+cMCrhIh60fkIc82qYGJMDgSeGo8RwPn1iouVstImpC
pSC2ud1ujH85w0Bt1BxwyQ3xCVLFo4TNWzJ1ZKJzXwsl05chYrfzVpWdSHmq1Bwy
Ur6xCxRDO9NXQcFn75P0Hy1YAhWV4Tf/THC2owBvoefsKFTGBg2mKv7lQjaViOOQ
Aye5VJAXfqEJJXsL7ptyIO/tbzlPp37Rv76BXD3iapD1Z0CU+CNcZkZeGg6JmBwL
3XV0wj5vCT/ssdrP+xZcRXDvfV4bLde5yIIByiPH6kOnxWj8Z2cTr75Idk5ox6qL
VBbMhTMMIRe4JCbERuG0Ag9rsHe+Yv9C4lDpMg+Y5UjeLKzo2X33ghqVU58QutAZ
GLGNC6J3CEBkL5q0BnA8F2SlaKMi59XfzV7Y1vj+grZTBP2/AOSWXHzo5cUqv/DL
YNkaJVb01zQSbvzhBqho5Ru9NpqZO8W3XCS3vkk4yr5uVhGvraHFXjQkkZRo0QMH
GDW2SltlHgs48juLmQMrIyL2DS29iAJVY8EgugUqyc9zIPVLt5NnetmKSza89wkL
mM1/RHlk6eZsKRQwpmloJPnyG7QlfAUm7YsLhnGQyCwp9L3sUDH0FSGtEnJ1Fg5P
OgpwzGCGB+tIFTsWUl0OUvIXr/HklZvrvsIQD5sJ3p4JXipK8tMSGoIRqh53qIhT
GkCd5H2C72wkxdyoN1c9lb+uMyuNc/+y4Iq0aoeHv6UerUhhepiZEdOBi1xnvOGv
IJx6dbvfZj9vXOfa8FX7tT2Mui5XyNZB1HIJD2XD3ZkOiEJ5BA/Em0pB3HFGLGVM
+Hm37tTYo71sPrpG8njNs79+9tVZUXETH8eCarHVNHaGt2tZqPc5mCUFoS5hZ50o
XqVjl6PIhyIPCcio7U60n1oLo1rMRjtng6TUHcdTva5W5HZh6OMlUvc2p8VeuB47
OcG65cO8sK1je9U/xCW+N99yjZY/jBSjIzWjxTEfa2mMY5TsTHQzuMiVc3Yma3Ef
B74GDIfbxnc5Ob1sJGmV+2x+vGmmf/6oBfJFnkSEa5bc0LuUjHVSZupWpc/Jun/b
bb2OWWp8eIK+d61josg7Jzwa6Io3VGmYNVYh8aNo7WaYKXeaUgw42uOjFmq+aA9+
/qJDXPKr0nphV/Cd16c0tDzKOF4HM/1EXTzA7Z0uKozthpLAUlELFPPinhXRPV1D
PwUUBxkIZW4m3BayUNhjBXV3+wgbp3Ah7NOyaogoqOQFlxEXXB3jDYiHsnSBcvbL
MQQ+e9igHNkX4xJFLs2SfsKonTUWPnw84DAAR6oAxppm2T+zwV5VlGWT6X70y4eo
HNiMCF9mImrhZkZzwmL9RzJ+YxYMlmUuLn9AfvVDRZR9o95RuVghwvFN4E4DkgFI
yS3RnYoOBXpkTpnM6zZy7REHnIV8220Su1IJhwhofGjFouERQfI+9JZuHtcSv9OO
SdjVeQ9xkMhMVp1VnucrSYoAsEN3o3LLRwhki3it3GjNOAnMCYvMFTBorP3Fh8TQ
LfsVxmdTnxL5sy9J7gIpfR53AeSJu4G7wpGP/ia6pxI+TNGEri87ifTvOmdUfWUH
tNCPpHKkOpQTdMjwfZIgesUiNUPpTmJWPGu9XSfP+tAXNOO+YyBOmGJ1cgGIF6yl
2v0+J76+cQPdvfvZ78rvz4GGhGJq633CUQVw3uEzSeO9LhfJxghiCqfxU/GC1DYT
N+6ssewBLWr0vcerLDeX0XqDXKyYefpemUINujvXz/lMplL94lDk4j8dzX/ENmI7
H0jPfijBfC4iOQosw1HTdupBSHXHk4tZJpFL1GMLHpYTA9fQ46Mu689PCwR8NXyy
gn+EsTEHedvsWmc4Ep+qSVWwf/b9nDSQFimnZi3+ZJ1Su1gBpZbp3MK1GUIUpkf5
rALez4xiwpwju0miKOpssDLYf7SnA5KlqkyY3Or5bwCZyN7Q8JihifmIZtHvzLL6
/sz/0NKImuDwZqYzASI8jMe5WFwPmnet62CcoKOb1Ns6jLGzTDg/gRBeGGwr0GLA
+Cb57udMbnwLoTKdM+zZmohB3Q5XrTT6C0PI98fWR/uZ/UqEFBL9+mKfN7eVfAZs
ft3reDkxKAPPWD/K4TODjuBnmsnV+4OHceiEeDOaw/i9pt1gfKYAJA6Xm3A8Nf4z
6YOifPyxIWEa1nMG7ljBz+YePIuhzJZwVHDlcFOd0sMs7JkrzZgqCGHMILMZjm8d
llo07jU3T8n06/itxikLNJw03HTYKCmV5KIIIeLO2JTN38fF00lGoqYSBDbYgdC5
dYwcYV8UK7zXpadXRF8kZ6XDPohdLao+e9XaSdZ3uZcjjewAxpSDvwv2HtPoTFrg
x7MEAwS6eXLC/TlQVFrsAq9ghgRXkYfH6+jACW1XcZxOLrDEIcwYAg2Ub3UXtE9g
ICNyV9krtIdrjLFhMjVBpug/FF70/uqB+eyTwUZzAaBesC72Fw6bQ9wdFcBsQErR
A1DA2F0i79uQofOMSrPyZokNIGr0du2fnsxADEMTY2xybusgxzOHqpgQSeUxb4Om
1hCmomRRGthVb6zPYa3V6uO7dv6EwN7mjz6ZHT4sjvhgR6AcULz7QKRRFZRdMrUU
u1dpnGo/xfgbIfr7jWqOkUBeSlqW1SSSkJ3tbuyakk0rAZiSFk/w4ZDhRrMAPRW8
pGzL1McxXlB8OibvNaQV05jc4ybaUgkBENmZQkWOXKrRpnggM2nfDcR9DZLlPEYo
mVMapncy+Ir9lzsMk8vf/BxnEsvRY0iHux5RMTW6Q3/ebUkZMwV+YRoTqyUJ6tO0
VP357gmFo3tMAJExWbjmY+BifYnUmtuc/xj8zg4ppOX+qIJ5zVKKyvJ9dM5+ZaHv
uwq1W4aQyMMYSbK1zqj0iDne8kRwqEQxyUoms92CY5INX/TSVC0ynB3965tq90Tv
5P7Jzz7icCMziwSNZOLE+NJ+G69L13uNj+64wXDz6DJZDuJ7NUhMpG5rwQNxr8pN
XZ+SRrHgceNWqt/9KGESXPi//pJHvy8mm3DYEbqV/EJw9VDar2O980N1qoIAJyka
Xtjov21xpo+5yZ42KG0CptOPaDyITqQ6X45NlC1yY6AYD6BRtR+ix/hHEdKnjy+T
fQ4w4bcxZILVVbsjZUJnMNQFf3g8NZpVgKslKizL1qga55ATiE/pzOpTHyx/zxCY
3lPr8DxwTz8lgzJp9pYgjQuJnYBpoRqNLc3j7Q8lOn5lbq/dFEq1xs4S31wb0r4C
LN+1G1QUXWOH9sIl4OjIxuBbV5yshGYCGiLiJSyK4qtraja5doECCGXtStxPlejb
iLkPoy6LwmU8/8FGaHEcEFH0sqdqwG4G1i/HUWuwaXO3QxxUYqjy/fxdJP4vAYPU
EufYKO5X+LxPvqFQ0rqUbXVJ0MziTi+WdPZ1N5JLAUTVCReVfuxyqJjTvCsSutyT
rxn/KtVbxthJJ0fJ4UqQh9vo1DUfg6JPjPCBgg9LkkSANSvew1ZXsovze9MV65D6
dCM3zaF8ioSf3hkUKNBB6h9E7l2s0ht+TrdV0lwUu+68qxj41sbbFTsyx6mV+4eZ
blI9PlW9wm0iEImk8su6AOKobA5zEMU9OdxMXhIzEZaLGQ/qsumcNkbMF3LzJo/W
Ps1YYIgjoyhTDwMnd8C1FQacILKwQYNeXHOVEDMMmhQKVs3+nJFB2t7L4ymtzLgL
+/sw3uNA4sCVy46I4oA90E/KRyhx4z5Pta4qG35+cZE7lPYELsFCetDDBjEEMjdm
6PX5hTh7JjLfPjFmxZsxswHiBv/52tavVzvH8tqh1/U4Ky6zfs+FemSFZshaLR0L
iL8kRqN+cfpetRALMe877iSMPaSdjktoSi4gA5rlRpLjGrc+5mWaZp6l+CEjShFq
t9R9i6IWac7qUReHmF2ichmt2QWJGTsEGU/OUL/H4fe1/1uEBvAQ0EfTRhd6uye7
eNIlCJwzDwII0CaokEAOrGD0pqPvzh09jnYG/TrpyglX+H8s1QTZfrOP994EiqLL
oGcsTSaE3v+Lep7FX5cecwSu1f/XiskwpizWVjyGhV2lJE8W2hK+SbRNKqPff69O
OcXBMiE1Mjz5L7P2fqyF3YFKjgGcUwUE2/rvjmV5/KHSnLKh8Nlx9oVeCJF55TeZ
nV3snUNGeBpvvnQ4FTU5yqGyBwesY8PBJOVXFR56oNdf2AfNuNFmloWRFOEpKcUV
6SS3xNcS2GC+MkzQA4jaHYGkSfWumwDBrCGpt71KlOBL5GzbYPfMtl7L820fI92N
7eb2F5Rvb0+lmvX0N4GsEwWzb7xJpfe8Hbh0I0QaG50a50s1+JoQtPLcqO8ntfvm
F/1IopClWnhe3tg4BJxM8mQCDnV7gJSjOb8UURtBudqFskqro72it08DUWvMvTBN
R/qdj0Uj5O5cdvfrn+leSsfpCFQPnK0vtONpALbNCBjNqcWO9r7fyfIF/Q4bH2u/
zO0yLa8eIuAvqz8TVLu+7Hd7UVJlbiS1OiRdR8/jnLDNZTOheOMu6/Oisef2e9dX
/3NMh+tgu5YlFHz6K1n6w5DBwa3dBtGveSjYB9Gs02P8CCwegWQboea2r1XiU4mW
OQ0NAJHus/GYSiaRe845Anu4YcMGizxuf8RuRv/R1mrwvpH43zfBHKoH7ZGjWMAk
e6O6Fofk0FwGcHck571SzTCNQyzOBGA/YqAN7hIxwvErxKtYkT3nOdcp9cstQrEY
5E7S0WwYXmySEiP39Jj+bh46qNLw3WjNgXKa5MVqmLKLvRpLSJXpLMhQr0uW2bH7
Y5Brebya9UYPMVCEiX07CKwg1xZ3tNExUK2GXTt/PjxA+QFEAZCAs8NhzYQtvxnL
G7yUxIR8q3REnjVMN4Fw66vRFNk/uVnThJ92ToeupHzL7a9OukyZ34lzMgLOS2RR
02cn0RygPKYnADQGNYbAhc8x7ptKmlfa5Xb5wBmxtJkexwF83r6I3uqfokfxn3PK
EvEN6DVuYCN569aJWtTdmtCmyNgaOGYZn8+7WTu8yC5E1FMhafQ37tbOwgLotTQh
moTzieogzNGTwbrQ8mdr7j5bSHGtUOrmG4kPU2WMg+KOBtEIz7muldMuj+0uDJpS
+MXcqgTdx+M1ERtj9CSRwC2GyTzIW1Gc/7SFjp7mcNZe2n5gc7C+P+PGRF7dlndK
7SZrLcOxOsVgdo08xnQHuC7SrqlxAWX1DErfbTVuqEUCIb07ZcCouACJWUtXaeR+
RUorSBI6Mlgqc8Ntjgaop4bGw8kZ/Hc+zqpxRZISTmnYHeLNorpKf1n+GGqSZFZX
x2Id/TkHau5PLZhbs5BdH/m4I3pNyUAOMOrwrogVicnnUDz3uC40wvK70ibP6pti
CVWGq9r6jht0Q3m979a6rtVsoZoDydbde/LqehcKdTYyVtGH1ttEzdVjZN0h9K4D
KqPIZXVKWS38PMJXAXZM7TaLQcXDBogyBSM35TlgcylDOenozvRokZqOVOeD5wWS
yQ9NZd4tYKkbpoC1lxcrNaOFYdposIWW8tyxQvWjsS7l8Ya/nFG8KFOiEEvfkFUL
uoYYXbbvME44o3j8VGaVghYZuGnV+sZepNF1jub/xZFmCQQ8XxOIIFRpHWv10E+E
NFYx5GX1XAeYIML9Ho7m5x9pKSXbyTOvKKc/EDgW0VBn9jDCSbmLzvHXFyO8srN+
L1TNoCmXj4eH47a0dModZMGAOVFu46+cyIcHh0JCE86PuHwaXvpHWcc+vX6/iRJC
ITHluev+hsbXdnCAep/fnlAPf6QCQjZxyopmxODeySij+g2KFQ1GxAB1T6mv6EQL
uRiHj1HsFUm0pHb+CTFxTtcpMuQpqHnXxXDzKfJpiNZZwM2pOm7x8q68vkC3oC6w
2/4+soOm92fy1uaHnhnk6vGsX/eKQTht1gtiBojpPPscEFcKRkyReJqU0IFA1DP2
kDtDUP07P329LT2BdxnL7AcDZYu8AaA7OilGZ9wxEvjRLmSUBDZr883u56zlpC2G
0R8vSCt5Mo+bMqIIpNpXEgwB8uaDLS70nytNph4gcpAKWOs+uYBGkTv9joBYCxDO
BnpnFH6+MLxVfDRtMzgqMdt1sBSsGmPQJv4XcqKXoloIyaI2k5BeEVK4qZDTNdlU
+2sojTmcA9SmGWTqtb/9zqooGkAPcqXxJtmw61pzkWz0mPRYLqkKkQE5HNAgGBfq
zpli1MieFLmmyw4c+9nQupC8k7Iif/Nu/YX9W70SyWUR4kLV4Q3UG/pPhXAvwIUM
IZQnXIkoGM7IQEaMdbzNGZBFVO+ixQfCKWMdcv1OD1XsvtU/4qI7SP6G+wgf5/NE
objsA+XxabFv/dDJZXctlrLwI251PPOAGR/UHO8apKb+XrsW6f4jXJl3okaQ7uCC
wHVNQxtAZ1gCTb1mTfClwwsOAlrXpf6L5QL88rwvkyzAW9rYxtXrwNKpOdxk4OmB
BeumvDnwWttJiplTofpnORFh+SlKceGy8tDFPG+/zAVfAiaXsCeXKZxkcd/azCnR
E/jS/E/S4ESGLdP1HK68D4y4fDxUs9Pw3+pI11OuM6hnR1ZDrrgSLyb1643Ufil0
BezRNBCNMn7MugEEZDi/ql6PWhMhflXfEPqVvKgfYIKRCY7zqf0/mgd1wTR7ZAcu
Csfpl7ZwdW+T0Oczr063iVoTEpfFvfGIsbgMFCG7+BIGDOgFOsM920Q+Wa3nGeBG
visloxIwo+uY4AKYfXDjonFhsQuGu9v8G90Fsp4TyFCjNpINgQOUGFtHyvFnRYWX
jTw2eB05W9b2nRb/+nxoAy6J/6ix+KiTtMIOB8iwEv4TCIz0fTkhEEL/RBOMKrPW
WckMGv7AT+kt050Akenp1d0f5o9FoW4VsaR08Tr1udtlysD70H3HLXjGePuXdTe4
swB0wZ2tAXh39GnCVHGFmHosWc1K3BGrZhyf4gP+7aQxjUs+3jP8CYQaiqj5jGxW
I2zzNHPiPOJfC6KLJxUIkIzky+5AUC64skGKit0ZDMpd5PLxEPc16AThAZmNhWaX
EgHgWnAeD6NobasP7xDFi+j3XYKNZEchFc+bTVmPF5VMWLExZqbjF7Gxa1OrPEDa
x0BhbHp/29CWzrt0dmGNHoJdnHsxTeLAZ2eoCTVWO8O7eWh+RUSRbbdhbKmnZ7eO
Nb4wqcKQUvSg2APbZVzWgfWhA7Xa+ebLZ4xhOyfXGVsCWiYjkXdlGe/JC6qHhv9g
ukZ1Wo+lIh/xClMg2NO1LnuZN2jGh1IZJs9D74l5sNWTS/iDdjtfe4M7wzMQk9UZ
v+ZKphY5s9ra9GMAWFzjobDRstEjWrPI+UX9Elt5h+lrfHZuEqXemkrNVM+wUBSv
icgJB2p2lVHhKDR0FDnJZzTNJK/ucJlEF6ZvbMyKSsuSOPoPl6c2lhRbtvkx+H16
PyISllz4PYiRcmNVy9LSWkYh5eikRL0WWVj0uUR2GwImwOMH2OpEtQ4BOnAe85Fp
12BTxR626+kHXIVHt6KAS3jFeNCDxCtI/zjh+pIZCAhjQ1Y40SweXCMaLmvWZiPv
gIbu7hWk9KF20IESoguJekIPDFI5KxSZgW3764N3kaNJxsbkf3Bpbf1/cOGBqRS6
RhGSAhFdltziGbGVStc61AB6mRwGPenjUedf0SiIaAV1oAfh4tLcbdvJNq/XfBRI
F+PGkgpvtUpnbLLAdoK9pxPRoO6HdbgULFXMbFMV2L9l+UN2fH6wcndQIHTsEfQZ
SLFEpP/GP6mzdvM6jpB0OlwyII4w1n7HhwsfcS0as/3awdZ9CgMx/vBpFKh9L7oe
TkiYLXi7rdG+tWtuw2A3M+GgQjzgmlb78vGV9F0nIKsnBv3SFK4BULKTtflT4m1x
1TMKmyUed099YXqf9Zjr1pn9VANhFxXO3HL7vlqH0wEmR6qAe9yzZyt5Vm9rAmHw
hgh0dLT+EkhZFTU5OOoIH37GarWJgr3B1BX0EB4oeZOmMBi3HjCdUpZVv4/B6m1A
aLpKT8//431zlAZLg6cEAw9JtNyZdQ3mxgRgNLgqjZckhhvD+6Z+KylbKxE0UN58
D6CfTo6bjSZquIQZsYqKsVEVNUSBh7RfyYM2O7UPjzgb9n7YklZKJY3GzreGW10z
pJR1PqEmRiWipSH3ZMsK0pMqlnyyaUmRBHYGdA4JJvTsm1zr3RAttCZxj1iJyLLh
j9UmKEGD6qJxoCluE7sOeU8oQS4d/uYXEk+S0Tq5tE32DcQjQ63p4eMUhZTvu16K
LjaxVeg6sluWS30Jf0ghu8Fn93Tjlk9Gn+haUc/1FjYx3uzorCc9WJmjNib0CFJq
enMBwVId87JjptZoWp1H9SRn80G546w/yGEhjXBfBAucSU9are8F8sColqfiIHL6
R47RTm6IlP0p1oEzoPDVSKVaJ2QoeZB3FYOi0eoX5IlVS4vrs5hpZS1v9QnAaANl
Qi17oaims7i3QPhpcbfRki87oVAGZXUmnu6gaOk+vpkJ2C8spMCA5tqcne4SdBp0
T2w/U322BhmPU3Mjoj25asPpJjIRK0B9a2DXOhTFEgC/7i8jME8ImhgsuSUMQObA
8dsGNAdw0akgxu5k7CXnaH6IxiMmEj6/0SQHYyxZvsUZZON+d+5msxmWYvZVpHJ+
JSWQOJGnKo3XumTsGr0dWRGUa1MLCfXf91ZjEP2kGEfiOVoa4f5HrqWzWMvX8nmb
tz4wYtDCw5hUr2PK6zBbqg+Xm+1zTyS4yM1w8wRGceLhPu7qFFdbza2rbbVEiZnz
R6WxQug3WAQadYBLLJ6kQ+JmYp74fcW8rNTz2O9/mK/BzRRLlodDKyvO0eJ2/uy6
boLGAt09oj6N6dCQXYHW/euAf02CT4W7dedKqtKo2ysp6vI6QN48uVk7ySnPDxmr
XTN78D0o+v68Nyyz4JsYn+PopF7E5RYIm/pyf4z63awrBLtA0smaN/M198IisryF
qAZVe7Jyqo6iGg+4EubOdMPeIq3yqNUoNbM51eF5wk/B2xTAWZ0gxyayaa8cOovh
MjiceXJsekSaUXhm/8EdZM7+XOdL+EnYh5nYDCQOfDm4V39IH3r6mHO828DyHCRZ
ByGFM3oKF5h+rARqKbB7rbLrCQkls1c9RxGiAcLjYn4QfEKpARm3genM8seQYOTD
WnT/+jEjhtZIIMO7IcgF4qF7y3D9mNkk/7PUmM6/2p/0fp6lEVq3i90+vW6u6/QF
2U5hpS/6/g98e1GMrZwHgm6t5RnJluIrrzRcy0mjX/nYkEoMnkG3A7WTUr1RR0yN
RUClv2m2yEpMEqTf8IqK2JsURqwcOXaGZoJSPUzNS+O0PFwkpNA1UxuTIRBOBO1+
NO5geXP+Z4JfhpFA2oS8gsny7K9nTLAgBPWqyRQDeQROypAgkia/psKsRi+qIA0a
M2JT/A5oxgqqWj2mUJwV6a3yPvd5Q+ezjEz2ZdFH4xHOMZQCOG8paNThdmPUI+jd
jS7V1bwm++nlj32bK3x5GwnRfaqI6yezD0KKwpaPXl6dZBh52w8D8edH9Y+AlfYZ
RVYG4wMmqbRfTJxqlu4cePwMZI3hggpb9m2ApPU/+BXeJmz5hh0cXjDnaZm1+FQI
zdBUDD15SK2IaG0pL5z9ZdiRSOxcd7L9vntGtnROpguAnj/rxKDEuKkq321/fqK4
+Av2SfKseX7jSCyiYnWGsbajP2G1X1MAzziaz5pyDPOY6mX54uRkQuq4LtBL/nhT
/oiHkQgfWsSxl7e3855J4lHC6tukRjlDuNEE9e5Co3+o3HC5tDxVfna3jjzcwm+X
B8chz86qRNdemvJjRCzi94tU5GKVQzpAQTUpyp4PxfSvn0R4g9hiGkwzBJw8UjlF
K6sGGbC7ucHuA1MNeYJ3P4P+WvQeCgw3a1aL+3+pHAe5o7bWJ6VPzcXRwRQ7j0vk
3anjFHwYdEr3y8fwQo1MRI2RjoXHmr6Icv30pYyKWvwj+sQlZsvDjWUJs9+yYTUm
PX3DFnNVTH6P5H+YJCuz1NOzFHjhPbar7gtt8UZQu/ZG8oxcK8em/VEZRrBuRi/Y
tkSb/B7FrGssgVhLlcppI6Fc1WGcSJBPUsvgBEvoZjIL/hpgJriG3NZFfG3qbAzl
m5r39E6AJCIC+UR97HJklxGC04FdjYzkMcXACAIdpFAHXeu7k2EoVtPweg0ws6Ux
5f5S/DwAy3WQAIzuJddDHbTMED/AcsGNhQcg21+MZp/KDN0dNVmBcBFkyAWzaA2W
ZrZtlt+K7l9OZQXN8TgPMaV+YflID+AUwwIFffBEVH9NrJAajTnfiHdukcqrcAG+
Qt/L8aSpNLxt79fsUIqq9PySWNGVBPKdEvqhVY8/pbVWtgZjL0ef+0PNh+v6QARI
d8rI4MhIQJMQ1+OdRpwOjN2iv+eM62rFVJrBwqLGUBZl5AYa7Uq9OMDck89BOnoN
JDZC9fm/5/KgPmUyxtvVm+Hw5N1Vpvcr2G4XU3lE8bFP89xfiopROPwL+o2VzSsh
QBQEC47p/IOC6Vm4OSLMURQKLt33JaCs+myqNzXuctQ7furtdiYOZNeAHrbT/bNf
vCqLTxlz4N/jPLHPi5nQ8/csmKzgJ0qPqjjvrE7/kdq2Yqnmxua6wPvrsY/Rts8S
V4o8n3eScktV4H63q5m5h/c4duW29kfsGfJ85zqQTG1zquL1U0aZbQ9FHuKnCD5h
VR5BLPE+A5mFHI6f8r0smJXNwEmPp0Sl0tkTrhn1rcTXQKgVkyAwe3FN2/lYENEl
Dm/NQ76SDJejr8fco19ybRCmKaGywa6rMK3u5CBeO2n4PJCsAJfE0aNLl4MvHmPw
C2lUkRZvGJvqxSV6b4kd0BqeF1ypMMcUBDmYMPpt4CDGSOqWK7oDjEdhX+Z2czIk
y1Wdpa9TWxV4Lq+jF2+p03BNvB/a7fFhorQZhocQVgOTPKPIIkXja7TRT6XJncgc
goyqYS97PlbrqOJcbg8Xn+fv5ELoNlN4ko2YNGaL8gu9SjSKuvhXIaNgvktuJdPk
ZZl52x3ESqZkLqQlLpYufy0a7BLc73C2ZY3inaSXqkVlqAJeDbBNAAFCydkt56aY
0YRMlhKgbAwtioH8Nv67GnA9z/639Qadf97FtG+OAIexxjFQK9RMmOOkRDE28Www
ZjxOTCZUiBIyIIYz8vkyE12EFcLzKsalOFI7wtrO15lrmXn8WHS+m7mUVRYGZVmZ
xdBCmORV3U5dDWKaKZT+XCMfToSxdXqmRPeH4BjlsUXeMuSHil2uEnh4syZDSlNV
mlpfAi3tA+Pqfgx4Y86ma/HJ+ViCJUM7M7UOACSahCdSrkIZBrEm9bzeD3RpxbxX
RwQvftl+GB5eyNq72l2sVQJ3EgwpgwllWk1aBDH1oj75zxmedbZhmY9jO5J043tA
bYVVyu4TcQq5Fdhs5wFP0LYt7mHCowoKuCQSFUJ7ahqNDyIWv1PIkdS2VdcsFM4X
OWNG6SU3NkNX6kcFtRYHcjN4ajhHPJCPsjReZczB4CoOFH1yZPvpcUb/lykRVh43
XM89vd1rbDk3dS2E8HEaj83D9E45lvder+dtu+DGMJ6cBO1UppVLP+gHqUMGHkYB
6R4sFEPtxB/tuG9v3a18vG+r8dw6FQ2BnlujOiNzYdV4dCCEuPZCpOEpyR5Hakal
Yql7ILWWdOdRv256RxpatkeN7y0HV6E6gotnwRZlqrW2DIvvJ+uR0mRXCi0GSn1T
ZAsb2Tj779bCl3zBRYVjm3vwZRWjH54vmS8EIu4KnU4Ugl8mehGV+0RxjebfIo6T
dbKjBrctLDLVq+CFrHYsMuX6RrQBx/XiBXuOUxsxfdm0FpCdzIVWMGY/dmH507z1
VFMyyuDNTp0ifz10PFi7Ov481XNuqxj+p6JeRA1BadamOF33WjoJXq61gpPrZphp
Z9+grxLgJKcc+kj41K572edRnPDlbCb91tAKUSzNcWsGlKxZf/hnc+crfFRyWGvF
SBnJqc3F7MmWf88npWjAF5bF/s3Jq+e6u1HRXmLbM0+WmJXXLbLJLprBDI8qBZVr
OCNp+ZXpMdFNdWvzvpg7uQw2EDrsF8l1rzs1aI7VAOvkN+AaKLCTmqrQNSxzhzdm
aX3DOm09AeihQ1SMV3C580XaeqWSDuKw2TBvySqfnKfPSkp6XF4TkjSz43IFkco/
DIj4rv8WIW20oOk5nKwMqJXoq3wYWRzOiDAL+hSSuKmtLp2MqtMoqz96fumsQ227
na/GcoyhqjCnlWeW8dsqVivd1ENw5CHEtvyQGlIyplmDiaysysU1aa7CCQ87UkxD
VMgDeEBi7Ju34aCE0Ogq9nPFxj0H3poUFUfhgVXnIpzhJrTAYBRIzlMxA8H6vSow
kR8Xr1S+9tTCmM7Jm2d83RaGkr8Op1y0rP4EU+04hQhv1BENP7s9xYY2RPtSMwiy
LIkOgyaArAJp/lOW3bUENOli0IPVUhfkGk6FaoELdO8tmbtDJjiKyCFAznvYF2d0
GIqNXSgDlvWuqKBiiecMuwgLwUrlJIRislknNaJ6mA5BXgmU8skYdZWZHlggR2m7
bU2eRG2xQ/NMGuP/9rl/AF+rorMpHDRjzJVD0hQh2/Vn+aUE+SHfkpwfQUKu9V0F
Mz0gLl1M16qXXU0jiDC+jx96hpXuxtedtlKAtQkQ6DlHvvO1vLBAR1DxLr2gezMY
AFq3pEHCRWYolkEWcsOXcS4JpycROc+wFCxoEaM5AFOh5qYQNLiGKpG/SucvS9Jt
etpL8qgWz5VXyeFjSC8c/d5aNB5FOWxvPbL/N2gLDi1ZtAGiUah5m+48ExaeWHZ/
cpLtID1qFAez0fwtK6FKuR4ZgFJUXe2U/l3iDNAg48rswdebUNjbAHdD3vZhF4t4
CkEfDFisrYAzzTKkKr4sNPhKHOu+GVA1LwlID5lw6AtZBAmWBTjfVD05hDmandwO
00bpfvkqlNZkqRRB7vCuiUtoHd4MaUzF1uXv/7YMpytJe7GhF3TcV8kxDt9V3AP7
UUpjF4lmWgUVtXRyshQXuKbCXA0mITc3rl8Js8DzirQdWz+O2OmdilkLw7Ahl6RB
vTmY6oEzGKF6t6mTMy2Pws8vLwWkZfhN/vw1xXAzmGfougwDWlAnV9CJsmHBcz9c
RQADWNhx4Gev+PlYDw8vx2fUIgrS7cP5FG97l5K+V1Cli4ooS2omDEYEnc1kN76O
K5WY68eihb5C/KSv1A8Mhpbx+YnyHpuTLmB6LNGZ28NDyEO6z7bqBbMJLHG1TGXT
y9/a5JZ+1MdmtmOf+Q+Z/IRacNQf4t4x7f4UUpFLvgU9oDObbhY+TZt3X4cQ6qeR
H54l1yndoS4lD/YqhdWLA/WA9GG29r0+Fj7AQRknYperazNwnyywVwDwplz07eaJ
lfK1PyOe4DKz8bxI+io85qRTeySVLea+FBHBF+gok1jvYTFM7TieJR5FVNP9+GKh
YATxhjUl9gHcuNs9bUrQ4NvYaNBs4P8ZFnSfu8CwrzjdrDuTm4Be4FJhp1UHPyuG
qHkhGOwp8y5FlyUwjeak5IPbbOXb4cMKif3c32Q2YVbY50B/Y9s8J6o+jO43J6dr
Rjl/V5OvbUOoOqsb8u3bH17+FBOvdsgdNbRWs5Q5/h87qrFa0spztpj8SGilzdbV
NmwdDEUNbnkkD2+p7dA8bWN6Uzt9Qw8oCqMpWarY2w55fuqdU3HMiF6jzO6jgMuw
73JfpFIMbbi6yFjcWg5wJyQePSPpf0puTF0n+qcHgsJ8iZtKOknB2XBFNEvolgRw
f4PWMHYPnJsFU+OFaGFXBXehI7BcyCaLlHUQWNFEirLtQEq0qF4mbQItIBtBh9K9
MiBBcrWHAz4CqH8hGzh3oN6D3cQYJ6dqx1cP4VoFmdYigCMTHvmJKRyjn5t0/iYG
/VcipbfbXAxMSLz8Hnyq0u0FR33qIUdutukU7csnKkzFW4KYianCkflgXSB05ZbG
ymPNDNUWvxzMseelyfwvvZ0a8SmEb+CrTZh37S9WaL7IIBj7WIxywCFsTgl06aou
qxTYewXjq1mLwWqrDpXrjSlkKT0Wb5OedhD/NpDwCP8WqCRESfjke+MZp+fbdL79
JAZpwa2DK6E2MxjdKuN4mEpe6YnJVvLxabEmwsmv2RyHktcobGJpItYfwGL4unpK
Ujnanopi/oSM64S0z+8P99Bl+ZMj5PZua50UxdL+0xEOGQJj5yTZ0fB4lbnzmP0r
1h8LSW6MRuLm3Q88IiXPP6gR1s1lXfQttpOWuZRxpS773EaYudbFzhnBtQ+W258k
6j4ILjSiN1EgDUAhXInde22KIff2ORSQIecwDj0qcIu1rjmIpCIv7uagbsm4TxHv
1w9+a+eLotCT1Ss/T9Xc8bGQGc8qaWR/o8IE4Y4sXcxmX/TyMdG574xtBYlh2wQi
qp7hZV3GsLCHfE1zO/6xwDAsxcHgXzoG/xs/YLQ0+3CvN9fJX4050r516leMaNHU
ZHll80LFOCHyiGDC0NziwZuc9cXoJrpNAHS5mMh6uGRHGUZZUjWff9HVX7Z0io1l
UbBWGCG65R4GO7PC4pvLH+AlfYRaOelV7b7/ZT//gyth06mKJR8Y0Cc67PU/OICw
iMcS+9SBhCtavO5dOI2iXT+45DGcbrbYEO5A/6F/V7cRJWzUxpcCK/c1w5d3/20W
JxYNHzSDaQdN8b25KyDwGe3tp4C8JyVVzsNgn+v7Jye/KY+fJXaLtC96dKAKUKXA
aMQeGlhrv0KmCgi8YLkhQWMCwVymA851vvPMK11CH68s9iNJTB8J6KyLkEwOoi4j
ZCPOf+5pBkwYjSy/3JNOI4kXQsNhrgrmF3ynwp3GEieOVDoeJ73UGkHNQx7w+Qsk
SmOxXx5E7Meamfpe/LnvhMuFQqoO6RgXLy6+oH/8QL+qLn+3hXk262Et9i8UCNGc
FmEpjYbhBGs/cYQXYUXI39rsKuWndHnipo2mX//flYvOp480gkeL9bCIM7UV+u+p
LXtfryB7IHD/GDAuv4aYOI4XO3XanRZ7PDep4mizZ4QUKyvldh9DZRaJ3+jXeS0o
Th4IvwDC9JwNtYgNrhX0XD+65ZdaRnUZQyyWPzyzhcXzKtU8YRAFDfqsFYZcXOZj
YVFcc7GPE5lXbBNTNCpxfn1hfmGSVIgg8T7i+1LboyrlKVnVNMniDwdawK84EeIM
Ez9racJVlz/XDQ0l5hXW+FoZV5Xp6I3i7mTqdEmWvesQesFGuFtlroLEVIiMQAzD
xqcGyGhVBBHC2IBbbTIcZn5QCFfNgVTzsQ0fWOG9JAZQrV49hsBNvR6eV/5m6uQK
OSkliqypJ29taMmhuc66pz08yFBtI5QaTMggSWbgSE5JF5B0dPxT6sDai+iE2FX8
7fJXYaxS0GCiNufXVJY6JO7ttttfOvfyts2yGq91x+rzZoVG2X1pZcqAlJBU7yNk
Bf+RZ3rTq94AgkMESmfC47VX047AkoLlcwknpJzCJkXfdH+JNX/qeDut+BwvS6zw
NCA0/9J/ILp6HeCpt1iD9uW8jWn+rV9+E4qYve/1kZ2v3unDud47vVTMtHxKKJoT
/pKKUjBEV6nuG4HCwVy9AMn+EpT1H7V8kaZqcOuRPXLHlAsyuwgeZ8Asa+c3TDyX
KqZ93ZcS94ynnWrUfT35ps5ltQIZaPXilM0ekuxvlASVY90eZUaJdr4KS0ZMJGEr
eNHtgwqlNCAFe9pO0ai/nnbnm5G0w+VUm4wo5ACubGilYZGjWRmwbKMuYaOnFYA/
GkyqXmDnkMH8IFCXb9vflYmbdaR1u2vYb80JZt0Ae6b8pWptjvEIENFhZnuONE2o
XZE9fWGIdf5MpTqoyDmDiSTIWZrVEyaOIKVkSk6uioSBUWUokiXw1QYM/463Msh1
de5JIQx0bLyqY0wkDnUzb7fLv9Gv4aJSWRyyN542Wy2h3tHbrlInUUhO7g1id+Ji
C3051J91qT3qXsiDnXxLlKeaOg8M1eWTl657MHWNuFmw/mt4K90L4+cq0jR6uYXX
g5aHFF3n+FBVHXU8rd2oRYg/6df+GIz/Ud2ZoPccIvX/p29lDxODpr6ntOa014Pt
eSoCCwJPy8x+rIBbqSP9GPQevD02wX27b0I6O1vZyF16SiPGkIQJrAuyc6h0oh0v
Tqb/dF5aHh17m8dPWYcf2fMwfNwhvKgPDkg/A103vYmb2tNPcO/xdUjXOEt9w0DU
1EtZWx/NQtn3fQmWlpLvjLHiyWHxbj7ngGosubtZR8EjP8azF783iJ6MbNS3cQ+q
+UXDIXowiDuZAOCz6SowcdQzLhsw/4a7D6z3VGpd14YgFo9T+upTeTDdUj9WCH1r
C8dmizX/NSZX7kJeRYE4u85BVZcc1Ww3EoHva10LJzgKG/6ol0d/NLAb7SYrvgmG
ID3/1JU9U0DIO95VgJT8mreTqCMoWCOCEK150X+PoAGr1ThC163NDZXc/yCyGvK2
eq6Bqu/KhnwskJwAWY+/F7mlUky44wBpmbJOLDmpcNnEqEhQKpyAD38pKhW+qcVQ
Hc3VyzrgAZXsIWdugWKxJ+cxUnHkPWMg9oACp4ay/qZpVHSIuZs8Oli663p3hg4Z
rhegCWG29az7dkzgnBP45XDjDOxEI4+Ls6t9A3W5NtLMcP0IopyqfBGW7+Y0GKZd
RdO/6sDXidMBTetDT7586v162+64i8Q1U2YmIlesyG0nAAW7SDvZaSSe66+aun27
TiA6II6f4pmy+5+/fzg9UXqD5P9Tr+SVTY/eSb9QLyhXwDPy8CTCcCjiC2DJKf9b
5viCtVbSA4AYojtdmUN8Lx5Q9I1aDFQgzmWsCmWD2ahXo6aoJYOlWUf2Qiz60Ood
cNJ+07Zo4OmgMDeJJoybyOYFkHw0PmzAhjQhgeftGVjnKXbEisUBAzviqKqbhBec
yxAINzwqXPihIrglSy/UpiyynUMfHmGMDzdiLyVQYFiF1oB+TRQOX8Z/CdsxJmdc
Uazroq6ytfZ4pK6NEOfPwGw9UsoIu4lNpG4MM/0z+YNejVF+OY6w/NfTHNG0caUi
VUn5Hujz/6PYDbGS1qlDg2USD5GDBifrc7JiRRJ00gF+IvkikSc/C05G8hbf24Jg
gZTVLFig7BAbXSAKqlMEFIZsMgToKzD7w3NxuP/6OdTJUbF2gGcgvv3JvrNBLexs
xgfl/MP3gjDdQod4DI/5e4uEtMWJwas6aLMs6PwsWw50aJSAvhLZHqSri/4A0+4b
aoGY3c6xUkteIjYvqglw0WKVnBSuQocn9s6Ln/elFCjh0WB9U1G5B+r/GoRjMfCr
nd7BVTX8YSny0aLJNt4C4YVFVV1f9ZLjNGEJ+Zz+5kB9OTQeo3B9d/x0lO9DOwDM
+gYT+Wdgb9kVFZd15bKq1LzfHXKEJYh1FAU6oajPUcMmv2ek5gqIX1Bq9ghojVut
3XELuKPSIoh5gmcJnM8w7+D07LYQJ/VGJoRNKQ7v/cI9HPIekCOd40MQW1gSCQ8h
Znqjar7BvMppTTKaw2Ufb+pOPA9rTuCKkDATjl6K7uIfccmT4RreJivkOjL64NL5
+ZDB3LZ0ocx+vPz4jR0wOQxapeM9YXD6W1qY4nxPJkcuDBMe7a2XXwpiJl1Q3ES3
CcNbYk4HNcwAOLxZNc3j55obbkcZ8oY+byMbmj30FwfliupBh6FPZJ9ybxWnz+XG
nYI/vf7IQd5H38GDuGil2o4siMwGEJJXPrfXxxYrT+8qy3YrKQRDWSbkL770EEaJ
SgVuZW2L9pPkKMvX+CqquF6kImx4WOb9uctD2Fur5TYIaZ+huYjjqv9I951ZR21o
RbWCmf9nFbNXM3ROJxHrbzU2iLdvqS8pJwE2z/g2V9AdJPn5SZwF+Sxr94/knPb+
pstXl10MqNqPXBgXmwKXVsxfPEVbUEj6Qj7G6OhfY1LqMTlwU/flLjmqW4Wbig87
DpI9/h49Pt718IRkF6kJKUjRxzDjDebqHSBwambNZ8oOltakHNLo8HbZLMKOx+yw
HPCHxmfGRFEsJ8TEcmO+R4IVzn0uw4+Ic4nFO8lzn1LKKe0HyLql4hgi5F34OHnk
pvYVsEg5ZJdkp8DuxuJrk9d/1fk2z5rVZNz2je5nLPNWgny1K0ZepdabHZgkk0XQ
yhVULouJcBk4pN0vvuDzW3N9n1ZNWVlITzbKVwR/x1v6KZ7c3RsjPW4DTEK4BvBV
XEhO6PbTtpPHs0UrRFJYe5Jwr1AIDpGdXFz4uSQy/gOOqS7ZCkx+JzCskowP1lRS
2WvEo8/sNEi9SwfZGHYmVF+DkGcf5XxwAomcVgCFvj3lOS7RWHFicADV1UitFl5f
R5Javgolx6KoVC3FXKPWb8/GCxR7rAzwyrqZEIjSanEOUrkJmK7x24LzdrdwsfxF
hfVAkiu0uC9gaxuq9pF3hiMRm66Ioh9BrvSH9Z+5HyBVRDUbLJoD604rtdr6KhJD
8384SioyJPjNiVQXEG1WAxVImqcyZ/luik3YBARwtdTY1tJFemRh70NjjE92HKz/
0n1qGYLY/fSJ0P5QNNAn3WnWzGTc0W/Hv273A/7rl/S0RJWuU0CP8dI+0VpQ+Q0Q
aacah2sgaafktl9VB61B3JI5ykEFu8gcMolkqeCYwE5C/F5v1VCklncYV7opA5Ct
M53mYD1uYRUih7MnJr59ASL3ST6nWnScS7zAFycpGg1zOoMxHZbpLHRRbvsquEmj
taNfOUJPlKqfdCI/VQrY9YhKfPTLVJHfOZ5BAIwYGjbQMvEBtJ4ohLIH3GJpLE97
J6YoqO1t/bbCXB1XAtmcZ4hXz1T1fKjacShUMLe5bfwomZQWwAOd/Jjqm1gOMxt7
gNnjj1G3Afa9p0AbnprjgS6I0jkSKGMkbjl3OluRDcbd60zcH3oH3ffcoH63wuRA
D2CGJUyNShQ1RWQglBAEbkE6eU5wdslzDM7jEE0ldF6yIMCuJhjO28jIAv/XomOj
xDfCDhTztUxUKCe0feLvkoth59d1M2eyXjCctpct7aY=
`protect end_protected