`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 4112 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/9huKRhRMtvnNqb3Z+UU7TahEoHV+T8U3P3ufru7l1O
3DlgtZzb9QxCbOjthp9+wDkjygH0eUfDrEl1ovhZG62J55FGE/WODgZGKqQ+wjB4
jqF/XueiOUeVZQirjioaYzoJV4u1oCRDaikKvsUh8gKChfF6vTFPz3W9bHFvpg9+
dAhzC6E7Rbs5wLQBxcDRRP05P6lzcHfXLsdGXx3yqM7QlPBlyH85si6MAdntkvfB
zaxy5IpbCk33lHdqjaTXJHLX0hTIvUNz7pDV38x8IIHNVegM4ogwc1SYYjIOuHj4
YZb3lR2xoEhV9LrbTHZ3T/Ahz41zC6tUx+InxcUIH/XDYj5kf3kBI7nNDlvbL/4P
wKgjTUhWTeBaDpuCjohmsTRqUOF6M/ciaKFd7VGH0VN+kr9HcBh1gVdjS9U0Np77
dtnjJvms+Q/wI71Pt8j9Bv0Wvpb4rJohUwosALLM+ugchV4HB+pEuU97w6g1DfbD
AJi+XXwZsGnRqRmpuC5mt/6fBtS7Hti2YIb5ppWfi0/75YjObrJQXTbujmHzso8t
oK0iqL/DXGGBtJyYeBJcWAk0exF4INhl4VEH9aB4Uv8Kx8Mb+Q+RE/M1v+4TdWhA
p+dd5hGnHHl8B7Z5GIvPZpWfX5OR3UdrRbO3zso8Ox8bDuETSt1SUmLwqjU5ZKQP
ggkCcBu8WQwWzqIMS9FHQfC2rMhnsJtF9BjqT4S2mBQU3tazPWS4X+Muzeo7XUlb
U6YAMxffXl9gpOrcbLtWgJ4Oo7lkX1zBpT46fY4tiYOCWvfdfb/Fci/rOSddg2io
whwen5wVnALFGPCw3qqSoAVqYx9fURw0c8Z7MWDWq5zdc6qthF/OnpoIZHkU80Bz
2S71F1tdCtwYEj4K56oxMbB2hiKAo6aCbgoftpky1pbzAKFbGX/0xBHIMARAsmpu
WO8gUaqHxvRrekGEU+KKqpbkuB0omZ/iDYTB27Dw6BznkfiEEuJQDvDZeV29AJkK
WSWTVsyTTeLoKlHWftwoJDiOL+GzHdao5+r9fuzvM4qu9RKJpGZ13ncEg9sFUbC5
0h0X7sVE9Jx0DMU4P6W6q8T4x2GlwwH1jNR+faHAAXOcyrQ0MqFSjONCTfobJ3Km
p6fPiLf1tGvb9yGpB/cLk+lomro37Ug6EfcYZKAUMa9abey4SRW/QvylNkHN73Mn
c1QDIqjxxTe504BZ+EQ0GkFC4hlD/R65OcWpU37QwHriI/0LqjMsyYU201NYxlts
r0XTvCFewysdmkdxCGgob9QpBCH6YkFyQfKdFr5JYcQEYhJvLevm0jbrPk8QxKX3
vc9Twy/HNmeJo0wbWFOCSSf4X2sUshr6C9KBhlPAxVeDMvhHTPS+Cypb/f2kwoyg
zAcxmWoHv+xXP+mvSL2oY5fu3lWeJGv4CQdnyQXNKp6imXH+sLqtproebDXTz+bB
KD+ZQqVci4pCfNAonLvoNGXLP3FGTMqrYVMfK1IkR/LUKAwK8lzFPBQ0qODrAiB4
ys+zy1c0O6uW2Kefq3KCkloKQxHqkJUzU6aTv97RIBK12L0QbQjsWI2TzBtlRmbE
8nero4uZRXgl8nPURUgmPw8lU5xrl4EK8shKK4SEf5RulEFSf3qMo+SIFk9HLFe6
2lAay2A36nlCySQZCVHv7EJIr9m/lc4TFIEhnfuvsEqlJS4SsGeLHQLrM+s4Uwfm
wJhzaSFuMiZzf1ekqZPTVHjX3R6/9p+K8su0aW9rtK8k+0f84qm0y8q/M0FZ76Ix
aQfi5b/+WvRbfR25FYqt6nGst3GMw3/Euoa8BQm0l3lf1eUov3uvTdQVqzM1LJKy
DSn6KS7U0WMP+gq92vBYyZtYyb1i0q2S3kJt7YUdrGIL8RqW/lECx2R5A6oDBzah
lHmFrHJyCJSikYWmFykvq8nLOgJ7YHNRYKOW3JuRr4Z6ele9U9z5nVOKj+c8Fzq/
ggub3Bxz5g5vvH0Gf16/64bXmchDKrosbR2G8aedSjMmo6J9GjlauJ6xjLQCZuEt
P8tTySfAn3d/uSNKP2ObJzRBlSsoeWLrIzL+NshW2CjTYEuvHYlKUtnQwlrZ+nWl
DHageprUkvzZnog3ByeJDnM5yrPz5j1VlZlprzyXOmu4Sspy9O1sBaZvU6bmVkZH
VYZmGSNP9hJYZ5wkGl/K+vcz6XCql8fOpiZqdwHwwywtGK57BJBW8I494STo9jbQ
XrZ7agV0MRzsjr55eHeQyfUB5SVqNMAUtT0sXTZana0hyU/eFEOaWBMth0BmjX36
L4r9pdlPrPb++C5HYmgb5xlbc3yeFX+8AxW/UxQ1ShpkdaRIY2G5b9ETuZdrimFD
GPNbaoe866AsrOjIXldJN1I5ANw/Ji4DoPxViIfkUaFCN3NOIEV4cvsitjyEw+4n
oSY7Gl5M1JACtgQVce9qoROI12OIf+k3kvV3D++rKkBjwxSJg6ussPzfqtMny97i
aNu1MSxIvOSWzFyxKg6Jk33M/qEu5aFZ+cY5KcU7FS7S0C1bzfklbW1JyFU+WWLP
+CmaEN+eGgYeXHMMR2pD1NyvXe9dBrJNzn2rnk2CwL8nrXGTF9GBDDQ4O3ubq37W
kpU7roX/djBZJvaRGI0rhfgs6SwTKRgySBNI/odEg9YRuWDd0aS+y1TKFL8DlKj2
AN/lMDMy0YF8CnAUe1E2iCiiBk3sEK4zwusr8+IJBGm7JEPQRn/B67WQXl/zdSop
yzUaCvA97vGDx0Z9yluZRNhlNLcPq0fQ4eCYzvdYE3mDFnAzSw7hXFqcFgsj2lhB
MhnHIBvykEKEYxde4oLJCTgYTLPw8gNEU0c22TfEUKd6s5IDtjdiUyPwFyLjKQ0N
sb0A4v2HTNYP76yWuu0xpGEiBbbFQirp1pCsJEvW4em6yx0KozyILFpDySvMSy0P
R4CtXttPwf73To2xpa5xgl2+88I5/lcC+VnwB/Z8Rg5u8F/LCu1tW7wHSvKj9IO3
XtW/usuXLB6ZIeSbkxGJLZDNEqU/G55FOwMEw0MBYDXl46BTAHyroaC5ie4y93Fu
apTRHUGYxOVELtjPzuMI4wskNw8L40H43qVoLlK7lxvqoBhk9MPdngqORiKjBFce
gxP1rSFnqpG3phq0HV/Lx6AMPZ2nQflrPK90DEYyrITw6ePpLKuZHTnA0pjB08NF
a7JzRq289o44UUpWeAx6BZrf8AfxxLz/tRGjqn1etBRWeR3jnORztXzkYByizQxX
wg1+e8/ZnyaNIQt92WWaoxwDMZoDznSZ7BLzRnb+1IRbMVozWjK5gcxUyVwE0Tdm
0xPIEMHsrF8cx8WJKGhLbUTTgYLFowBEQfPm8hU0lJIWaTY5k45Xi7lHIRv2zUqG
1YbF5AzGvz3k+P7B6i4Yre2H5ZO9+0TZClBBq/jCsGciwGI5GkKIxEuW9nUejbK5
7tP/aafmjsnSWtiFeKKTOAOhEenjDNbCdPms42f/dHsvRvytAGKrstk6eyMfS51V
TYHZH1VZyCYLjOeIu3gpyOOvSj+PdfJ5TjT77ytWbyX6bHqRqcnuMJkTjDTl5nBp
eDT7n8q/CQ6kGMn0rhVOkIMFv/jCb/rcRo8OaLqSShv0SX4788LjfC86cePEyGrO
7Timj6hEpt3v9H6oB3i1wOs+Ag4GGSDYcMkhTSyKeLojkfj/m13L39sxT5n9rbSV
A1iKZ4LysaQlGhMjuqxLaW8Y0mSrff2SlqEu6w1JxIt4HzWgTfeYGfECki4FJG+j
fkGrG6TVaKYJmsm/d1g4nMGDxFGkbJvcROI55emKLAZWARmLEblUITP0Pa41bA8a
77RrTXDQvVAYh4imKXrQdMYbTIcwtnfugM+W3+Kbpq7Wq2MzYceBn1Vgqhn50IrK
uERMUbd+jXI04omuFg0PLycNZq2vlbQ/wgy/D3xE98SbmYmXryaCwFJ13fz5hUm9
he8Med+OgJwUTnLx9yuqdlXiLdx9TPTIlQtdeYRNXnV9QwQUohpVaDQtKZwVff8/
Bac5jOGpj6q33j6zglNqOzGqbZbwhUtEp2fc/lt2LU0WSel1e02pYdIlDqOhi7Ba
x6y0nkBSdyUB/JcVhcrz9hzDEYyhKBg0C5YBDrOxncsbK2/RE8APKrAXM6oIAMRk
SxUJMfLhM5xtAwysI+uHNmWw5AM1kEYEsPrwFuXFMok0ilPHa2Ty2pONWOEjgb3p
0QCvr9LyQruzoLf8JuNWLOrINLdGUP2dsubU+xFZ8VAjzXOZjwCDFXdb+X9AwpGL
5iRrzZx6BRr+N2mem+xlxVYL942SmX8H8algjAxOfEFkxOd01sN48+PhLrsywtIL
x5OOHdZmFZZ52Rla2iokuLsOf+HyUQhp4jctd40fvBZzSyG4nh4PX3mT3ajqaF1E
NspGoWPUpT9kemWvd14blDHpuz4m0uAkfeKrRfgmxqGCATatxnv717gUTlRPdApz
oFiydFYz7Qa4CZ6rx3xSPCs/LIsN1Y3y5qbe2Yewler6P0ae9r35puJsmrwIjPf8
uf/Ju904amF3plWy2wzzyamtt1JuvxIdWxi9XBkyP7Vrbld/t2WGK4PSU2TsKPEi
gdw+w0YzUaBI5q9BpX2tejxRJVknGPL/GlkIvo+8yRkxE+ir8Ks0ZM4P6pXQCM7Q
fvcOt5jDjuTcJ89nojqWKsUPu3pxhvUR4dRKctio7SbrOshhDLOy9mM2mn/thICJ
vKBzO4l86Ey0KNQjiB40Qc1WajqNeYHktPyFPQmfyry4Vii8KuhpotjLdsjV/PDx
H4ytGOL/FwKSt5SRVv3n3W66+F8OC08NFu90fHAscqHcDGWFw8OZeaXuWbz3kCph
6E+5dHG7FZBF6CeOxCbYa1bctGYUZV0fkOQ33nbH6+WKH6Ls4aOp2AFytgjfX+Of
zAOWm9XIA8guPxv8CY/uZzOizcHy+4GA+6PWyu57LMIzVN8yaizwwPHhP4RNygnv
DbwXXEZzTCGPYH7Y6/T9j/59uzo5BWjVk4mMZQ+sRczyO3p7lq2PwkN1AMhescP3
Nf2FZiFgnCOXwF67eyBXQp6btZ3+nrEBEA+toutuR8yH8WkbD1kY0YRj4FmlWbOL
kboAYNcDklB/dvL6dwMkvftGrZfKtODU2m+c03xLcq6e0oJ0NBozMensHOwGwaHV
5mzFVFlknNuSH+Q3b0FBEMiJS578o2Sx3lDa+PtnS4eQZ1gNAtQC+3Us82tXbasZ
1tWXfUonVQC+wtGeYrLsIrzzwhL1RamlbAlyooKNI/ymFRo2jDFne/7hcaygxNjn
3BJx2YVZxtbZSjftJKlSbsAN1PfomT/FUvXf2di1nn3nyKqMbbyescWu2Z5ox+iq
4GAo0qBdysOBBZQm23+UXeoGjMr+4AJ1IJcRAM/1ebT/jRAl3tJIRYn6qd16Fvnn
XuYq0/vomHbzP9UP0gw5gTMjPmveiYiQdFuwV3rBepE=
`protect end_protected