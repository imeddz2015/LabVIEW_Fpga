`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 2448 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/59UwEX+aE7FohaWu0/8IpTj7mav863zUNIsgIH2BWb
Abd9opeuBjbGF/waQMI2vMJTwD1ie1YueHc3nSNpEh4OXp8P5ybZFY89uyGz3ztU
W1EsuUnchJoQgbHZ/sLbgtGRgsrAFn+ZoIeGN1d6RAGptBAfb8+m5Qh3/nmmBWJ7
TNr4fSxVi9Fc+2BiuGjk+5459YjsJvqmcpm3NRJhx9GePCSIJCKV8o5rwcCKcgBU
sXxNBkTzaRNOkRfzRc9NkeGdfMnsfmuuAlwKy5blQYKtzNF/ZaUfVPjXkLOp9tHQ
wwYaxC0nSS/Ve7MWzv/fICB0WActhIDGBwQNYFHFUrGMaLj8BmuptrpK2hlzNxz4
kTO3ynUum1tCt1yi4W+wg8U7hyISeXX1f2UDkkP91057MM42cQ69glnMYSN9k8qf
mBxqCizYssn5mxTw19GkenrgCj8iUisdT5lut99tMHSKI4WrF3tmua2hBA5vs2C7
DnkJqqvfv5pEV4IX24CnxAFBEryidohgMlr70upqDul8FT840cBlc7TiE+upZS2q
dk6yHKZmSEZLhsh2SNFQLvB2EY4+DcU3h4TLxQ3IilkxgzPNsrmRsfIjfDV5t4Py
sOVTnYUxSLDi9m4KyACXJkVS/Jk3dipPiApfSaEZhyXQBf91r6r4SVn2qmVyf/uN
DerGE2n6GCSJt2z14DXeRo+vHP5+SwX6alVqt7Nzn0IHE9/ENnnRffJM1HGWe0zL
wHimqYgouihBQUUa1ewrxr95AfRwPrv4Hc9SNhSI8BhDolQp2Ovw1dgnyptaDeRJ
VT38/HMJEiHoh0ENuJLZzOGH7Gz4YHJZGpzjUaq0IRic0DmpDqHcB8FklkZbIE67
9/tgh2clAOzBEVQZBq0yZeovyxu+pJxvtSgwN1HexjzA4vlzZn7UCfwt0i0AxwNz
/RtK83FAKGPCIQg7OEYUktsTkJ9SDumSsLpp+cmPxqjLfaQEyumre+bIhw8YivxA
qSvnOI2k+gaSvHm1vzGRR79dHS9cDfIg6jSBt5Zj7CPrN4eP3oStz5M+8kEB3j/d
J6wOJs6AAnzU/x45vu0jgrlvW4vpEHEI27AzFFjqyhBOa0l0OCahag/mIX5cVlDm
CF9tV1n9qNpmxlRc3CGPYrsO3xFN+b0PEiKJzxzdM1V/hc45ZA6jPuSizICUVZEU
shXNSKIo+NLHDOmQ3W74Is1b/2lQs/S0tKNt1IhCQ89AUTd0R6dPevAwuGl1ToNs
ecGF2JVkmIhfVCyzPCXVGhglnGy1DwFkCSopNeYVMkbeZn4ATveS+X3eslKyRQHd
xU+d8bWJmN6tLZwuT2Z/q/HbTldCf2HBAwrBzEDsjtuqgd3Vgf/D7XGew0zueFqV
EmsRmzAFNeAlNzQZkWV0LWnKavmO78wOI502kDJtWx15SOhcqSgeD9u0MooJgvFT
1MlCcLIIGQMg2RyFhZj28Wo2m2pV3YrfS7Ean2MoxZDUuGTC8g0j1xt8gxLmKAsY
Tob2iV2l+sO3MgybYl7DF1SyB3MmqaAecHBzTeF1PTd+g/O4VpA6g3JMabE7t8Ag
MHW/wuV33HzClsHyxWotGMANaB1CaGkG0KENi0zz+IlMrCs0KmL+mslMSFfymtfk
xGSziFH/TnZAK2PJhw4eJeWeeiLLgI22Or6M92jqANqKmLGyAfM4iz6mL8c6IUUO
iFLJTnYpQNi5tMhPcf2PMPVqlZznNikZ07hxFQpi/0NFaOlS3lW/RXmHlUOuaE+p
zDAWIWpOV+wJy2ROsmAl7q7x7kPB8c+Ngzw/0Yt21Tl5CeWuP+ohpp9BAj36i92J
TcDSn42ea6XK+Sg3iv8BdiQ/2DNG44FvlSVUtnCVun2AgKHOwPsYqd48Gp2myecx
gqQ01ynIdrTmaNUJnHXm9Oqsno8fbX903YAV925+EJDuUGuA3PSAb5shExIPp8iq
rFUZY+lpDlPQDl22f1+N4wfsLNfxop0k3907Qfhxm94227kUWp83Iw5x+Qg+gytL
0A93+NYQUaWzvove6+1vOlV2eCeShHzDw4503IS0upAvodUBdjJ0rP8PE3s3lnxQ
verWg7H4/2OHsSkvvGXpTw5ajmTystAdJNr3JQdK7UiD/pK315frjWWmKI3g648/
V9geRPwWiSRa8OZgk9f1argxI2JT2ynzebeHbLDXdmgtZOgQ1O0Z/rJM9M1KnfP0
GxW4GK4OcOrasNbi8TsL4+9pcvuOSIZvhRAiF8vjwZ0/tnm1R88jXZ4+F99IsKRC
Wd6Igp6RB/cMcAXevfV5kodVrnkO0Awpf1Awsu/NpCdQTjeUjWdrgPRjH1b5Ioo+
/JqWWfrZ0fVtDQlwsSbhLrgX7LVHbr0VEriqAmfEqTOgPeVsSxUwcVBnnHx1Tid0
Qm5VdomuxGXFZIF90KT5sHlyRghWbj4yHbkxhed+WQRgwT+j3kHP3AB0qDAJq8IA
ic4aFRmyVQHjVH+gH0hCvp9iGDYz5op60CCe++1sk3NWRGB1qhzWAn0qRryTOJku
remB3QsLyDsR3YNmjOGPx1FaSAuXDSFccGrU+MAKc7q28DXHr7njcCXyggyJZW7I
TLYL+1IRsLoY0crI+rTaE7T3wsumOm95G9Jh38X2Vr+FxtNmpvLB6Y+Pcou1ixDT
76uQx3mr+F8u/JZOF7xFzZUI+6BAc+sMxv1EFcwA6lFk8g/svxjvxekY6kX3UTbT
avSn3xDdVXgdiGZM5UrzU3rUfZvaj04l8Jq3BI2jJeW8YfwzLVTv2ZSiltww7qpy
qW7TfhbDnlXv4EUw2a6KiBgHADEqqozF8sxv2yS9OcTwHET0zIwrhLgmDbtwMm/+
ghZc09yGgmE9cWbYSmq9K9SbW4fpTlMwncwAfHAEe/HxeA/sr54JC95PyvhgVbh4
hqNhyIgveP84sW8wFKVVcjMhESfvDpAQ1iqOyk3HCUgH4H4KWOy9LYDjtQfevx29
4cZCv3m5Vrc2/vS8HG+8n4xkXq9LJGX/fMOAS3XAYLkIQSw0m0O0mEAs/TqrJjMm
BIwRlqPXjNPam4OO/gtjfmoa0+K8Pxf/IYB45Xs/HAh6NyJvbvg3Q9hFzfpraNt+
0HGZyGsj8pSroZ2IKTiD/anTD1otOW1h5YGib+6z8zH1SImbcg7ClaRFGCcgka5z
eCG9HAlUe3wfJ/ILwQN37SAqmbtzCoF39ccc2cwplnTFgoS4GRc/Ws+fpznxfSZy
`protect end_protected