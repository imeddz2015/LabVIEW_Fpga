`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 16784 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/59UwEX+aE7FohaWu0/8IpTj7mav863zUNIsgIH2BWb
Abd9opeuBjbGF/waQMI2vMJTwD1ie1YueHc3nSNpEh4OXp8P5ybZFY89uyGz3ztU
W1EsuUnchJoQgbHZ/sLbgtGRgsrAFn+ZoIeGN1d6RAF2wAESJmYP8zw+p00RvjZ5
G2ATm2jrAjm+J6bPpiDE3zgrH9qdtG2uCt9Nr1qpxWVy6kQgmwbL9hDe7SzZfQdg
PdByaE8N3gt4eMh25RT1HB9UajVEWp6lompunHW5VmDFwoHLTtEqKUd0aEf2Qdft
tKw/Tow1bXwePAZH/AabJnzGZi3NtCihjO/ia+KXIvtJA7vqJLMgRS4hk1Y6lmIk
kbcBW+rPPDBGxqWxWVLKW7F98qVZiPS+n6LruDI+1kcKpJsWnqAPg5pQKpbLX4QX
953b3Xm8T+BeUuUB6zWpvTTMgV/jbqhaqI4aV6Ojh9omd8t2gjIm4BDSeinDCNTK
QC++mJY4oXaJGNbD90WJYG1AjejN/u06t5MlqFU7D7p/xnPBk38hL5njciswDtap
KmacsJY10TO8Jefud4SfuXvNIQrzm+wMZkl/dA7/06RUl4K+SX8XBV3IeU4FerXt
eL7oarD2+IruyFGztVK7/t6c3Rh/GmIUDb2341CN+wqWWRP/jucZJ9NypDZAI3U8
tx4Y4Kv1df2ga7GStBwLWARZZUYtIIxbvaccWuOeoMWut1B7qyWTq7G2HOrMuQuo
V6f9pFq03NuA5hAWnbwTvuNjsZ4u0L6iLX56aDFTWv2LE307u2nqy7oVrHZAiCKc
l043w07aevIE/mlE/UdX9a1RtKltIPJWnRqzCYp4t21NEYuyfBrzDR9lBnkYDxmI
bWv43vo2/FiyK4iAuUNI9YmZSHL07vwewBDDxQWrqUG9jcZX+xLBEH9Hh97+a9zp
hapxFo3eaDPvQjEXCILpJoEDVmN7fQXPefSRBgrEyhqo+znecKt86W+CvUmg3SbP
UmGa1kkeH07uHycfMN4T+Xh2k1acd5tl4tz4kwEhIQHoioSbN5ZIUjNItVbgst1A
EagEURao3CGSqp1AreZa0l3dPdNUgP+SyWQNRBAc9UuPMmpnjyY62K0N49gj3tGB
l88Slj3v8wAaCqlz+hsvjwqUgc0b/lWPFQvijN9weKcKul1wJmPENwGTMF435P3N
KtYME08VqDuCNKcOxXH871lilZt693APekus5+bSWCuHMUsEwrExqTJFXYbqvy6u
LyRYPUtI7K6o3J6vRrl+YRhYVAavVJ4LfEbZd8Ia/NEprzGxznqPGOKZ1lhScGp3
xxVwYD7O8wfcpvOqO9UbYnjjhgocmW0ySMyn1VQ6WnIJZz0saOlYxHRDfY9KMphH
2ZJYmQb9atKvKKr1OJ0k6HtSmpSeYSfRtonxWGESDxBes0bJYs5xOLfh7WpqxYz5
3x0eKb9ffawy7+4IaxL3rX3ume13MArKZtHnN9538D28AdPxXog3sJNGr4fzHvR/
GB5ksPxhlqqHvp5NUKh3L0B+imzc4MOmnFOYLvJeN6HNg37/hZpN4Gxi6BWkyeae
1NJGUtdxzgVuDO03+/kd523UMjxKa+wiVA4m0bpyVxbCmnP2gP4abBnCwRWeAQhJ
gsHGy6qcM3Xg0wFD2aIhBctiGVRAYkM/Folo4BD3g5UFFqtlqkZVgxuakTXpYgoa
UpZbkhX4uYOZYlpwp3DCwnlBP4bXzZnFaLO9ZnPiaBP7c1ZLwNmUlY6eSognq2Op
jBuoeE8AjNbw97/fvJ7xHQnplvwr4ph6MjDlU9TWPNGi5CzUiqUuodoU+jKi1GcH
YuypW3rq+sIHDoJzKa6mYmTfCeSHBrXxT3JBxaC8XHfxTLY+nr9zEgQ4OQoxYPrv
/HwNA7/586fMTuGEu490Mu+NoZ9HaKCqtqARDZ177u/hiJFMohdHjGT3XyoTy8Lq
j39Gde6YmSVbSqfuW76mdrt8yHrE2jDvZz+b5A0ySscX+AcKiaR/njlsJ+A6u96+
4Hw06LeWI7Ra0WtyZDbpfCZONiXf0eGQ3TlMPoeBx3+1qVC5eiO3sbT1PXCz8ONj
Y2+WzkutE02n/JFSpg4G2wuRP4OHOBue0mJGtI4PJWiNv64FuFZZ5dfP8INr0o/k
pnRiVTs5K0lilURITSLdrlqXZponm0iL8vwyqAsoWY5FW1Yi+cblb+tkXAWH7ASA
jZ5xZhGhfxvl0jF08zrPdqz10FG/MPtzXcC8WX3XFg2tU3LEk/pDJnJrdIJRoCMd
B0nfabDjtQS5h8mw3J9wZuU77aPRwr499Sgczv9UhGbs5yhjTCHCzOotFxUhiNk2
hyoaRjbj1wyjuidu9JOyylt3vHrsK3/u4naDsFvrpmP58d83f80SqvzOs/oK2p9e
FQKI5i/s3F91JW7sesPNdf17TyJeTSizDvF6xSpN6KtpY5E6OVkF4zc2XMY0ckgI
+4B/NMnNElR63WGUe26+KK1RyyzWkxpeGTNSdQVn7TiAvJXzmsO85VxXogGadpZe
8SSrfic40ihgZPQzM7ZWlN5ToHbnr/nOrI8i6xixv6f3+s4fteK7O80JYuYbT3L2
Y+2wj2INjdYhvtT1QX9ApD/Q5b5kN8heJXDWEVl/wBX7PHuFxpoaxjD0u6+Tqp1V
1aGKF4Gzil/QUvgphO/UcYToYqBzuqakPUurPASW664HmWt+GaosTT2ZBtG9esfr
c9kd4AiNBKbrJANgq9sujjT0y+7dIipStyVMQ9k1qqzWEXo/UCkcvv69IsnY+724
U1Z8MrbHp6aUC0DyFuTSeASxoHWJRM5e1kMewNI3bqS3XmcD3kJVY5hL+TkzOYd6
rzrwcU4R6amHTl3EWfw5Kojfmt8NvcR9+evD0DwMqO2ZfcwBSq9H9GmFr+yKTNo1
nIQxHCn7gkPTjmVEVP3kRTITx/Jv9QhsgN+e2qmAkkJxrgBtroyza8yo/fKy6S9N
TpYbiI8xHTi6+PX/Pel5KeVZFwjPae357A9jAUrfGy5khLqZ2qKTzXkPiX4ef7Bo
x+ZFgQN+VCDxM+8ppJQPqFo9BECRo7VqS2dDKHXvSEHLI+ESjQZ/+hIjREs2BR1R
pchCCedOp15pzixWSXDn3tAFvm58Wm/S7zwMW1dXotfULP1EwxFv4NqSo+GeMbu+
f4y8edsSoFlRKE6KMp028mamxMzudFttQAWc2Ma0y5VC2vbC3HsqY4LrsNpnpCSp
jehx7xInEyfqBEe3rW51boMedvfQcZ1cP7yCUVJWF82+TFYBKoGJ1mV8oDUAPBUu
O6h2ImuKZitFZnpiQvR5n7ys744fJ1c8PvD0gW2BhidHZ/xXOv6XT5n6JP3MAy/0
Mfr27nc/j+3jyBiTwJJ6ov5IjqGFX9ZtbSlpGxqwxSisbHYrnhj5NiDb1/x8gppy
ps4cRP0kMy/ztQS4hOSM9Mq6bG9vq4lJK5/G7WTc9RoWYesmP7HtIYvzPtVSM+F9
OeRLjf3hwRE3RxWGCdwMaTjf/kRzBstaCKFOz+54VUZua2IE587/fDUg6eE0fx4m
eKhW/oVFVF4IJq3n25fFPAH3q72+bgEymGoZgU2Yw5Y4PbWJPRKBkK/RJHFtQYyD
WtmlxyoprAnhi6tWPrIy3t8w8RMk4crRz5hi9qOnPqvtw9QH6TcJ3cTE3quO7HVG
vjQEHIfJqUFcKDLsVCrNQIJURHP4fyHvI0hI6D+yEGMQOyqFSbH6Mx3JsETYepYa
lAydl15Qb1/SqcHOL9lAi0KJMJN4qMfkQsucdtqY9fk5QCErtcHR4tn+LoxEaj1e
AvURysReutJHFCilQgKqpXvoOCE7pNnQeAAcsRQR1XWhN+7t2WQajkmDjRo+lv7V
bn17Qucj9dBCRnHapObI57ys9o36b+qgDRmu39ClSlXd3MZL4qOXE9TZRrUrtV5F
VC9R2UD1z0f/zw8PQro87gHqWFcxqiVg1TcgSKFfy36s1HVbK0zhqNHq2/urrmoP
+mW2aiAp9OJSQ8TJo/ATDwl+u8wxVSVT4Pog0AYNlvFc1YBCD7kCnLt9vwHVybMO
n2o+OzjzmS8jUXt/nxdnvkcoi/OlwRJiLs89S8J7vZoztq3QHIGXKOUGK62QOpow
qR/qcefwoJ2DYuM+9vUH6A4aSZW5lKz6ete4t0ykCZk0PijD0l+9fXE5Wxqr1Zp7
R34drOv9DMKn0QivlKIasBU1iANrErqXMGjn+N8TI7pUh65u2i4Ln1ZHL/5BdRIc
cI1MvsY1bOHG6QO1ABkUJ7I+0k3XUIuDX6aEEtzD0oDqSJe5PXebG9DkzYaVNpJ1
9PoXHyRQ8cpaztcbXlXx1c87fpyLyw2i0UD0LzlM7qXD9rkDL/tGWn6BAJ7ELU0F
IlA4hHD8adDydC3P7vz9fEyq9LOwcn407m1M2uJ3KtVMGIWVCbSbnbzTTikLcySP
ghw2qqvL0/ZZyf/joi/7rZLAzu3+w+8jNlieNY3KKSfBzIS8Lm3z3gafa4ey+Bph
k68U9Jph5fadBwluJPY8Rrce/aJl8MW8dRyUxXxyGc26/U5eqjVpR4Ed2qUZ5qka
btdCk8A7IcUcef/AbU5tX8rKPLqq40u1LsTx3zCgc2Ym+oZIOSWCIeh7yuCWsr3X
ZGDeQe5GWZWrF1n3Uszl/jPkv3WOk4N7ZqGbnisRpaUSgzA4t0ctoXchLyShHhCR
sXGND1n8GnD3+Y1uPL59vdmIVhTGprt52csAMO5N+dueYj86ZdsmYzTwxKO9mS3d
Lxu6dtulXClVLT+g1iZxiXR/kcSAjiP+bSmN7psKFkHCnxISyz1TVGF2fd0xCeEW
VeWDoWWDJIj9VhqnVhcDbpLDs/F6cFZK6WE18njC2JHWVBks1sOrmyF0VNoOVtsz
LyXivNYsSp8IlJmC+nIXJSQcLOl3nBZ/xfSamDfr4VAG06Lq1Ko3xtF51x7ZJKMX
byvf+8/fXrZoTvFsF7s0kMDCv+Rw//97OrJQRbARyK3NsQ84zpmSbIZkTyKN8pRX
XcCdaOGx22iP6i0PEmRB7WPx2AbFZhbUJO9SoA0CQQauwgEzKXVMBFkkVacyE0ka
TNmVuuJv4kmX9Y3YNidoU6rwn+CF95K+SdBcTcFnq2hD5no5XYzk98DDEHnScA6A
t6Se3755S7FQ+FII8d/+v+MMj6VOKMWmnqgXEISTThT/aBePaGs+iIZbPERlfhqp
YGTjMIq0yyjKBYfAg5P7C0w+Vw06gQZnOnIinndGPnJ9YSXyBEs46L6c4ak7yGi+
qc4PFPD7i0sm5cu2B+EqXsllO+TipaePjkA5+Z/82AYMQ28hJPMnMQbCdDHAX3Aw
4LBNRwXtAFndGPB3BjoI8APDKe4ZwHMP+nE707yi7kGJFVC1a3Krj/kSSySt0u/4
OUTumtCz+c+4yAoc2slJ25qxnvXF7ELdF78sRN/jvUP4e6cA5+AOZqcYhzzwsH+v
KWs60cZejnBUUHsUus+b7HWdi3DPcVuwwDIJ5k4TtiiC3A7zd2PsiJ9rIS0xLYoS
q2AvbhwaJcZcXCU57UUOxhBuzHn5Iy7ZlT3OpsBhvL7Rdd3rDVX0JRL9TnA2xuMQ
YAEh6W7fT0gNfE5L0FJlWCXaMffYQzh4k74nEkY+rx9MZWsRIjuIvLTR6aOArvzZ
JWiGZ4aBRowdIpX826a+XKkxURKw1/gftMY7Em0CBHtQJM2qnECvA9HS0kIFJpMZ
4/ny+j0vx5t4nEM0YeU5COVfu/Nhb2kQNDjmI5WRCGYZiMnDf1QqPd/80wj6T9y0
UOw/in7cMSbf5MqBiFgZjcQ75ZTwgQa+jXgSI2MztrgDK+F/X6dw/nscGCYr4urm
7SPQMewuvE2fm82t7y/pXkT86XiWHx7BuOOf24h+RYZ/RqTlIxZmBn5M+J3GiZse
YMiyf7Rw8zsEgrFWDUxAS3Ei6xSntIVOtT+GSrxwszbhbcXWsGdMcq72L9pIaIb/
3zuOIfgnhihX4wz7HqsGvcMVlDI9qiCrrdt9texaJiTs8pkPTDAx6C3jMAsjna38
dTkp7RbKeZf21PUAoU/a9jJCcfl9svlYiQk5MfEXDpfP4hf+FIoNKPWir1aaXbyf
NGNiwIBglC7aMO+LSDZkkTKcPJt50FhL9JVPB4voJ0UaiLMECabwW2SpMXeEAU5P
Ii41Zi41WvROykDORynsHTAaNtNIIkaucDhRKSdHfge+K/SxQlAJu87x4eW4sPBm
ibPmxUZzlnq/qeWAfI7DQWJ/DYb7zwLR9iVikRhSFdB5A40IrSXEMrKx8/j+Cixn
a0e2Zu5gCZjpd6HM/JLY6Z76Wy/ls/BeDLgn+i8ZYpnqJZ/dfUh2o6vjwHqx6/tw
yRSGPDdNKLxJViSAkdJqMt9VYpqRxeeRSDBqiv18e+d7UeI4KzvqMM85O+QdLfcl
QA38dm4tWdDekQc7QxlyK5171Ibvcgq+3CjZJHWyq9bJvzeT+H0SJSwuybL8P8ZD
41BcfRnE+gcF13NIVpXyxh2p+UFpoGTynuEB8fisqVAQeRLcrdQx4UB7lEX42+Xy
mexYG2jbkUr1RQ1K4aTyo+4d138sUz54e/y2DM18fw4n58JVlLf5vxU7x+3aMT2l
pF4dLlVwgdG988oxOmEJEi+0JKEa2PWGq0SeZiMpXBw53SorqIP6qmP5c/BjgbWU
xMfH0Zejr2f2APrFj5xe5Ai4D62+ARaxgpL7bMEgvz6wUY16Eywpq9wuRlF+g8s7
/gOVFVsBN7HqGWnkAQlbdBHG01r+5NMqSCMofpP57KWblm+k4Jqp89WHvLvdVVW0
kT74OL1ugPIngENCTK65n8GMF2p5xEdgCPU57LjGkqYtqpJ63Yu8YhFC0NuQOiDZ
bZLy5ZvgZsLgFBTyyx/I9AhtTcNT7lkvXVJ//5RGHzWX3+A3A+M7+Q1U/PZGDOuF
4WG1CE1gWlBIC7QCBBwpnfFu7oy1uC49WmvGGu5iEhFCaLpza7zPdnuWaskri6nc
eEYavaYvg3YkqvEbFIm1ybzRoWLHT2anvZR+hj5WBgHwHfFz4efmb8J6Ew1JBzcV
+Mlt9LMcIy62kPUHKHFW97GcQvH3LiGZO2AtxH+yf6Y/ofGDR2oxlVl73eCr3cO+
XHSgodtQRvDDansH2ARTYPb0oHpy9Nrk1b2EYUcMYo4d7BxJCW7pnwMRtfoYOM1/
+kzXalYoG5uYnM3bQMNFOmLUCcaig3GYu4y8PPuhdwXuWDXszKa8wrjD87apV0uL
/CxRIjY7RADNNpCkE3i4WtLaJaN84rJhdPUGpMghRGnNKGoDGr19xj9Wjz3oQJ3k
NiBX2ODHrzPXkHq7aeFxWvsFEXklWXUwEJXMcsceCZqC+tn64DIPqi4x6Ur6eDxv
VNP4em7MG8Lt/DiA0n/O62N5qP5AReiKwJsR8kpzlKkQjZ7P/43pd/D8HYGyr/VY
h7gIs62YriqFijB1R9hRQ5liU2daET+HUI9IsQD0C8HMtmaVhFlVwZ2j0SdFT7B9
6Gkp8I2yOw8edItfuCZlh+tnRHswaMz2fGkFAoCxJ1ded8NMwNmIvZcwqOnanbOv
o5LNFCj7IGTQJrRYE5PfI5cQ9JxNHG+gSx/DvVIdYs04nKFIaSqEcL/imtzbyKze
8npqrI2qzpC1rEwMrhJmC/WpBhvB2sEwKNavtNq6uCzP9CWoSgUCRmsJ3CW++XG3
SBg6oK6ejHrZDfPtwkrfhVtvDm7v+SKC8dQYGvy2HhUr9IHCnhyXJ8aS7szPSU00
byr7mklBtTImO8whZCNDXGpyj9yh3luqprcg2sha7cT5VSP5HXbP0Rv0XuBQWcUC
vgH50jo/1sRT0eIN3JUsWZhiUjO9nShyv40mV2e0zCkX/kONx0tjY9+zK063kHpi
n3jclqf1hWdZsfiupefTpCetacsuEr43yQBDDy57JRfSmArWuZ39rTYMBrE0NXVV
93FC/Kh8NRPtZJm+Qp2Uv7S3PtmRvn/uPoFykgzLl4FjrtzuZolwyg7hMIDbo/NN
TP+QM3kis5W+fJL72ifPK+YPwW23SoIFnHLjG0AGCmCbJ2Sms4rBj0l+8BFnu181
8fuQ5xqfybl52RedCLqQNQgI0tul086Ul5wGQPjZfjy/etnE7SMw2n6xA6VHTkzy
4T/uCNS8plPZvmQGzZyQkVAYy2Xu6bZ/y09HMEuLK1NZIy7CSUqMbGmAWwpfGhQE
EHl3G+a1ad6Kei9EbamV3N0cXiowqV0807PEkXzykPjb0CVfLjZg4PCMNSIxnwho
1KE+tNdgDtT5R+ed9ErKaSsxhtRbBCZAW/VsLvbIbHp71Kc9luqEcrWPSruW/jN9
2NQcXaxDg5OQHAe6ppU9BVH4nphwUpcIOfpqfIfokenh84cj6FL1X6r+V5ceSczH
bFtz7q5n3AXDleOLVHvNI+bDT5CASWebjC6omYplNYGsLqh5+5OdicJuN5D/PeUI
9Q8VdOyYDny1BMmr3DAeNQfzOU7LCR/xjcyYnXqWMmlK0lmtta5tedDqtPiER+g7
SbgK6B+hFButw0C04ahkZGll0Lzkx3r+E3JCF4mE+1SFccjilmPC5bdZ1sB/H4Mw
tCpHYLQhrTqywXKzVn7B261ec0cu7J9Yzu0qw9Mhx3CwG6RV7tD+QPHG43QysDVE
7xFk+vdnE81vX1yj6gnTu/UWDlbjkE46WHDQK1VCqQXmGmPhjX7zTSTRopbNsYQB
1BPt5Qlt3TZ7eieb3h+ZkG94FC/uyti5gVXAugB1ld882PAIlrfcy5imCGRO+Hy2
bj3jZMRbeLs3zzmWd5xhmizhiFNpBnAUaKriR1GSQ+l6WZOD6CPTsCDGKf2pvj+y
fEhcVgin7HIv4OfTA920gwCNrf+Xbq6aWYDbVsCtGqUfFaoIVjddNG+sLX8X+0aD
q5iNaXz49is2wM/nu560pxpCdiqCwfdIVG0QOlHWimTA3dVNTFyfjKPBsSqEXIDH
UtaMtoGGTKQdQ1WLNJRvOSVy4wyHgFVyz/2IrX6cmYVmcXla8lxn37OsBfH1RRot
pYGTVpSuxyI4h6YKvMtHiMeaHetz9OXp4gYi+VBxQHS8wCe139O2ghxOnJQGmtRz
uv8m2G00ol9xdzjvB9WK0hC1weHcfwNx27l2uaX2ioPrIXDD3U6KT2C2FZ6RNemn
e2OBwibp+UrZDErJUToguGqtajx3/E+FHHtCYaKkQv1GuXkO9WUZg7xwWrQlwRXl
6KPdhBh8v1xc/DGA8+h90BWEPLE0P/OnBEiCEjyh0geANYulJhHREbAWYx6TigpC
kcKb55Ic7uc0FtuUnmqm6lu3t+anqTasneesvAGyeIw3oBXtasn3U4Fh9C1VWqMf
qAAudt8lWmKlphcl7DSlNzvWOx5qCmvtrgStZ/l3zyvKFEUYkWY0ttii3ZfXBjE9
q6G12I2yhkETBBAe0gaZBSqBzOaVLga7RMFkDkxE30TNs0/BvRVOGF0nFCs0rHsB
Y9la1vq4VbrF0SVxVNxbfonGuCd6J9Zf0wEG6Kz8Lee25m7UOWneIA/sMOulXXv1
v4aFMb/gLbtZIwgoDaFMx4VbjRHr+PY9tY2vq1s7Rrox+RjQWA2TpoFGR060Yiiz
Sa77+g1HXhOCOZiY3D0Kkunu4bSWGlPM/GywNudwqsU854/M4zuZ3tXgGG/v5yp8
oF99JeBHMsccysA6hScbNcCLVz7cqGsGAa71D0hvS5zCvTkit+t7iwgmo36pWwIb
4ZoFoYuiASs5Uw0QR+6IwHUh469Ox2xrG6yKyQlvldc0GgAUWA+usKes1k0kUSu5
GiyJCKFnRnTGb5BCl24ZLfyk99FhuuosXGcRBs89V7sJoGXACHY634NcPN3PjQO8
B6VusoglN+4FdNF+JsJC4xpeurevK1K/ykxq+7K1pEY1Ibaej3PXRN5bhGu1Vsfy
QVmFsiCtd3cThh4kdTCDXs7SzrzHiOB48lSKIfkcxdukjq8J4+MIJbuOzduPhFH1
aucAgMvJvPKU2oZJ+qJXvqMJl1UstRw2HRC9ZKcMbxmDvxCFWtGx3hvMHbq8MX0Z
VJED/HCinGXPXB6rZVWaOUcZA+sUL0sDYIObLFiJRcT56hDoQvtjVEiMH7F1K5ny
+0z50mNYU71jyHPy9fxOY1wZzYGD1LKCmw/C6bD0jsueG2yU3eJW75Dfm36Z7R4/
y8egzDJf7DI/EhhexyKkp0LU03JVjUpmxgKWVQHi24L3rjWTcU2AcHqqr1bDG8wQ
m3OyOVtgsTFoR2REpCN2CVPfoXHvCXHELd7Fe1IG2mFnROHl9OT4QkAVBQ/ctir5
3EWpwG0Slp/A0yJmEb9OZkm29bT5anUei7WdjumDz3qLINdm/TXnJxZA7bymKK0e
4P6tmDcvJcGpb05bdA2JNWVyoEq/OXIRUo7Xp81TCRWEwsOIvxbMdf8VGZWL/xF2
5dFQ2TOyvRzW6+VLt+kRhI3UNnzRM+TUOgHEaJO97yGLSRySzrp7kxSmqFMPml43
6S6SQNUd+t/I5K7KedWOo19/GTBjFRVqHG94OremFZy7gCqvPsCYIiUwEuc+KnLU
ha7VPmcZpK/bl4gAsyQ/4ID/zJlCGVT9C39fw1xr7hCxW/U2X1A+qQ648pjxCqjy
EUh+/uQ2+A4zyJKgPpsIOptqHkFTS1aPtddfiEPwPwa5hS7nyqSONQuB3Bg8AJ+b
p7QILSyXMjyncDhyQBjZl3FeZRso/kSbSP6Hr6cJHj5w2+V8E1Id7qbqSA5IWG5F
Rlmd86+KDWams5y/Aoc4oomhQSFmgl/QBkA1d94FNeti36chF/+Ze2MlbvnGqIP+
qDIbKzj191g7JO9dc5xv0H4NnhbfTnyhuYBSg2ENe6Uik0Jz/l9Q9GeMqTOvVZ64
7rkMPHcC4KtUUlNWEI/LJIgRE4nj/VujPAUdHDCZzs22koje1u4zhUeCEnnk+V6U
phDgt1JTAjHmh/1P5IQx4aDqHYnb7V20HTQHb8vNureDQXPl09irdBG2Qk594UVa
OBt7OYc2JvfZQn0RnomS8BEXTaaVnk9E3rCsgG4Yjls0zwzM+t8xPx7rbKO1wXB+
Bl3+cO0BQnk5HLvJBcMM4NlNoKvjD10TYLOA9DxaR/+Gu0n2S7DQzNWJ9d7qxzuj
2I2hecvtWtpnB/UluuezuVWKqR5EwgewwM5vE3ZhbB8KqcIRqbEWDCHpf7IvVlW9
2N5bEBwHoTASos7A4IeHr5Ftmhb5xlyx6o0eAVPppC7hJUhwLDL6OgwVayrmuYlF
glvxdusI6yZRHh5ccM6WqNFVmSt4+Mhg87UXyecjD3CeBrwakFe7d0VCoqPA5bEZ
QzLwP7wRK/HdQG/FU3MKT+UkIJHJnEeo0Mg2ImgWFeA3wSlu8a/Tpn6d/jzpro3C
ZMdaoDmXM/JRN0cFXGS/BMRIRVBhJpnOeHaLfRA0aT7iIbgoEkPEZ9eVSnjXUFAX
Metn5gQngVmREK3s9jrFAWs7wlECxqwWmDQA13lG2aCDIHcEwf0uDxnIOz3IlvBf
O9SDyBURUnPzYRFHIDuYQcAWIntA9Odtk7STzeA8WTH7GfjSBjkMA2oKUJ+MLv+Z
qBDyWWo5crBaWSHAnT28NbA77ZRFOk4XVpDFohj1BdxKfT7CqVUcdQ/RUE0wzFPC
xWcdSN5RmViJpNcvXRk2yWyQMidw43nHEjKXTiXLApsBqy4argRvBzLu6zyHwsMb
M7gQnDxa6bxpT4ewZAAtMGySFzxCUoz1/tUJgS7BTsOsRu3iy28tJPh2LWMNX9/M
QwZRSbDTX7NjPAiYNLUs81LVxBv9wb1ivHdU2pL1XHrthYOQzn1aSyYtsbSkJcyc
QPezGHJbTjxRyDE2aROv4k5e7ad0dQ4gUO9uX9k21WqFc2EOMxyO8QxfvdlLtPCJ
SueKor2r/wD3zyg/vIeyYxmQqqjNEiyseGT1wMZspegG/Z6Cw9df/ytF0lazPx+K
OV1W1d3ikUv4AZMGHE1wc1Vg7V5O7Jv8RZaEGpo17OLEvTVjO+qKX5Sga4Pr9ysl
piCnFDZFGtuqZDGP5IWzZIijxwxlG+4/uYIY0O4LLfvZSL7vfeODzOa+yN2Eoq1C
h+QZx6/nyOFCHxfnmDSzdkZ4yrNQfj7hU1A+dl4zoceFOLGGymz/7KcVILt2ZV3D
DxKqqrytk01kTdLv7UQAD43rHwPlIqFXIEOmQxbtm1SFzkixLHHT5b1H6zw6SPWI
BwLodMr+qPtu6yH1JJm7BMxOlnAz7PjPtmebBwcXXnJt75+EptSJT9+P81Sg0IFT
wyo7/PXDuwztidctljs4AS5FHrvwYSrCCihcSt2QBNa2BKkyttIye+sxLMCvvyzv
a3aFXHvhTcW+co5WF7XbMCZALS/ONohOHezD79C97PoEJUWSIL403t+fVU1rKk/9
oXduPPtOz+2AJne/OsEhHqSmtO2sAcObiQj4n0evQO3BB0id+cTAlC5XpLvgjesZ
3SQ80GfsWraEK291pNyLCAotXaw5ZA8PbWzAuZGGZbN88zgEfVQ+/21bn0K6QgMb
uPXlA4EB96uBHGyF3xd9WXmVBjsOLLGWefZ5KbVUNA3JfifBtypEdAPMnZn4dyMC
vG2l6DmCd8yQ0cogBFURnw5hJf16wNB3Xz8T9H4F/rOPCYomfGCf4xCsCkoj11om
P/1BC2ZKqrjkgPjP+EFFnqnrSwDorlKw/10algpkHNcEw6crQ0qFkufc5vK8BZWZ
F51bpXwkwUtkCIZFgVDLMBq0r2G8etWADCE7EAWJCykH4b0YOaY4bHrGJqcILdlt
cHG/y1DJkwB5gWhD6gOhgg/a3h0/zRObLWLs20r1qce2lVa/0QxnT0F8APoPA0kA
DyfvWwKucEDaJQZL+h/8ra05qKafkMpkq0owVtaKciREus8NwX1FNQXC46CtCukn
yec5zqxO8FCb5aD5OgC9UdyYaMGNX1YBB33QMLP93Abc9TC5iLhaMTFBatAeBNIg
PbGMk+Z/C5y9o6Y/vDOFKWcvIslfgKvHTu+++R45vpQwSBQoZP3Vbygip6rmtAWs
dajjpGffCCAmMQ22eF+t3lvDtZhGyvWMTqC1mZPoDySrrBuRVfKkomj1o3vVXy8d
zC0c/gMBEm/NhH7Z63/owLyPnSryh4Uji7aRfdEXrooc2y0BKrrJcUNI7O+Mv3Q7
6L79HdgEjtU2C3NOPqWNMizNX+AwQr9/BQn9qy6cwduM+dQz6/t8Gdw2e1ksi4Dh
YJnR3qoZbOI4x9TojhbsvMowgUpwPKmWCRzPGymS8R3b6lIegJcpfkNxHZwiP5mH
7IdSuSaG6+sMYIuJbWqV7a17+C7ZLE5gu6MkxWqq+rYjxKh2mHyzXH0q3F1Otd3s
Myg9XBkWEQoVSTdxwi+SbIwmU2PGwuG4xf9bfN/6UmJN22at2NR2kmygyM3QgI0v
btakoDKUu56lYotjSLNrrMhgqTFhPduKb7qJRc1pm8GRf6KMvJDbTG3HBbtQPuVK
9USShjAyB7m+KHaXAol5OrN3x4jfEE5NaXSL8ZQmunYPQa8Nj2hQ8Drw2pUXK/XX
uBMrPnaHOuxtPDD07QtDz1gLwtBiKTIBSkXwvrDhIGn5CTT9Hw0FtzIU7fbDzj/A
H+9O5uVrnhmDv/LzHz6DuXxBvqVsgbe9WQgaWCGyXL3CoFhiKqwPVWC8YK/mMmkS
OuIR3xPqQo/R9cVHHn7borGCEXnlk8WFU7+LuD9AIXvHxAjToQfs8+1vLBRTl4WR
o/n3KNMIkcX5sURk8JUQ0BWgrsIpoeMsVFQ7oqycalCzqKZ8/5rZaQRjxqmsIbVZ
QOfqMrYIA5vw+9NzSvnHEWM1IQZZU3YLMEzy2Xs4sz41KSyB77mGndnXJnL2g36D
DQCrF8UMd04KS20uATlU2T+KoFkPRXaV1oc43JGelNTTzXJQCyIgaquNADf2TY/Y
Ee9XHiNgtqQL6qYHOpWhE5+jFrGrKOtU32ql/DyzIhMxGI2/Z5c3iY1Uc4+x+8nz
wwlyj/gMlqeD0f9XFpmorFbqeIYiRT1q4x0sY8nNcYR2h3rQ3/ZLVjhWk5IwCOaD
phSGWUM6/5xhr7ACp/m7/z5cvmdMc3hd//z/UQn7RxbvPjPJ/i9g2TosrSNHKjWl
t1Yhst9Q4tFkB2XaJLYTogfaXpn7UuDi/Tc57aUAwA4yopsGRFJlNHUmkg1h4tka
jY2JCupjdYCT1RhXbISphSAsQzR1RkQjq81PX5gAbO/pyUFmpkK2jFB1wvivDaBR
nHFma7dqYhsR+5IgfAVF+TyY3fyIEXUHmbRl7Qq5g6UTDkrzKRgQk6W8mM1FJf4u
OFG0ga5W3ZDf+h5Y6rBmjPE55gP14I2wfree33VWojFI0zfD0/LUAO7ILrX0Gjp1
cke2CN/VpOyLfwg/qYnRDrpgAMyEIAivkIghCRBwYU5hRcFzV/u/UcDuOGSsiSpM
FoqVW9C7ISMYf3s6hTsPRhfJUq6nWaZlaQC3igvfqZ9ZRCtTzDvox10h3rlEdO5A
jgtQdnI47YhWeiVgvmstyAeh6cbQ6MdY3FEurmvl0RiBqNOwaTRnWZZ48Qaiagtw
e5ZWfFgQElwKisdSczp+eyvGfquMEOcU5oak7OmZl3rwulC6RCvLKLD9tP1JFw4b
9dTZ+xLSLEkP+uC2mG2NFmhUt/+q55i2bNTxrViRi3JZRu0t2G9QQgO4nV+OWbfI
KSBYme9n/gf5UK3FckTk2kkCPIfH+nzP2J+yjpFwgOXCLIbsYNKwAIa196wIsBsA
znvhX9Ymz+mKt/p+QSWTvoaWTb4lZruaWWpxytyFJ5m0WUKO56RvIj6VIpsnVrjk
OSGRHDFs2O43i4z7yvqXh5Vl6CfwhWVi9TmjTbKE3o+h8xMPkeUqva4xnu0zY02G
rA05yAry0lt4yeeC8cPVbSiZtJ0UJ71CzQ3leZxrTFlI64ecJ5QeK6ISwtGYz5k+
bnjPEJjeThhq8s/amm+ANEcTbvDoLjgk27eJdVbXQT1E53Le1qta4mpITDqniuqk
aA8GM2Vmcq2Tpt3UVjHFzhPXIOnY87RtQXcLKIDNrgoI3y6wSaLR076fGg7ytXsA
xCEMpHXyPVCWHrj4Y6YVVc6rk36GrsIr02RxoFKmYAR3nNkuS7erD55X5TowfnaT
O0bhRaK6NCC/NsFNKjHjwsEGW+lWh92bxDLbRraQKnqlWPl7Zqzy2CzPhTOqnnfg
mVucZIGrKwJ5TNk5vgaLwUxru26ebqLwvD9yaXLKGfRh++vT4cRoMFGpKxZWBpfN
SIA+eX8qyNPSl/lnnRG6Og71VjzqN6AXa9ehq8ay1pjjJByYnFfJNWyU+4HbUqb3
ogfv1UJ127vN10LVo7Zx1SZH9I0TJenI1a4rsZYZc75SHqhBeMOCiIRAGoA755BC
PiRpM3CSBmH76amKwf4Tef7GR/WLIKxCyZuahg//858tK08UjCJzfeRMsve4ajB5
ighUD2P9Dbg8VOZTYyj2v6v4E/yzkH8+cZGOBkg1bjoshomyk62HwYZ+rrD2Rz1X
ntQTlZ4bqUNPIDXUvFVX6GxTFhmw+YeW9R2kArWcgpm0WCCIpu4DjEKIyP0CGLAX
x3Bstj6tjPFlOfEfOC5aMAApaOivvVJGrs4mej1rffimYbpHQBQvgoTTNOHavlis
Nt9QH/3jUp0TQhY7MR2UIEwb9Fqmv2JJVdMDvitAwrRSK+pmjnu+HyMIcVLQsk3n
nmCfXw5/kXdjqyt6EtPKp9BczA2aS0Jq9BHyBoXjErwR16x4tnQc2AzhJZrTRj8r
qTzpTtAj9mV0T3KHmMD3U3yND4JhNcHgMDy9mUHaOKTZX6u3/nhwjpPtr8jvxK+T
jZreUbixeBZ+yHKXBOAczBV38d24jm4Tj1mNpRF9AhHDNfcRgbtaG26rYeUtK9kt
Py1P8KH8EY2ZJeucc6cPaLaejpweFQe33bF6NSt1tA4CuOMXmfACxEhK08mv0X5D
+eXFMGX5xjgFkmfPpa28Jqpy+XqL5Mws8Xn8iAGGZZ03NimxdrTDUIV2kuax/x7d
6/811Teb2nqsAkfrPbMv5kE4dXZND6JvbMnDjDmdrLpDWzvZifOxIcBhDPHCZOkt
i/gUe/F8QuJM1B72Ywdj6DhHWhaNCmQtfYpUuP+/stHSXXKW4HaFSQp6l86H1RFS
IVy6CDO5cIOMHjwm6mf4d+zCxGgnxq6zWnENPgUH+qHqn/pqja3vi/DWMJt4GeJW
pvRACWxwj9vZLrUJiyqArqkAQ8P1xRsjwUyzEEC9Ky0dnHt76sVpOugTiRoOHUO9
Hsho9UA5hMg1UvZJdtpw9tTbnTUtX0+Cgjc0H5lSEBfB46woB9nqYVDW+UiQxmMm
k9DMhblqbJ/Ug5yM+pf14GXCRkMnPF8GdcMUnX2j9H/K5P9WVkfkphLCSf/ZBMEU
8ivDVO3HQHTPGlYF6aL+amiv1uaVcUJNhUOqw2oeOQrkUqeMLAJSVZngE7rHFQbn
E/UBwqju73GQawMmNjH6VFSYO+D7hhNE7/8gr4hcsTA4lXDKyp7Yu2DNwF46rOBq
l4aeqvVMFdSwUqMygjqbsoG7JqvFUQQtZm31zf8739MlMBFxu9pHotHRPOglPkQd
wwpLmk6W+SD4YSDR9DzsloGkb9WBh9uhuflFou+EqBy2yPzJiQ5mU8riVvhdOMrK
nsUeDT+B4xqRbh0+brleLZpd6PBcXnck70MjJ4oZPmWFDZQlsx4oVpS80seuaCyH
+sPbHNAvrdOOF9H2VUylI7IZPKrLF6nCgbn+xGefVY69k5Yf72NI/jD/UH8EFmag
NfY5Tdyf3FmDU7wcRLerhNOpPh+QJ0ngwrq5YqHBjZs9nyMtKdHESNjFroHvrPXP
0asv9NUhaBHeq9EoJgh3CSx6KcW220BQKoAUQ9i/VU8kV+aWFdfLGzkNn1HJ/jcW
3JWT4SY5G3+qbos1mW00/Vunpj6Pdnd/LH7ZJrm6GNAyIFU4dQ+bgYCGoGQFhTgr
EePok8Y7z7N8p88p8plOP727Zj6dfQDvWUA7WYLICdndXNw2xrIpfHIYykJNV8Cj
jOvcN666DaCXmbczkJDm+kPmYLZV4GExgjQBeavuvm+0DTJErLeMgRIiULHXRP79
joNp793GiSaPZgWKK4zxfvgQ8vxFZPWzUpxpjvuQnUv10ov6sbOVz68XFGhgcHF5
rkVixoWkTYuEED4AThGzVRrNJlV11zQugVLTodTfFkszfBuhnyiHB8qOCRjRoJEo
YVRqplXpeKC+xmk2Hi766My1zI2UQAcjAidBVNVjc6Wdc9Ft/cYO1iaiVr+E/hSU
QEWkIlluMcdHdbKNp96DzA+cpoNg5CbCjuX7y3OK32beyao13YUT/xHqxoHrhb22
7NVwCSjJmW2czV/Z7N7NKBabOWAF/iSPhKJ/y8ffMqi7an+UH6BXldmlR27rOb02
sek+uKzgy0UCJSGforg1GLVCWXA7N66JNLH1BK3b7socPFqqz8lyMkaOnXC3jPVg
bC6wo7pazMgcWUp2vAj1iAWv3ZIcoN3jkJxb81YyJex8/oKtfT06lXaZUR5z0/Kv
orHmkZ1WjQbtFZRuayF+NpEG8fcZYWcPJAc1hVFtKldXe5cw5fesOfoQzz6k/bmy
OBQxGtd22tWZmFAMeFIunXjtn7OBXAiMsZ8Q82+hHh8v37q95y9RSpYMNdKFtI1P
4tyQKOtdi1JwL3ARqLujFUa0ejlK4I8zG817exqj574WBlg8yMJ1UDDNMoTbOU3b
pLVQgwtJv0/RvbbtwPzSEayShYZpECKw8lz+l3/wsfHsRWGeSvTBQs1KyLf/7o15
g4JOcua1nvit+mlnIv/St4Ck2OOVlOwMlc+IlMsR+wYIRa/Q6fI7zBJUk3varf1G
cLicYW3/JijX/SBfU0Ymdn2GxLlwWbvCRAjcLZsUag++rJ9BKi2mE8MRdIKUzw5z
tspEzMVxxiEIFhADeyEXejnKyKKBxo/epqNQC0zauyM6dTz7phSslw8o/pN0JKRQ
Up18+3WvdvynMix8aRjGohKhjH9SESvP+A1UHnnCt/SzOswi6bndq3nm8xp4oGzB
KMZSNV/R2PbcwUBMDRmCc/1itAQXUQ1Qe/hbmbSNY1yloBU1xqaAFwnje58b5szH
wEiM8M5KWzRNQgdp9DnvVdyHwUee3kPvUibS3OIHKfiIbpx41ya5ywblN7mZDzo8
rxYSgXxr+TfBmy22QCBeMF+7xJEkohCfb/IdximynYaCRUV5tzz1h2RcNhFUIiMM
PMsF5XHmUZ0R4OnwxFRNz7bKy6afQZIqdtd/luk3PCwKspuZucS3UqHLa/3ZXvYh
Auoc+zZlaOoU4hFNlgNUJRQ8pSHvcsGXNd/CdKXBgoIKYlronwLA7srhYm3PdX14
f55eKZwH7uzzCebodEmUjGcPlrvAO+t6m6Zyk+1ECDptEwoEJm8oJC1wuozqcek7
rt+5SLw0K5L9dvNkl39ihfC6U+4BFVjPByFBK1q+AV+1B1Tkj/EHf0m94N4Ibn7h
nJm97SjyMPmwqMFpHT8TCVbqYaN3rHpS+9EBRdzFrJrECjOUbhMWF2Wr4MxsH91V
oxTTWe5LKuuMT6xLhGNyfqXKzbqVvuTHZlVeuuEZoeDU+rbtCwTouenZPTtUUK9s
wu5zxDNPwVZYLEny48WwrnG0XI4L1P5qvHCwBQdA+iiZyvRFLncSwBAmh/n4xtCX
7mXUxovp7sEDx9YuMYoRa42q85AaYFmLoNGW3IhNNQJuHB+i+dfML4pLDzPlLBp0
II6QDqmWqRGxJc+id7JvNiffsg+4oLEVnTg09ev7v00dftMJ1UAATvmC+y++nSA8
uzg2cqTh/bg6ZoD8H4vswALbfOhDv58P0j1rBIDvL5QqkmmyDXRwbKuyoLCGoaRP
OUBEWqnsKeuuQ1GYLYlVfxf15k5hmGEOpHWZqxzngn41LXADAwXbmZZJ8w5s5aiy
uUdx/dSgqTCqPCM/eRfQ2jiqBDmEPJAnwHih3Cn9UIBvDjEgCWjJ8jRo7s6KvRbC
mwA8eCtm83nHIEJvDxdhrNXomi4k7JseOFy6Xv2N5ZDfJ9M1LyhJlPwBiy5aU1bI
V7eK95DqNdGk+j+TJsfZsFfkEKmKmNxjOFTjlXNUwKxWdnPr+7nr0kPy2ZhwPf8F
J/fRyYEaBuEMNvC0C7Vq6Dz7Kuq2gv5SEfPkdV7yxv89Zlg4jBb6JcfP9uEhGBEC
MQDOsX5LPZMqKL/LCygKoVU27mOPhfCRHB5oTksL70JK6oo/dyYK5mdxpJEs37tU
3jr7OS127901SFwyjYNKTO5xa8nNrFWAOT7e/OtW3BpOb13U/bRwodhoHwyv1b5p
uPR9KagNoMGsg2iPDVpy4hmHmo9l1Ae3olT/DjyEwzPqi6N/Wwpm7tr0p2272Hhe
yh52H4ByT9EWYEPg0UwRqy6HhWNzU08CnF/5LMnhoVINbU8ClsneLsLowbOF0L7T
Qqu2Gr0koi4NBZNX8837k/uaqhyw1pPTuxjbZH6HbW/qSCbvkV1Yoqw1UJzf2pvd
2xRRP7aIewncB/RkLK24F0ei+s5HatdJ4qy0C2bp7L+YZac2Ar3OJ2AKzGmNAKJZ
XEr8W6sbjB6VMiE2MRPraVXF720Jd7U8N2PvwRP4iBW4S7XECPzo0pj3JgGhRDXp
AgOFyCTcCt2c0fmU9WbEHbUyvEDYoe9VrgMY+NEWVrojC6e8FO2H4sgl6pM3Z3qL
yr/1/uvyYPvXdcRtkFXPTYxI1eBvGE4tyNC72s6mULphKljNVW94xUuAgvsKU2GH
WhMdUYDoGAcZVhRUf2EfBbEBMzlyj9KI6RNsHVvCJt60edrGctaO99SJrc/1/He1
0G4kpvOxWfPsiMIqFK+LkUY+d8a37GNWyKlp/iVH4p5K8boP66r3lBkjH1WLeqWp
gg46PCdnCpUglqmXa0o1tOTnY7xYGUk7by0NAl5CaH1b6L8WwtLcQ7hnIFvEl6u/
nfqgHPfJ/2YfT8HOJ6HjXBUBnqvA1DfzTANfknpYUfmrlUb20kBvN1I0sYkhkFzI
wRsZtSwHYVPvBw0ij0YWfcbeRumuxKCVSvtmxa03gT4/+p3yHuG0/EJ2zwRSxEhk
AK1E93KkjqWbxl4bw2NiI1G9HhbBUE6vOoYeRejkTzeR/L/T4BMVXo/P+sp9NmnY
8AoV3jfaQrg0DrWqDj2mC8KibM0NCdCCBYHv80FruOhg8+EvwCSKnGFVFeVbHt/P
FCLNaVPEvIosPmBpuzCiYQ0E5LDxrDsHLGjAqyBhU+N8eH2hizmGGW89/Sx8YHuY
rnXlGBYFzLYp1QzyctESsPEmgPMhSjOWnEE9R2PvsjS/bpRPkfGOPA5PSpDDnStM
1OZUtnAfasNfFt7H2jtdBzkijOOnOKwTJQmFp49mjLQeFHa4TMfic7bVZ7Tm6XG4
HHwOsKC7uwUtzjfJ9H9OjBYOJwl20x+Q3b/cPdwJ7UFfW1FRdKXzfBzw7+cl85I2
tR3JptXz/PP23D7yfZlbJFdOLtkT8btWedPvX+xRbOjfAeL+l/g6a/uAWueN/ujn
H9TB93tPkn4bAA/16F1s2pkgCjnXlE/ruAJhFnY0i3nVsuVBRoQMtKt5RsAiWPV7
Sw9Of3Wqop3wNwPqtgTyv2nTJMC2Lp9FqOEZhxf2G8I5qVLps4fSTDDMAAuzNasA
2oF6WQV2cQZIcqwgNmgdxcDzA4kgss+Nrgdvi3ZWrfRIFotGGt5bQmQVXi72R66o
HLYapmgAgnsF0dadB+BrOc95uMqBDN9EHcXlbPaTchmeC+FdbIi/0CcNwP/CoI3/
iSGwaaDNQ1uxwFhBVlyBvP7KDXmecJ1hD4m4izUHWlXKwFsoSnJXLdDzJx4hs7eW
rH1pS7/ubjB04q1kZwQ1349uxCrs94fDo0E+Qn9La7v5iWP/wjd8ohMsLQhxR/Lr
cBW+eh3/+5KDpOsW7yHcacVP21/D31jfgTJWdbgRp7oZ7K+wtQuiEB5VO5NO2VFy
8R1803HGu/xMrdGRA+W8mpCDkLA4Ul3rJtU50ewd0+H4SgcPYUfZJyZK60tBaKt+
4lMRHHx5TeV1Rg9ts48W8cNOkXHsN4U/roC6RcHa13jbwiHnlzq3B84syfprR0va
M6xA3OcRCrwFabjBZs4eCDg2eOTfl5jkVwlMgPubjEKcUEv+NkXbnSwVCKZU2XJP
G+krR9+R0q3k6tm8fwyBF1AFhX3yV3z9Rplmz/U2Os+ESy9AJ2QstTj5OM0OM6jx
3YxaOHAha+PWoagTockhZ8hE55iK0kHyi03/DMTHt5lii5tOCpxLuerAt+9sFtKX
pvCFvcXkxIa3dybAsBG9Gt5+FFgCl9eRWBkd8T7tysQnr2h1q7PJPmuL8Rbn7lD6
IEc9tzxNaKb22KM9SD0A9UgI8Z/fQTptiMyb68jh5QwhDY2RGKWHzf8qup5YrmL1
ddJCKf421RTlnIKnDE9E0fNeajYZoscDLSkiufI7Y7GA0ORnZWXoPrUrbK7BPCVb
yDU+m2hXpzhoV2gzSDpLTl0tVZxp2pQViQyC71oRGiLJtD0X7aFtNiAn3bjrRDtG
4woVW6KC/B2nZC7LCeqS8pIWWzTPuQy8Zm0NBBeziWuMtzaQ4YABp6AiLfWRQXE1
VvkI+8d3/5WDDmWyRch4IHb+0+M3PDv2cuGHcmP6mghADtbPwqBf6ghrX8Bu2Rlr
IHTzaOKKnKYwSPwCqjybNRXVr6MPPPmL6ad0oHHbHK5C4AvoJTvD1TWC+pNvvOjN
U6jCWM85W0zIOxhs0IR7GPdoSIw2cYFqMJKpuq1twQz3AWqFJkl4YYQuUJdBkcem
m4mZ3e0emRE4PX40iW8JnuJTUr2hB9h3GlhMQ4YRhwr8w4j0CvBP4i6qfnugiRUv
UNMPFaBGZ5sF0cbpJfEJc1Hl3n6JgPtNuHnnIECNNH7b3Ic4qCsrGP2RTmJWMGZm
VQHwKe67BaBG7ED8cHhvsXg/sDsujqK2Ob/j18Qh2paxw36XnMunsqRwksa744qZ
2rhwG3I2HOhtKdHN13wo3EnfEsB/OsyQ2urivrcJA4TqXoH+hH2DVOMKGyYXFR5Y
gqIxnUEkQRRMrxMYr438ArO4TZuwTD93iU9zca3bZJCwehxLBoDNiLCx4T/Vrq3L
3w8rg25yobEaChCzMzcH13VmiPUFLyLZofaa0kbCwYVoJM6KOyUJQkFUqQm8WSLJ
YTtN6aKK0D2Lf6IfxyI8qN1SYZa8Y5OCFyJV4aRnkBo=
`protect end_protected