`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 10544 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/59UwEX+aE7FohaWu0/8IpTj7mav863zUNIsgIH2BWb
Abd9opeuBjbGF/waQMI2vMJTwD1ie1YueHc3nSNpEh4OXp8P5ybZFY89uyGz3ztU
W1EsuUnchJoQgbHZ/sLbgtGRgsrAFn+ZoIeGN1d6RAF2wAESJmYP8zw+p00RvjZ5
9+h/UViMu7NTQPSMcx1+4lmsWbK//vESgilpT8xz7cIzUYQuCk8fWwZ9+Yif4pGs
f1EW/N13fmEPf1GZ+tBj8zvCcD+ju7xJBDkt4A3i44RX72JFLFD+Tmoubi1OuQsd
j+QSukAdgl7xXV+TR6aKepdWF5bQp3NPoucdTC823E9/+CJ3Uda3jXZOXtj3eAb4
DnrEuOKyW84D6BF1ywhwWBX+LFoYLUazt+GHNBLuegTgLPClp3wP8KkdE72NX0wF
pisAqmheA/yhqVj4XaAHZcEQlUNF8p6THtIwf5X2oWX8p3L6gj+pjJgyOWbu3CrA
I8gRwdowAfjQO7eTFyhkp6LqUCgYcRKZ/a0cG0ujo+MPbluBSTt6R800wGVigtoF
OWhMXd8Usw78FV3VGTwgPgg4+ke+TDFXgrRhtY+2+IAA4zjsnm8FrBH80Nv9Egdm
g9W9EXDAinfhHMSZJ32I5iquOUlbadRtFRXmwe3PbVofo2eVzTywCRXkbDQJibFU
ZbMK8Swir2DLTUznq2ERi9iYbyujblemByzy7U6UOwGyeiPzGyn53chSx4BHeiZ8
m51OknPEG20UUDK5NbRoVFI0QFgBwGP8MoHufHIyN1dqOpM7zh6PGqDYiEWQAvcV
ctNKc7mz7nMSwVzIJDEcVJBgoLh2KmIawRaJSsZnwrOHGlrnfwNTc2hdxizKQv1q
3fB9YagzZnAjEzQHXTdpUEwi7M4i+awZmCLYfEfPg7/CDOIfUSGs6MzdF9d6fhWG
2CJgnrgHTwl7aL8ghthKHmKejEd8n7krrVTNE4gGz/J+Rxn9XcnJNUAffmRmDvcL
xp48paLyzThGHt/xXE1wB21Abt3D8CDLngS1WAshTmdnvUzN24qacXxLnjt7+RC2
Q5kp3a83qIGgK3MuK/Mj94ugwlw77SLe2pSyZ3Un5rSrW7zn6v1iEBIAox2h5/ND
8Gj31MAG4pdtiHekJGNskCMTxQmtFXEwI9N57BuvLlVy/pqEbFnyxNC8sRiLuqki
0v64H89RP0rktyIjrZMNpztvULV6UW6c6xqqQhJg3tUawD5Uba92EBQAVrWTx34l
gdi8R/E5KDaTn8JnwIZdcNzFGMnGSgEbk/zsWF31EEHBKTBZvybB31GDf6DOvwj9
rAVQu5PAr3A054vz9vu/bkt7PeZPH6u26794dRexgvXvdULcPlKWueDKkIoObNfA
MkmCcoVSU9pSpbkvCZZl14+EvfJYiFrv4D5ltXnkAAcSvAkBINr+iS/wLr6SmeAM
9xtk2GTep84pRfSRjQRXd5v9h5sEuwpeOoN1abX9Hd7acJ2h4H/ipdxV0cphCMTC
5ToUfAdPbzTDRv6yOYCes8GSi0QtCq/uCzohCBy7qqTa/q0RTtUyvGAjWdokTrER
pgnyjnwZZLQXVfAUlsekID5Arl9DC2Op8V2dE3l9MI5WlRtFNr83ir8AvLflWZJq
wFK3Esb7GrVvkLfQMyVqIyvBza3B8n/KDjBLrkJdqefmtpCY5Kg29BuLR6b6ISJb
LwGEsr/eqM8YKgUvvYBQu25CTBWeAOb1eKAec0oNj+rAHwp+M00H/5SfMuttb4X9
uSx158nsig1drQMzGjtwEaNaEWSA83VRxPChzdcmnTLQpNy/YE5dR5rNp9lTjaGb
Zs783R9Z+qLh2K3Pqgnw526/Y9EYie5RgjnHUt8mGJRyobF/VuiHGIiJI6Zm5ZQB
Jxwp/LwYfH7g/7tPsDEakToUgqDvMYoRbW6YvanPEeCypgXuiGu+8skIsUEU1o8c
/YwSpTFcFvjDP1Fq9GxmOgUBkfCrHXwpmah8DYrt6aCfSWdKro+fbfpbDgp20+9i
0U6eY59T7Z/sZzlYfUwiX/I8q3jLCLeJr9U+YyIupxBDzmSd0obvHWse0LZYoLJ0
+poxCcokmIlfFk1smFMtejSXA3F2UuwxioYcDm2ecJ9NZBonlsW+Bs9O2Rvgu0X9
AWDik9E+TPKW/al7rgylt3sIauyZJ6xD7MIsLXqs0FuHgyihyFcnEe7mg6XBdkpW
xOxVV+UQUJ4mQrs4JWpJawVWh+FDFhVoIBAmDWt04Pm+MC8zfOFZZObGpL25Cp8p
0KzLxhMDWnxMnHDyKHH8c8nAtQy5A1RVfksyaJ94ODlX047qcadqGeARDMHJcYqH
MwIyfjH7nZWgnolCfUZlHCuVzxaj1m72WfXP7TQ/dXLpoSSEWsKncwxsLgiAYq5k
g8AuQ7F6yApd8PxA3T6sCR9maMQiTc1GF6TZ8ns7fJaiZNMBaI5Ru0B2J+eRrX0B
IFZ4Da/Dclc4PRf2mo7pfF1wRG6+jdoZof9Txwda87bl8GimO4iujvC3S6Cf4dYC
H6oLLeo+ECSxpPsDZE9Tiqgm6prlZqpZkXMJfkmTKqyqT6AOTAvC4are4y1oRRyA
R7nJuUms5Cyh9xAyjnwvq5Au9fmM2ltl7OUQ31pqQOqfQ6A+rlF7eIws9Rila7ka
WAVjS3xbKz2apBQQLfgpAiJGnBBbx57sGngSZys7bhpuk1ixPrYgMO2mOCPdIyJN
+7UuQvU5udIg9oKBdFhJuzpx830VkOSqjeTv4QQhUqxf95s8R0mPMUFRfrO0jeGB
ZGSi3GR5ZUehAbQ2Z6uzhXz5oOfCMBvKi7CM6L+Yq9HmIftnihx96+ML2k6nyDpy
Nx33eOFLYG7gCcWFejy7hzZJB0Gz6U7LVN/UpQX1Dvq2iK6L9wyme7xY4ckv4130
R6XfKcu7svBR3ar5NMPLn7kyxtS9V+2cckyj/zxeV4qWZ2Iin4QStcSEHyDdytdQ
3aoLAcjFeJFEBp2rxguUV/tSnO4wjyWIIUbrdRMOdnpbUcrk9wxgDgXj1Wj3/8KC
rwiF+R1saEXmugfJ6lxfZJ4P/hOLLJLZYMbgKweVPBlbQL1Q81JhbwAcBZIrcc6d
9A8kWaLOwPMWhcJHqhcMUU5TKj7IKuhjj6WiwleUy5N8Hr05QLIARVzCYSw0ARp6
8F6KJNc04rD3ynKSPIbJeIAq1QZ2Smta7IxhOQqpI1mOR0aEXEKxN9QBuWXpqmAA
at0UHNw6EXxY7d43IxB6AFsLxyHc1/4YhMxBWv2JU6em1n2P/5VWK48q+nWJwMA8
DkReCf3nuPubHb0JcPM46gk4WZihW9IzOYYuHggTlOp90JrnFPs8WEjkSTYlZ5MH
swhZaRZo/96G3Ebd0I4wvzMF7igx44y129GFGCD/j5VC36S3BEn/5B3H2mk/XnvV
2p/YqWmtqzqTA6GurqoQTfXyN0La3C7z2c9HbyCPaxr8i/7U8YI3qc9XLpIwwqt+
1FWYJ4RvZhF7qY4Wmq4lifHcq11tOjsZepYzRG4S4h8LmsY4vBBAz/E6Qka4Jbtd
i0DR7MEHd5fMrYd3kfufNyGPzYoYskcWrhG348F+wFi38RTvMQIU8WAcs7XaFfVt
0/Rh4zNZFFm36/a80X5PcHJE3i8m1zBPC9w1Ezlt4XXqEdYHr9W5b2ifVN8+WFbU
iEFT4sLEC7s6dXjkQlHzYRyOUT2t8shz8ar+N3fsv8zz5or+2C/yT8+pUp7N7LsI
FFUIRNeXKwGg3O6+uqCy4Vqbi6huiiSWQbEqr04xuU3KHXJwUrktmEZ+MzFVoJxQ
Za8FCgHbf3+7y2A1zC/Tf9WP2zFx+7Qefbxfx/n9ihbPyS79sT+FKlbkaMvLJf2T
wP8QyoKQuZvXM5tw5SRB4X1DK40+v4pAckPlYAYY4Uo/JhNuV73GHebb5rn4jkKf
BLMgWKqzxGHCH0v2XFA2FMOZDs/5PYixKW3xo7jhz9qDnx/dyPzGiTHcW+IWiy5y
cqGC/XG+RxkdyrJxDE6Uin4MFIinRKu5z5iAhkr4kg+ifQmGZtPgfPEqVWekD5Hv
ZINOyKXJqjy5FugB5EpNCD6oI+hHZF5xAnBICer3OJKrhLpbzsr60F66S4kADcec
JZ6MqI8o8FfAeFH5plgZOi9Ou5mm74J1zco/WVBYgY7vlqHV4rMiW/Oc8SvWvc5E
TsEMU7e7iFNxEMmnMSJ5yMnvz13bi+fLY9FPMy5XjWaLwIKWnsMQbTc6G67MBVbZ
iEVWxkW4o9el9/YKHNybzt2nERAaVMDqpbGGHmP/njckO/fwOY4+WA4QH9zQ2A7+
hnZ+ZGvup0xn0c+pEQlInhun98+VBWx3H1mOU6b2rQ563SP+D4S2Bx3C+YchE2ks
9N8BHb3w4GSsz9wBgdJI+MOH87nL0OpbRQZ02XWpgLonTbg0xAZrlSIzgERJ984W
iQ/kOfNAYKOnuR+Gexy4HNvrykKg+nAZPsipPpNVw3dRduRbzwCV7AIzDIL0zCVX
kZm1SFJxS5PZvTO3O3fDLXM+4TlEvxdaTGTlwkw3w4t1Adzr/1r5lojoMGCJ2c4a
rx+aJgCwBDe5nSH86GMrHTDBWR2v4aS4975VYCfuLxzECcal1k1iaSTYYbUeoo4O
jAUKzmuY9V+87IqcIZB4xFUCWsdRzAYXr46toZ1tub4+Ns8odQZoaLQlLtERH1lf
aq9jf/HwiIDfnmGiE7uDaD8YijaTnDPoBqy9rFpkXc5EfeQC9rCte9Izzka08RDc
yM7M2Tho/IBP76JD1c9EdNEXhFSTxBmEOBHEnwnOM2DJ1lOaA4gKxaxb8oP9ImG1
mmI6e/Lp1Zpz+0YXnhxNyVcaUoLL3piCRPAYpGqPx0V5IVXv/Isnnvagw/NVQAQ5
HdAuXYtdjKy3tpFnGgn1xgxZZgiD4KdU45LjFy8E8SA1cYg0ggsLaTVKB3ZSPPGc
/XxRWSugd3pzUyTW+y0mPdPHOZFcV3bqS3MM3tX4FaYcC1SOovdRow7ry1EKD9AE
f7sJunbxxEfB+ZSCU1JGUtX36HpdvqBiyCAtCLvNnMfZNEGYcR4ZJsFsgP6i+Yy4
1AlPm4C6NvUppCkujWqACJFwWiAAMxTXntALGiPNgTiN3LWvKGGxMdt/eg1VHE9U
q01U/7y21Rg98sEUUsa0cmu1zZFcxsqmR0q5bKBmKA1qqBsw4CHOcZfMr0FHmyc/
W8MFBn3dBzUTfNVFXbicljxyB6Bi8ZcSGijB5+O8+B1iKyMVsTYMmNGM44M+tgRU
S/DX1T3TzL9ceodejvSKfVEwAswjRFcxwUCZXN3yuy5BZlaiWoSG9i5xic4A0KR6
OdYwBV5/xQJV4HqpZckaceetfvQuqySLk1V8x3HJfXcWzcxeZVlhDQnG6dEkR6yV
FJZDWUhpUQXDwwhP5RLJwVFMqHO5M9wAbjpWkbKzBkcYW0qzX6JLrMe9XUQqS253
lSj8MxJEytsKO6SbR9ThQySstFcycWnN75DjkIq7zmE/B9HovZ01F8ds2xzJ/PvF
KXWrCzvS+LTHHjcwxlXpltWOxnz9KEGcAOGP7qFXnvACz8pO+C7FllaYm5N90h5s
7MVmpMOk7wxUPqaM0D4zZ1BipGAhpNP+Hcasrl1B05E2i5yoSpaIUS+uYOLXWNnS
8ZzFB1Cb8OzvC7HP1RW38GPBaWxjjZ5bV8R6ZApV6fAxfqGShKnCcg1lCC/K6ard
Ij9toRqQP/wmALmKFvuOaJYE9afBjwkcMElxqcsw19PoiOPFZBa6AaZURm3mmvnI
fwHpAaum3uIAOCvWbul3uWvcBsdXikDn9Y8pLIvc/gPduZP7GvSgIV5X2UVBjLKm
F+AvWKtZSnOBnFgtOf+Tr910m/6uHtUz2+/IchTV1UJsj5oIkDlpb8zzikkQ0iZg
CSCSBDMVFr96SDsUzuKECKUqGO4evgQlUhELFFKANN7b79g1YN/5xf2MGS3FGjA1
MQ51TnEA6wjpzLbbIasCwdZclbnU0Cm9EFHYr5scbHDU83A8mSs9EBNYuxmDQIWO
ptCzaQflp4HcI4NRH6zAnkDPyHf+XRKEh8ZJ16uSUy/Behv0ui7EkiVeViEf2IWd
B+JKx4iwvJJxIp+f50ZVZWPPECdvMCLjeLm2jbaXD7BVjwG7q+EZs3xuxx7zWs2w
RRCgsmQxRcVhCbydSKkH0TtQlOPvY5WvHS+9ECHoi781NdZToOFjF8kF3Mwv/LWB
3Rl6Uh7Pd26pE2n6yDwCjalEsB3VAtdpu99VR+KKEd00448IAgOUFRWhH82sKY2X
Kp3Hci3YHcqws1sa/lXoYhW9McXFGm+zY0wU2iWxr5NEXqL2RSnvxhZZ7mccOjkm
ZAkns5kwhAFpqHPLBT2pCkJ/Lhb4DLk1pUmE96eZW4jqksmCuIt40cbVM2D5Q7Vv
ugXzbOBXmidapvl6tCChGE9d9ZlHz6ecW7JPtYMXlWO9eYW1n67w/lCYismjHq7i
bhM8wgBe1aiozq2arcp492RoqvBXAqoSTFJ/mTXyHcaq0b8g3cMY5CZEUBL9Iktt
ptJ+u07XZyXGb3ANYl9Ft3+iNEyJeUKmXfi/3HmbzNsBkTo1YDfkgcgtHHIwxcdR
cLA3wzPHXK67Jd9WC1JoO5eRlRKVncPLe+Ov9R84Dli4NfX0slnH2IJ9zRl/hj0B
re/NPw7mMfrgnzNKWtqgSRz2oS95cZaBCUYedLV8rpn+xvTcRIpwEf+ne1/vDQjY
YvyPgu1x5ib4btGxiul+GMVRazghg4yx8OBe+Z/XvU6kr1WWOQl+zruKDbayGWa8
LJzB4lBCnQb75838QAQQWxgJxkTzJSiU8BQtO+cNk5kBz1adWVkOPGvSFv5qt4q1
gDefTe/oYFfPIGbAPx3nWd13SGEsWQu/g8+KLmhV5cLscgv+a/NQIb6GG0LwZ1eE
21WIDG3VslKxr1OSqjB/aeDlq1+fG8ov+IZK8qPo9HlzEjINcYaDO2XXzmtjWDDN
PFAEeNDDafopqgw3puhe3F6J+S4+8vTqpGUgZN3rE9lWAo0uaSY30IJcSfcY8Prx
YeYeIqmlvBNAaDpHelflGKsXHQjz4ZOjS2+Vbsu5dJhSfBifMZiKkVN0AMvD5hW4
iUr34X0ftN/ZZZrQj8AuqQnSJXohQmRNGBW52fFRrJbX7zxDBKXtqp+uGt37F1GX
lVWqDdFt0nRhw+Qb8vd9XH1Y2u7Ctm9u4xdihPM3S+CzoAID/eqit0zujccT4LBt
TTN4hasHTRpYInkz7mv5Cko7P+MuUe50guO/rs9jElL7MzzYn7nVFF9ImehIGOQh
wlCRFjHPF6zPadDbs79hqo55GNxUA3NjQXaFfDsjRLkGiXahkLrXDbDGk/mi1wSs
RXSUUUjqAgeClYZeXoKHFcwhE6aVDjEgkIWKRQ+p/cVoJWihxhisKw7s0MhJO33i
1o+J9TLPHm/2XkkT4PhTbrHlyfJNGIAI3Lh4AaotU0TEtCShsa0M5eE1yqSzsROn
qcGz97WBYRUppAFaO5ZYYIa0+amzeQCRRKSoN/O73gxXamD7bZHgD2fXW1flWMYc
eMv2xPO2n7k2XnttF3+9gK1ceyZfrZFpnEJet2TDuBYdx1CYCZKhGSoabhfqmQ/E
xjCybjswAfoCqBzogCF1hD85gl9xKxe1/ZmvOdIrEORlUgGw195oZjCFz27mHHJj
S2/gdYx80MwJ/+cKEwlZ3vZblCuvI2wM7eGwsvnM6H4MiqtYwSLKXpon43QifgL8
vctuyC7S/daSm7F96B27DQFnFX33PJn28xp/msBjsUYYRioup78r753XXLzlcDrd
N6cbAxZ8QkASzbqjofS03rVV/diJ6M8JvsLjp+5fadhbomPLpXOIf1Jkqh1tncVv
JadCQnsL66ln96HpwCz0GW5Qr1gVYXCjAxLNkRUJBnS4cyPKBNofOuDeE5OwLD0Z
WwcfRdtrJb4bMZ9UPWsIBSNfql7bzvocLxcoClMiKaZD3KxUI+sfW2LFcUD954P9
bG94UCM8TVm5rPcCBU0c94zF22xx+A/GCngO+opNYaylceG9ac+272xHbEjlSXcr
x+Cqrl0fV9kPi4bL4T6RMw/6kmmwwVg5SDN9Xk8fAoh1EaHpXDRZ3qm3Gj3WX0fC
JpC0FRimb55143XwYDhexIGMkPtsh6cuWTEKkbFmMoF7Q/+k9D9rqjXTAUMYhdIc
gazkYi5TymqVVnHgrVoslm0zO2/w/0vl0u4GxoDsDdsCGDCJZ0WbK6ro1MNpdAnK
U3CuP3ZfjBAOg2rlsdteliwcEjSbsxTh4oHTeUcqe6UtT0sWL1tzViJkdTYYLtws
Lj5hRnF8Fqq0EgZFHiWQvwPTw5g9vcvXmFLHL+8vpUCdcfSiQNKtDF4qlBlApyRh
zwdjBFWbfvjkfDzhaTuGWLOI2JKktTALm/v8bsziDAVDF9fewvAy6G6A9kXNNZsN
2zNtP23Sn8Zc0Vq01NxV6l6/oQgdcNJv3j3RY+4rLRscsR95+bgvA3V67HyNyv8t
67KJjvaWjQTQR4Y9DU2HzpzyJhjS6wWT+/Sc++mLZbjygDIGcqDfVy2oxswBntXo
pbVfLlqE++fPeF4xztm9MeNkPj0djNU5zml72gs8OmDtfbLd24SX0fa0kK3qgFh6
pdl6PgOui850p97uhtElhls4E1ftJgUt4NYYS6bVerqoaUqRAV4pNoORn1DymNox
bJ9F9pvnfhpC1OEOqfW7rwXzeFTIxn5pP0UPWC0fLy1glsmLFIP+bfnG8RNh02Bz
FfwaOLnFGn9p0liGhkI4LKiRM47eaW3pg6+tqi/FfF3tMzxyLfqIy7KqofYkFzli
Pxe0OxKCzBTIxmkRRxbwgPyeTXNtQBxU6afnJ0x0jXCh0utyRdSwDbS5JfinMh0Q
ayfJXotTSREKD60g4bQGVQkpeP4aw7fPJ5PO8fPgg3aEaBShX+IaiUTerwWtorJY
xDGcynEdw7lqYWpx3GOf5/vGEW1RhLOaZXeqhv7dEvMfJ27JCmnvnq0o1n2Bn51Z
2kbdvlf/kUhzNjmB3iuWqS5C2iyZP+hrPnj9c9b2wvBp/vIPLClwkH6OFhhuTpb2
IORcKf5l9hCPH2s6Kf9ZrIb2JAooodsehVwzbPHwlmoISso9wwcMVzHFxDbzFky5
q/fczgEjjTE1mS5sXjWvpi22gYMEHmsxehULiOe8bKy4Cp099zhSPSV7TTMOsCz7
Z5tsxBNifUT1WzeXK8LfNmmgPq74tkZGSxYGIRrJ1S/spy0YG6eoTr9kaXbNxaU8
H5I8bj9F1qayDtFRZU+yxaRuZFnyQTtAgl48ZxFyZzw5wjSRl5kUAsUf2vRoeWZ5
UXA9Kc7gpHH/CnwxtLS4I6OsWqq3lk701lOeQqPeGKy3eYO/g53pPiFgs6jQbaz1
zoqZ6zobdZcPuwPhoWLHcQzYG9FOPcUrT07W7oKex6gwkXaEUCt1KaR2TEtxoQXm
K7h3cK0NMB+QYFfHbdrMOCY5P/7qzWPM67zPBTor3UC2stcvhmJ7ydos8kjooWmj
QBbVSVcCgrd5geVRN6Grq7cS/SUz/5IifXwDez5yBpMHUDtvQkU0p9EzpyAF6oF2
6ULJGJIkvnlAxohQ8T2Z98xPCKJJluvWVqR04ZA0xQabTenZWoGSlOwTD0wHqK1c
6K+SbLCIIKoUjEF5nTV/A2yG0sU2/4o50So5wdX+XEW7t1792azXscrHLFLybGPh
cRbb8XG4/ElAdQnWo1VG93NARpdpyoJG2i/gG6BhYakbgSFt/12bVEUnvD7IXJCy
eS9Rrb4aT+KmnGXcCzdKFGk2C8XTZ4sPRuf318VnyTls7zguYJF2CYUQDagUi50Y
fotNZWpcv+eMO7AzkxwcIZD/ig3c5pMk9MQzh0imxeO2lXHC2tT85SXDY4hNIN+F
m5Rj378PIWTNIkT/PdNdzm4zcwTwskyodMPsjPtAXLNh4hWWY+Ffgk1DvjxFj/k/
PjhHzOpb48GWdP9KcE7HUgLNa6PFBK8hjKZAwmISeGOzuvDV5CN8uKevh1MnbvyB
R9rcF+vILBIci8wM64h/uRj7NVrYUWsq7m67dneCJTx1LrMBJIVlTbZIVjW8/KT/
FV3GiJguRTSUbqIU0wf8o4TfO4MU5n8oWbCYE526oAs9LSsc4RUDK1chGKwIUTge
mbnddEbp44viO9AtPipg3lRS7HMklC7pBmKS/KeFjZmxyZkPQA6OWxnn2Zv48yc0
Unun6ZFsoWYm85AENaU+F11pN5pWr+mt/tfu8vayWf4SM6B6MzlJSwpFdV85ZofZ
cKj7uAQjrjb1CMfKgnLad8VaoKe1l3QPDD+0WfeJDYLJRZk5D4snD1H4ds/GerGl
eBtnCeWTSmkMsSCVg4GpmULIXNjQtk6UNCxKQLsmp83oBvWu9yKtdDJ8YiDfidq9
0TakFDjNG1RsP9cpNMde4DQsALxjeFbPt410QH6XjicXX/ANl8wPuY8J5qavKsOj
SJU49LePQO/2shLv4l3VDcDMaihvYqPtWxw7RHc9pdOAk6H9glyZzrQfwXWcG4wH
bOYVcybjPIBg9UPh/2kJPrQB9GIoQR+5hrQxa6Fe5uU/dIerHNJmkoob9urmrHwX
boWGh/g59jxf7eG+h8CBHe3LYFOcrUoUzhZgezEGdZ45XHYIs7BZ97EXtbubRqKN
+P8oebd2W370m5R0T6DwPArZm4N+DXWmeZnaZxxShAqzo9qAua3RLXXjfjuhZOrL
Hcd9vt8g6ONTgTHKMfdB58xhlcaVKM9z9wgKfNJ5n5ycSZWOa4EHek+h8GYRiaIN
Ut6woMJYVyjyiXBanvqZUi132ZPOSbLWhJeGKLMB0V7EYDIgwV2Hxg+Ye5WYO2vY
Bu1SoKHvS29rZoOO2bWgDv5a5sWHgXReC8BpEvMKeiCHe9Dglsyi1KMceFGR371K
ByTrVi76lGh6U/SxV93ibmcf0LhfVrrJw7B1vTTgOG1kW2OgI0tHVseEQW7vxy5B
p0MVf8a82tu+OZkSUxEYtel1hsA6dnkrdk52paLih0eOMU0Wsjd9Z5C6W02BoBeq
Pph0xf4Mt6x3pDV1NvgN18L+kpKbMcimCCAdf//y4Cb8LEJ1CUP3uYBjgzCp394W
aSkGlOb+/tPhEbYKENhSMvet/kXqTckXkwN3I15Qf56fZDxsPwuaNFeq0T+8AWwk
o+hUvY3jmT2jW1Fkqyk5WJPKcQwWMvy8BMMs/j/8tYM0hEURgepsjLzstI1mNYGB
aHHUucs65Pnwi3LM+g5ykyMhnm63mm7Nd1+wsPbURPdrX8m3lppO1A5sWs5tayPU
Ao6Cuv/bwKiLlOOj8So7jJT9mTDzCXmVtoiQXeYI/yZ9ii7btq5vFht4OUB1GMja
aXGQpyqrLzmgM1s1OH38Sj+0pGmwj5tEtzX78nP1Ci5QmGXNFi1O0MYbTa1ykT5X
PzfsF8c6vSewWvwohbstBYp9C+1DyN7CRUlftIf4j8g3/jDWcrly180gi+lDeLTC
Rgh2rFyGy6z8U5wK0Ynn/P8HUp2G0vMbjgcjFJXUwJ8SqKFaXC9acc+Qp/2+/LPQ
/OuxNIj2PXohsP+YiGnTqt3CnwMT9FWAG3O/9cdD6PFc8wqoTWFPisSyuFC3Y3BS
a970tJS3YgzzE8Hu8Bo8PFIzfpaMHgXgQHb2qHjdapAJOXwUWQ3KxLJZx+grNhWV
8PgT/TrSS8HyYuT8w8fr7Vjp+VVZvBm7XkL5DRusmm03pwuYlyDuVF0z6Yy8W+fa
9z0TQ4ZTQa8PtSY82gbYeV7Pj8Z63Bru+/daok14ioYssTHmlIEBldCD1QCtUZ91
KgJYhR808zzYzBRwrnDJs/oP1dOd41fxuQxKmRXJN2USw/l2VH78O7HIVD5uHMtC
W3+zuiZLf+SOgJF7nN8opDB3h2XeMpsTu+3sx1RBcIPGqq+vP23TD2+GCMAL3+N8
LNHoAyjOICCJAqIIm2xn6+JTWJ5QCqdZNTFZZbwEuyBG+5mfFLPOaGy9uzgtBR4a
L/8bxVMb3isZqAKe47T4Bw5DvyI9bc/gZw427s5uJ2LX3afHrgYCwKDDqgcGdz/g
X/o7D0sG7/aW+DNevmPPNfcD/OVXnE1Qj4cTahwdC0GuziYaYzoLDPubtwUc5tt9
tv1SvCqtS3rKp7wQisjTaLmU0sGNtp0qkqXDKcmXVkTrfwoRB8R2PjwHIGjz5S8a
E3T+xLsUekpgEkH9OUpYHsfidOIpCn1lsPtYEJ7VGupceWXNHgghfMXYzR/Tqs1k
fJGmcCA02wTMXdk6cvibNZFjRetIsyZnhSOeauKbHgRSswyzEjKMJHf9OS2MZaHH
zs3ChmFDZ+4w8C4TGFS1YegxuI8WDZqQaRWw91Y1zeV/wcoJzJxBgcvfGvya7usd
tMV9OuwJM2fnkVnsCvAY763diIkRFD3lNFbaDdp8pZr84cSqTXj17QcFPkHP0iF6
3wQQjE7nTmCWoj+NB6yHKcP57ofgRiLTrqDeuweQxlzW2B68MGu3+L27c+2DdpTv
QEm/HcLLwp4ZyZGaKwLcfslPv7PHLXnnHgNhLt0TObq3i5AhE4qwC2VJ3kgCXdt/
UizYPpQnBTAAXi263mZfK3qAWob7NPHX2PyweHzzMLgyX5JHOBdzYB+7JyaauSDK
fro5vHdIqt85lultazBvDj39hh0sQzR6tOGhZS4lqMrbepXAp3MUqiDTZZ3in7LM
ZsQiUfcUi4f8lx3+ewgSvvojVc67iIBdUTovU8GYFTHyOPB3NOXuWLshQ/DLcSj8
bnKtcpa4HLhpr5hVOG0xEvpCab5zo35uz6ZJ20x4jnJ6J/Tg0/afKJ3hb2CyvQ1J
jQqubQYxBqEXXnEmq1Jvuj7jXKnnwaE2/kSWUvhADSliC5l85qPnYdzkgNT0awaR
3suGhP7OuFkWY1zgUDsKbkxZ/cCZXL4F0sPUAkN4ijOehYHV4jGsP+QeNOoR3/eY
YtzyBaeFhcLrIE/3HMBTVCOVfs3hU+Hn8L0Kbtaz7FxNV6ahH7rowjEBGhCAacGe
4ZilH68FUa+3Xji3EJA9eBhuGyXDNCHJEscM8TzHtcrC0f/GwJMD6kxD9y9r5Myi
ME0Anoa2Rl5BUUShlqjEHgh9ujGYkBkBa75I1QVH26cMeCsP6rKd11h6XHjGt/Cl
+t0a9ePuJNXdrHBndR1fFvswMYHdphSR8K91DqyYAXM9mhRHOgs4qWgbXdOXySyo
yFuIGfijRqutV5yDYpdXDrGKwS7CM23ATwzvNxtSToANTDoHmpn2jmO/rbsx7niz
JA8A7tvRJyVq+fi3EQaKQf+4VtnJJ00QleYLfOAJzA9ElAPlRhwJOX92a9tPpoQJ
G64VQ34C0+awKttc6HDKs8lkCRctOPRLkwVWpb3msAx1T3VGDdna5Am2x9uBm/Gd
4fgYNcqRihgLwFE08uOr5GKnyfcymBDDP2tIzyE3nbnXN4zITM4zmVSCXSi3L01s
QJeUNHM68ZQfpsknwbsz21wgm5m7ggDAeA6kR/XaA/YnqAZxcp4dIKFueKlx80n1
tXR+nSPiD8coMIZrKAF5Tp6lR3etU/LdEef/1Fd0dbmExR3Jdiq8VE4ZoCQItEgA
2aRPSFjFWLE1dVaGi6NaPIfgahLq+ryVOeEHwoE1+DRctacTS060CzNm/YOUB6WK
hOZcrap6+DMb7d+UJ/5JC9VOcM26YmVwjEi5PeRls706cg7nLa3rzQX6Q0e2T9Dl
VHQ6/iXgHTFIcdLTBSDGVUZyUGcb5A7D5L2jEWoOIAzsUrcm0lPF+9B3rBwFec1W
JE3TmDb632zT31r7Pqp3a9Y2QeeeRuGxqEy52jFKOOSpdtI5gn4ANHEFKCkTe+H8
VqoYOEQl6HarhrH3yPz41shT2T/IxbeSF2QdscunxScf3/Axy4eSdvX0g9M86Kob
uK9VWk1EQpbtJ5lSLuVZe1VFomJoevo+FaBL0gETf0M=
`protect end_protected