`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 2832 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/9huKRhRMtvnNqb3Z+UU7TahEoHV+T8U3P3ufru7l1O
3DlgtZzb9QxCbOjthp9+wDkjygH0eUfDrEl1ovhZG63fJH+b6iIa2eefku56VIua
W92V3G83KPEXU450BlIYNEFepOQ44WMoMppCJZi6bot8OKCjr4YRsbhQQIyaOmtz
1HnMeXBfvmyZgjqpQsw0WROxUWhICwP4j9fmG4FUqGvqFKJeK8xBn1U6GqIQpGTM
jLIbmjtrH2WTE4xaiIRqVbmhjk6Cu+5W2utlidi0P+zPoLPWLNshll/KOnIveq+7
eDcZecEmDELJod4+FFGrEJCWkLwFvl0bAxtUEEFSaukfeITC4wu6NQIzfvLHiBRo
7bZfq5eU3FkG0qlcBQq4Be+uUxt9TXOxM0tudiKcPGIsmQiOtazUz1tXzGzBD8UF
QdgAmRjVSUUbCN8Oou5cYjzwNJQeLvEdB6fPo+yueUozEmp1IwxG4pbJC6OtSDND
QHfSzQppeyxIF6+aNqzC7eAM+c7sVG/5i/TgWrBL9Rj9q41Q3aLbnpd/Dg/2owQe
j0Y9ftTPeGj8OD/kMFhgym7PGVAi1GwpIAzhdhQ+AjiymYL7OfIx7uQE0xiwH39E
AOyY+m5r/Vb3jt8KG0Pfn50ey5ksTnesnyFmK3vawZ09yHEQn+bZu4oF9PaFrsry
azDYhVEX9csu8hKEvaVeCEOH1cHN5XOzpc2HT0i4fmuRppZo4DyibzgkAeNdsYLY
aKr/jYoweehWmMLT/0F9MLQD9XFu04ytyg8ZtmFOvD1mD7J1+qGrNByqynmpYJO4
FxAuay+iaU4aRbiuo3QKB0oLv83q044ZonPF0WH35WMvoeA04CnQpzX9ggaKHM8f
VffEk0EQI+XvhUYL7jyevAuZokckLtphK8zPlOhmWcQ12fZA9mab6fxneNUTYZVJ
T933UwVcUV96RiwzfoDUfu2/YKB81MXG5K3YnaxYbKK6lwb1GX7hkbtYDY9K8Ox3
zOHO8rjPHU0f1GZqMPTTNRj/lJ2argOrIZ1xiOeupZXdpNb7AtjTk0RsAHpf+G9U
4c4xrLuELP7l23ZC6FBbm1PDeKRaMttSYKdR4uwVb9vRTYMgcqmLUrr6/x8f+cNK
hjToEQsROSKDf+f5IO2USJ4rGg12rbdRsEfxOB+j/joG8/vGfX8bOneBgg+p5NTW
0TFav2nNkvuTItEauYK269ghb1VHDDnFnJ+5WuqZ9WXSmvACy1Wl6Qg+SkShtOrh
rc+C7v2GvHH7hlahE3IpMJBjCVjfB/dTA2gT5tHykp8EbicyjxUAjyKJoOjr2IG2
t6XS6vulyKW00uWDdoph57uCq1GMgVkJ2slQU1dOq7AnxMOwLt6KHnxkkZbYoI/q
udgLGYm8gtDyv7uNPvn+d+NTvQRgiIwbUKseHU4Dud/zTvXgqyaX1s+OeVt4OOWK
0JxoNUsO9DjoTybmtNxs678PcIkEOKFYw1fu3xQy1Xzu5kEfCFnQA6ZwYhpjCOgW
KdSCZyGsU14GWbYiLYHfNwiFuO17sBLHW6qxzWiUVNTqMePqUdLfZ1RkJVYLMMRt
6BsoUgol0Np4uq8vLhNex2dn1Irg0VmmpKLbeaj+ePy/84wOoEPfGEqDFzT2AQer
Z8O8tFMFOn4abIxA8hr5pDNdAu7Y5v7vDlxV1c3NYcCLbkZtNfGQZE0QXyw+bikl
pNf2sJXP5PSV356ecwp6DIOMxSlNf5MhlRqzTXk9RsSiySRlM2TDPmnH/Rbgsy0N
W66c98/j8liim/HgAL2lrMBUSOXyHA/BLG2VdeqHRg+/28r7vjjeWhKLXJ096uly
WLWszzA9fpeNTxMTXKumTTsknrQ1E8rhhPeL9xemN9KLxz0wRFaik2qAz5I/W53d
8kmG8/OR6art0rJ6udSdxKSKBjFQEI0N4puvsDUwyec0xxN+BzespiUFq1GRjtFC
ItfofeJFTj2rFaGnTEdkMo529E+hu0ZM2CpDVAIkv5l5KonWRukLrjb5pFp5AXOP
pxs4UPN+G4lNANpCQfCItjFaTlfDJxQJ3Qa/EMCiYewsTm4/jeDSfHCdB68LF8zE
dOhy9JY4TcWd3O5IVxNIcs8HR9KhMIe/KC8HUXs2drVVIkkfsOQ6YJptJSCK4QvX
Q+lwD4YkyKIVayJJxVt8wBJFUcpN8dMIntPSRlyXCDepkPpxQ8fpYvAuBcEj8Thd
Bzjgur86eOJIUOd10V6QZ2tMVCQozWzTUKipG0x/8WUsvMzUr1v/thdW1dZRkZQe
ws3tgn0gzJUhstb0VPgx5+Ou5jy26fLH4h2qOOiT9s/pWQbUQVPBGBvdNZ8wRAqP
lQZvry/VpznoBvNNZFeag3KuZO7MeRBfoFT/XfhQfk7q1YhXqeDrY2NK3WnQS/XO
LBT6+9iFsynKdYwZKYat+M+6wx4aqNFG30SLHzimrns3/YxzKL6+XeHiHRfdJKvB
vAnVQin695sCoEC2k8cV+ew16vWNGl9SXZTlFyDfCAudEH6nvJ+N5jhntZHZ7bJi
YQqeJDJhKKe9yReMgv96xF25Ir9eDruW0cBTKdBBe+NT/CJriWYsx8613paOw+T7
m7ISUytID5RSoFF6usFtGZ8yOxCO39yATnOaCLh0MyziiFX0ABFrNTh9jU3K9vd0
2Ug4pNYnaD6gojX2krnk2VhOt0lpYSVBV0tqiDPbz2676KQ48Wf7Th5IyK8ptC0w
7Z3o8zJ3cIMxDOrPqfTbqlgtpGhZR/K8w4s6CBY04y7EgHDATtY+DlF0yFzyI3DM
80JpOxURGoaz3qhFKdKf2DpF8JF/NWvvuj+zl8JSaBeywZJ1PPNMwJLKrdiCdbBa
f4gZIG+Sp6BizKJIWS8Sc7aCKP5piFNNKBiFo9VJbVep6LwbAO79/7Zv872TEIHQ
sSTeMiYI1/RUi3DdUjf7e+WEywz84e3BRKs0g4MqmWOGtt4CA40Ij7rbMLmh4aTv
BQ8+b7CDnRTg53tYjapfYwt6TaoX17FtwXI6NExNYt6Qx3fqqQchexL/+5OBYOcs
GCyy+9l/ZUtqclxMyMi1ccejK2MN4VbqrzBaC+wPKytnAReL3JpFZOph2BjIe9Q5
zZEp4GqyDJtF1vBhumpS1eUoXll+avyQvpIuh+HrG16le6yUO7L8ymszYXMtSWU8
zmwwh2Spnx1hW875RKSscgssiq5F8KgtyIE+xhBigXWzOD0o6bAAQQ8cIu2+pZoq
c9IGo7/tip8O9V9K9LXwQzlyixa6vPwG+wT7VobUqdFmYe2pKgejMZJ12O2plyuq
zmQ9yQhkP6+aJNx6SYVXKchx9un3rlyJ1ysbnELxl4bvYUPycPp1ZUGLqu3LTeOI
XO2uGQDkB5nhNt6BSwaQghLyQdfcZrxXgkuouEZIgHG6pnkWxiEzojlZ3Ncz6/S+
ZeVSzjNy04QwltDNBnUIr6mX8Zdc3z+d28IXWynHzpewYBJMlRgbmGFQtvZ/QVGB
eX34PsQZ6QoyyNRhMeIN/A+zZZOtb8a1Fe90wZEeTE08ReY6M/0QUjnFo5tQG1Uo
1bDR6XDsRrLQfBiWiru6LGA2PF+U7G6SjpLADOj4VxT5cxv2svOG5PYORZIugJqb
ytu/QaC9fZtIu/vSwhmqAaGDrECiVmMNfgwXMfe8EbnQyQ/gP/uwnVkSkPX1bWcr
UdFmfzM0U6I7mpJyagN58u0ehZ3kVzCCR8ojH11+slW9bVhsR2GsWog+zRKDghbL
`protect end_protected