`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 5408 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/9huKRhRMtvnNqb3Z+UU7TahEoHV+T8U3P3ufru7l1O
3DlgtZzb9QxCbOjthp9+wDkjygH0eUfDrEl1ovhZG62BUgtYl/tdbgM6dq++Bvzt
If44Y4BW7I4BL5ablkFirB3CpF8af/dV2Er/HUFcB/c7ksgkcyaeAI32rvbARD++
DuUdYW+5KGFV0WcvtPnC5ihjuEm+X1q0BFcp19Xv17Aijqxqq2sX2bKBJ1hnwvuy
U99NGowD4NiJtCQKb6v+ZqmXvVWL89PLfn5VyEl+dqrNtG2p08UfK7gCZqU4985h
OCsev/aG2vF0cl3ZBijyDBNYu7ITSfjGRegMd3Q8MkAkAbxUkGLSFK39cF1GPf6q
2xg9DwhvG/OccHLtAdhhA3F5cH/SJPJv+9tuYFxSJHx9lNQGpjasLxh7xfhp9lGb
lQ8B9S6wAOz2ubIClCQ3+XRkBzyzcNip35RXn9Kf6w6sSA0XMSXOe/3kFQgZwJZX
Mp/2hkSCgxN7qtKJym9D5dX7xwuWbJ/N1cvplmExGY/0JEIuHvA8mWAlhQWW5haX
FHvBYZRsp+mH3gNljYv+xmdbkzdBDtXLpQLZDCT1VBv01QtJCjPY7AxCukEX+0UE
FQj6BdpSzr4dyv6mutNw85Vp/zpA8X3lemLR3ecAK5trA5SG1WEhnRERyDvG1Uo5
cPeBDakeAiGm+IKd3StmH8PU8QwG/0rEOCwDO/1a2lVU1H/Z7BRtnMms4wxYYrzo
nBpJDjVL/FyXja1Q79UeyHZRmJS9f3kQlnIPfRRi9Br/xNFG/VJqa6Yat4N0bxrB
4RstpuRL770No9JB5BC9Sizid0jo6TNVal6LqRhtGTA7V4AK+ecwm/2kdy5XhEhs
YGicmKq6yJ08WjJalJGCQMxEUwlv1PmVWPJj+/papCxfpdHzj7B2H+gEE5iP8hAC
q9DjkbwFDdkiqjKCdLFp4H+gozhHFh8pnSNA4v0cmzEqgtZXmbc5eI4x/LhyWHX+
ETsoQf4puuMjTsUZuAz92Z8ciMmJCntWwNWBkCvwqHeEI0k7gV76Ft1c2AexOnBJ
KVC7I363xVAtv6GMTXr+ojCA+bkrs8veWGJ1rcQi6cGasc1Cjnbdnz4psGNrKKpz
cwboB3YDbfa2IYXxzSENHor0P3SLzSUimgnH15cwRSc/cvk2D1qe92Aj70mjRhqL
M46TeHfqWSM9hZekLvA9P61Lg5ShKtG90ldjvjLjdVTrzMwpM/MYY7sM49EkTjaY
40eDpkJC9uZ8zG6gDYC2/NsXnVHY0SrwtfqzPHn6MiG27OSiSS9NSEPxcNsgZ5b1
LSJ26EGNzGIzEYPhtakztc4jZKFwv5MIPkWyMUzLVFry4Mi4aDYx2Tvcos8ywQEr
cEtHcx2bciMG4ahulrulwuh0HFg/snHAs8mWAzFzTCDYg4GU+TNOphQ3bhFjIxV9
d6SMoRCAUU1J5ACCs3bat6BCUeLl2DrUsWQtRk2InNNzWzmngMKWIa7r8LMQ1KCp
kdnzkpvjd470VjEPaUhUngglUspDNTXC1tBxYXWASdgYksCYvul/rQCoROSKq27M
SNkvNosoaaQe/zogAS0FjEloCHleU5+9HqQ3qfbMbANrCZgFOc1M63YswuvYdhnI
qCfwLXE0OEx8Vyr1jzL2ifV09YOPoHD4ysDOhdF7cqI8PSkaa3Ae2w0MrJrJ7+IT
agf66bk1gziBywlooVoFc/EbyBSae4qo1inCZ34pIHzlA8Z8tPnWtr+amLYv6PCj
Yqsfy8TXxYmy8L0fH/w2GwKp4UlVPfkwOih5N/fwNZQLbns8UwG2xW1HzFlu7Ob3
jzYMx0nwPVnnhd72VCTGK13ui8QifSC3hQaJJutvM6cuTZpO8mhqJuJTmrRjk/ET
eKeRw0eqtHgWR7JmlYb0mX1MWQ4F5mg013KyJsz7vl5m9xHEpBY6IqW+766r+HRM
L+3AtA7i069Q7bA+UB1Y7YP8xUVog8+Qc4myp5Fs8XEhfsZE3VUcvyaOKk5Avak1
craYbcrvzOecEwemdKLC5z1cvx+YVMrffDreM2h49XQWF8v01DT2FRBNEUwx9HBn
j79pJykElFSJDz4tVSAl0BjShykTr2I9kCQ3YiwZY7IoaGyvTTAhCz0ugzCbRr8q
LhmMfvDdqUF2P08BxcI773WewG3iCQ5PEqs3QFdxTC65EyHhVeJfpx2CEL5Xch9S
ovY6jAmeDaMz7L+cWQxylaUc0tsgbXxjZcQR5IsoHqAL1Z63CP0zkRLCTMGiZyau
5rPg3VzLCCkkycTWrV4MBkzDW6xVXzZ7JKuN5zFZPx052JOWZeqwN/eKMbMa9Vuv
LDwMjL23IJLNHUuuKK/E4nNFZBn3GCipLlkMKPb2wMrRLA9amNAWC8gQ0+uOEUwU
B1+a2Zj30qN/VRxyK0fJg6bgRmHhvo6EbI9yrSNBxWJH19Fbbfo84ynM9BBkwKaf
Tz9Yin3wdeqWTnieae+WrB/KHeBRnbl2kMkIEBgQyCRiLQjgKAdDx1hHnSXmE8QR
dIi+OC+i/ZTFllZvIFomFO1GPoZnJ1HfH0DmGl/YB1PBIz/OHyCxP7OfdJNuUhTI
bZKG43zn5tNuWRbGrIMHgP5HQeLEv0yFyfQSbu+nxHKj+OhaUZJosxzmaUuHDhRj
/mWESdCD3DroReK8WBD5DrIoEtSQ3/C6sQnWybNtx7IN7mrX6xUj2dxVK6OBw1/Q
4YxxNtcnk/X+UnR1OXXpJQ1jFWDBmN1yWteGmfS//lL23fSHHsWb/VRb7PcQbhDC
HayDRNOjYyBzvXX4koTOUNeqxDsBVU/vqZWlwAEx0GVN+4TZ+JWmId/gM2eN3zEI
QmaZdiC+YqPAhbeFm/Sqi5H5n6gcDU3xzm18h2b2+MBuc+2pwizxoJ39yEWR2Gqr
wDhu9Rn29yrhIFefkwhP1hamKmtSQo7hPFjtPLavK8WldPaX9c1+zK5P2Wi5gONT
DDJ10tGKNwth92ruEy65dyzTgUKKrLcILiLQ2qmSW0v4SFTF6AzHu2nXC/M0W19J
+pZhpzN4NLEHCT6874VzzG9si7RtfyNrhvESP+FTQ52OsMWgXgCAiOK5MLpJ+J1A
DCJSKs7D3sWtzBgwu+NXHWf8QnrAJgryrY4ubzfxe16haKfKLgt3lYCWW1zoLwkp
WNkEsDJcGXQ3qHzZn8GcgeEjnQ71qiIuQuCsRbKBMqZjpbqRjsf0D1gdyAU7RJ0R
7o+I+W+eUGONKEOMc9VmJoMe/apHM6+/8+kHzU1iccCkuMr4FoJxRU8kfVTl67/E
+HYBXohXUiYTAuxnMG80DTP83CjErRS7wLimW1G/UidxhP5S+eju07MCNyWkw8NI
6F3hqI/NDyKNsuOESWrz+LVjE45Ksgpgw2gaLn8x4h7QeNHeNr906EDMhBTalrDA
ITQAbfUJPrEyBHbop5feH0yF0NYmTddPxo1V0PDHgn8uomXpQsd/4HvtNS9oqzPH
YO93OhoAKiipFsEIcnO2bJFrfNKT5FsAgGPIB1LCK9tEGQsf9btbdBt0NTpF9bSW
+yrtPr7UVriMf2gdX2hnhOrNP1KXAewtZS6Lopg8xx5pPo+oANPy+ONT6Bvx8BnO
sKWcu+J92BRw2Zd/V/dC6UAvAkUbsrQrdLd0EKMR/JAQLqHmPMrL8Zjs+0zACRyc
6o4pm+FFH+zfR9psBtFmJr69ZgUCLp8rTNwtYbCgy5jG7X/gMzC/T3CKEz64znKr
GOS7FyTW+6EAjY1acCwrqxWbuyCu0H7xZX4blLyy9mmFUvQ8Y2Hvs+UudAFz2UHC
5KwSDoyF1Xa/i6os2U6GKZ//wBh4QULES5xiPNFk/PlbF5zGWsJm43UaZ/N4kdQA
Uir+DfJqsw0it1x7ju327jq2pY5RE2P2gvvtHosmNdFRS/7A0aNW2tespMyTgIs0
79HJU5OhbyGKyRoxuEO7OP4Oifwim82Fpavib4CupeXSpnByaqYN8gZyR4+veWIe
09sKwh2cXe2Ku7h+S7VzfyUwZUWF/3eYv97eT2cfLPCrZ1LyNbxpdX2LrMvBL+HM
nC1WRqwRP5cPlB9g5ODiQkBjZ4ovb/UEofw1333gs8OxuYtDODemUAbr1YoVrxIl
jwcH+5nCvQ0MhsNuFapVnPN6lE2eEpBjiLHNpDVJsomsc6kiJDEPiIuyFIm0oCgM
MYXCsLzWVnuLM8RU2sck3wnm2ZMMKoTW0xp2MMy4Cxx65keD8hdg7MgHXiKiZUJA
RerHqPjYU1tqechqCcKA5nT2Y3Tp1zGnB+yhjMn3FKV3YN4De0EptzQW9WDJkhjN
euhj72z6Co3xK6KhFWIYf1MiUH0t6zF5GTbLvmX+NPGxXyhkGAR7mgih+bRNEpF8
NMF72B71ESYZ/T/kCfLpljrTzrbBCAZTnWMh7hBLc5kdU/TuQ3Mkb83g2fXcorIc
4QKMbyoFTruwSPAcwh0mFvawI6VdjoSSy9BML+eI4rSpkNnsd4b3IfE1SZgGQv8D
GNiIqoCy89BbQhY+k051dTKsb6hL7e1ocY/3XVOCQN5PvdGk0/oTxLNxbNsNvmHd
jvdSSa72kK58Qe1FK7w7TCkB7jdeSLtbVt7MyGIRdQBINR/sy3Om60PzFUViveg3
aa8TmikOBXSOTx/wpogkvJ0Q2KMe8PyXWcmOrFL0y0G6GZ2ywppNUd24tY0qRlaA
4BAu0E28LGevn/osytCiW6dph8vkhU5zvdAvc+AH3g6sOoNVDn908XCY3bMXtNjq
GFVUvXFQLomGCO1Ec7jTW0rHrMoOF5HR0VCxV3CrrM1jvGtCZVbjjeFWLYZPoURu
7N7jWLku0Li/BDK7cZsJAQBOvWgc7q0DfTIJIepcvGWhf0saJ9/RD7mIHn/a8Pxz
PgEA+PO0AY4RjVU+0P7XNq9X0CjZqeFKO7tRN/i9GlY0FgcUtfnHFplJi1tzjJXy
TcM2li5c49eQrg8g509sCqxYYIKyzMkaazxGFVbxWcTp63ZMhe3fyE1SZwHs81oS
oDB8tQIyw5MV1gkpG6Y5m5IlwVuW5XdVmohoDj3FCEISd1lbgLrVC2xarAHEC4bZ
lH2L0IjQ5wvMtAGhUlmBequVV9IR8tGYTx6E5LiTUYo+cKvBdjiU3VVhSJ/K0Yug
Y//TpAIxJodBI4OeDWlVYhbkLk75xUEl6+fbjcEpGHtP6/ARhuUa3FYLDCc31JpO
iF/byReUxDtXBUi/UWCujIU+Gf9S9MvOTmDsfIhHd8NTvk4PPd4w5q0IeW/tFJ+w
edVVzhHl/ZWDHxiknhVMvlxLbV8ZIyawbj61gI0Gokg4rRxt3shUpJ7jf1QW78db
OMIF2QsWWqhrQKEcJ195b6W0afKcplaxAXHWhPN6CResY0FaVZVIbak/32bjyH4l
bTWTUIspfhgLYVzmL1nHd4lPnm1Wh3R7221O/lacvSNBHCKqQwfwu7Kw5nBdM5wO
zqW1/pkWEt52Tz9mo74fp6smwEsVOTSzItjpWDVZk10QSyh06LzqI2ZmUmEcgyvQ
HYymA2XPdBgvs6vY+eTksqRlCzANHN3sSOL60RxPwuUvskGJiBjmwUhlRUwThO9B
fDD+qNt1PRnsXKvuuU5HLJhR7NgwHJCS5ItqyC8wcRFghY+4Y3uahNQ8x4CWRV35
EljJH9X7or47DiXNlqO1o9XxNqJQNUT9sBl9Mrjr2a6OQwjTTb0botJ9aAj+Ypwg
V2CZ3afyHqWFcgs0gMPmme9dRT9HHTxunr0Bj1EFczIfxNlJnysrHLTKrmOxin8s
TCgPHvMAyn0IDQ4LMqPQbxr7zBfbQRt/LnvQZUJa5lSDQGkPRfM0KckYTE7HG4iS
gHMu+sDtMmMKKfP/mijhYz3lHufKWlMUU2BR4W0sgOYsr8l0c6Zh1dkeLgErXVPq
ZRmOrJNvlKDj15yrrBXWdaXdCgCTdqbP9lBnoLpLZdvEYdLV3SC+CCAFDqjRiH/r
3scju5HEDCKPt2NZ8E1wBqChhY+vGpvyFJ5ozhjfUFjZeKYqiurQp0+IvAUZPont
OIcBDvMgnSTEuelswNVYeR3KWgqt8D7xOzF9jZ1csbYTKp16GmNZYJa2goU3NpQ7
t6s7r5TP1ka4tg7556sIqZScKl4ES4980GfONIW65iq4tsLwgMjyUkJ7cl8vWZLL
9pdXyqBiVKIRsIfa4j4TsJsgfTkOyrm7HwPOS0EasV7NLhK3mIMKDuGnEETIOe88
s/YuSy8gyb5igRxBORi+UTRESPNdMLpmva9h/qQwIuO1w2UyNPVsVTUge4kCXi+v
UbpPZ3Tq2j+dyiBmVPpJxyuXuxzmxAH0ahikKQvWn+LGwdxmDlnKXLmmGPUjC9rN
o1V1eMiyRtR6R5AzkrA40KLHtqVZ4f5E9krL81e72hxeCH8vrfncVteAZiKwZNuN
4V/xWHZVJVsd9lpgvrsFok5B2MIzIaW40D+6iCkykonJEFx2wwj+bdnBm5FHO884
NN5UZRvc1nReWbhjbgiTZY5AfASIEpOehyMNccC68HK+LCRP8BQuYCgrS32Edl1o
vydiCSHG0d0cFKpU75SPsS2mR/VpVHuqqjvOpWTQkwB2BgZU0bIjLqFapRQNgI5E
5NVXOG1YGyQXZSSumTzQbN3M2A/5xRSZcwLORFTdNpM7vO4GoyYEns7nS826prj9
lCr6j1knnZRK+lWdKPNeG/L84jb6F+GS/YrqoSwWvEOSIxFeDHEtF5xxZdDGwu3K
ngU9kkXyLvSJxo6NqixC00H9VvJMU+f4oagpOuHe0JyN2xzgaX3tvT9Feh1QfCNH
XEcPRQ39wRQPerw5WQ3sljw+W2k/Z4gk4ndAs0xwUakijpXFPK4qQCWEAWyviXN4
b6VGt/m+k1o347fAQ5F6OH4HE46DcC/cQEordXrOPLtZuY9twTzd5+9RRa1Xko/l
e3TEWFTln59ZHgsIu83WR9OU9mEkNuR1pUXn1o6Ot0KbzgGUFclrF/3RwAI2q7x6
rOIo+KcNvkS1yHW78AfHEpjtfn3wO38qFM2p+N1UOMKNDINAHUdpej4qxJiFvxMD
5MM7U3nB1Vo7WNSdDFdykTgX54CuCKZ2ka+XeOAci0yMHRmR46L4Dc5/RKXmk4xs
vVgM3oyJf47xqYMhYS79I0YFIFfTbRtBB7TiXCoW8qY=
`protect end_protected