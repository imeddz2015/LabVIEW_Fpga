`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 13696 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/9huKRhRMtvnNqb3Z+UU7TahEoHV+T8U3P3ufru7l1O
3DlgtZzb9QxCbOjthp9+wDkjygH0eUfDrEl1ovhZG62XHZ9McbCWEv3wbOUGMqSw
LxE0C5Wm8ZZyO1mXO+4ithDUQmCgYaypytj/94VkCL9D4bTZl1LHt/LOyip8UoIf
qnkWEoIpbskPyyvpnrLRd6Sf/cZ7pTBS+MmOcOXTAmrj1MBFeXEA4nnR5n4nba7M
d4LahXnM60JTuVS83VANneynowBHjJG6Yz4yP4DlGCrFwNNUQu2kPzqiJy9sihX9
cAPXF6cIXM+K9f3w6/ZHHpmHGZ2XQBgPWZ0ZI7rkNAKQvz8i+OK9RIYXp5yMQmFK
4+C8UkGLz6P+3jwzzz4V6m4+b0G4kEpfreIT8U4Lo6BUPmRuGN71PR1wLFKnupCj
z6IuDpWC/VG8+NL0go6BwiUZ4bVB2Q2mpwhSOIrSuUMQuNrJ2q4Ocvg4PbNdIHIL
FC7a8YxbI5a1w15/oBoD3uzd/7Y0qY2MNs3HlkQUGboKzmhLthSdZtQQ1gVN2dbM
DamFsj0IY6BcpzkVL7YUevtHBSeJD/FJ8p2AV1WZ5jqJp9EuZjtlysZX3m0EEMKf
6B3/nf0+ZuUrGsjaqOKIFRgH87CXCe2BWcVmuz+QmfNTVIeNuzfqPZtTRGgy/4rZ
bmhQIl7kdYGC1bstnbTQ1nponcQL5p35Ry0wDXzJgJtPYAuDF16iLn5kOc0nQYCp
zA9b3TQ3ROxqe6FhZwkaAOihclEbXtO6huCCPxvCoNF/+LKs0D4Do/4xXgY9S6ih
m+vtLNAaZ+rndvmAKvcafe+HZFt+PwEGyjbD71H8IS4g52Z8ljJoKY3HE3oVYK4D
4whDfzsxbFxwPEUJz8QXR4/SAY7NEpFzCfa8rEngXE2s2++78Np6cM8X795rfnFy
rQ+2r2JOay1I5gHxzKw21PnUfzVYd6SVteEpuqJlGcRoZrMAb9r+62eS1ba5bTZR
9f9n3kEUmTPm/Sh/dwKBJxhsGIKdgxITToWjChUWxlCL9ulzy3+0iZ+KMs+FQKF7
cwFABULMkZ8zEcuryYlAg1RprQRBbYhCUbBm9mrIRruUOCgkYmKzdDTSlqdDy0Lw
hWbNCzsW4aFIEeSRO00M7ax8xMW4mVFnAGIlzW3f3Uqwj4b76H0ockn43M2KLBwZ
AlHWdS2H9ilHbtwVxTpx+W7RGNniTUt7456s41+QM78bkXeuvhackmFQVVPdad6y
pLsnQCuhJc/Y09StMHtt85Ku3/kiUZl4ayt80nmp4TdepSQF3ncyyhL5r9EmB7Bz
0kTERR0rd9fZuvKJXcMqZ7jv72ive8xpz0uW49IkLs9BqV34dIn53iC2KILA2ZI7
e7YjsDDV1I6RR/cbVHf4ZeZK9QySFXTbsNMryIuqi5yTMU9fxd1MmVnEpxY0cu2f
YHNq8GwtWM8gW/LnDtaCqbCOlVJ/kZszgk18w4P4DclN/QN83X0ry3bc5C8az0rC
iESi3lDxyb8mnpBGdPh/qQfOm/JVUJaXKJlj5kd3Lx1wD8csRy/LxNfudALGZvv7
1piMXtJmBrACwTIGN4GncmgbTPIo0uP8rJRjVkll5knyP5cONPSKYtfYVGIYKTNW
6CTQ3S4XmKgUmP+UXPSAqhECxF0TAno55GmfSiuhHXKnumTpobCl+/KHA00UNESk
Vac3tPI8AMZAHq8ovhXQ5ARAyaSeZXUQYJXbtWJkHuquB0BFFhWPMdvND2vFBgpH
oPdyr2uPhrHOS6gXJmjGwcn0VuBJ75VMbsDbI/FolnHXBcK7Vpp2JcGFZslSW5gn
tO4CvAc7PqBuKm8tJiAr26eZntEQPa1oi4eHIOxb86jKHBRoMcfMQM3x7MZhZpdk
zRwcMxqaCWoYAduokif6EfvSG4mBBIvcquGTDVuri1mwhKkFCRjvyO7aDNKfYoWJ
XcQEv73LLpw04vJK0GZoMeCBAfgfm3LJgj3J+tkVKrPrqhK//qXCHW3IbzP7UxaW
+UnDIQtn6zJjwIsdgJtpMSCyezTcRTnU2N+Pm9B6V9/SD6zH+PhKlT/ZkTSkQRkh
otw3pwpscLm3JrqlBmAreNktV7pH+s6C4I7VP1YwhSINndahsz4HHNehXcZKSvUT
IbPjawWeDjyfCOBubAOKCtdzzcYa+jjVislZcrUZnpYTsqZkDroogASIRgqljy71
s1BHQbdftiyUoiCGkwz5XkKPKuwCBi3QrBgTLu2Y7dZXI8Ocyx6BE7ZqwJK3T0th
JxbxHF+fE/4/4KdV1VGH0BRnT6o6gfR57tME5WCQc0Wl5/4uYdVBSwJ+9tnavG+B
o8GPqtHf47dcT+dM/r4otj/eHdfPDr1D0n+2QI44vemekRx9qGwNUaZHIv0OCWvp
Lvc/7GHnvT1CAJhix0J7RuVvpe3NNsDoHogEd1ZH13wKmBeRsq9sY/YWv+zUlNQ7
ftZAhIkPYCiFKdV/FLpMaTwoD/Kh3x6t9k+BTy/s0GdG6pD+lpNKGXRbIIZZBdUy
NY2P0yP1rSy1xamCmU2bpeWl4de0FN4CI5n66icgzs9AMKw8gfembwTwC9w03zU/
L2KonuFwfD+H7MAKFtI0GRmDHlx5J2DJC3EySGBK0NfH1vwPMsNBvVx59A+R6oFd
1RmJcs9F8DzSrWV2Ko+sUBG0QWQuYL4eMYqe0o6TZUGTqYmrXsjso6KGA/Of4qdJ
6hKsfq1eotkn7+sAjGoHdduxdUfNR4t9rZrVO/RjBAtxPGLTmqOFSr25MS3V9yS4
8fXs96D4u3HkG2V/owmnQV1kDjb4iLOvEgKX9TuRHHHfz31iTmKlsgYHvdvPXbA+
IFd26pYGCXAngzuA0yfYJ+9flOmJ4oXr5IcgZQ9yyP/uva71G78jo8/+HaFN/Qsm
bkw2xN6Z9tv7UtkWLB2PwfZpGMCTyfQUP/ibRFWtrKdQ0ZSXHAbxDJxuaSkpgCKl
dlEv16zk40prTcwHuzT4NxaTr4x0qhv6rE7VkYDlqFRlJ1Kuuc0AqxrzBGNjB9gn
yoOHxIa000PJSL0tM0isbQ5ZH2qeZZvkgs7tCXvHEJQPmCQgtnrDP/dugTY8Tf43
J90kmbbUC1HLV20b67gl4vwl90CsXr9btdToWtqoFz7If8sf/htnJcREurrijG6G
354pQA2CI1zznhEz73nwPtH7t1xwOqFdO6S2aOcG14JH0QX5OXAhvVAJnhS+qTjN
savmWIYVif7D/XD1jQ2WjfT8opgMKoi6muAmlFRuEBtNsjzs07EmQ9yC+9Crte+t
ehpjC6TUGSuw3JaaYfNtpEkqYfOQImNbh4oMtLY0g3T0KpwmdQvv5D0eSQvkgawR
d7i/ApGHmN30n+l/N37EbvFjayWiYPxsUHVLubDaCVfGawHqX0afzq71ypgNd/6Y
q7Ra1i8yolA9io66olsjK2TpOFvW9GjdmzUKGynGKgRRjVxnoi3176YQFoO4Q5e0
dRNWASBf+iy+zVk7aQ/eMu3uj2Ts3iGZL4cslNazZHb5kTKKyPleEXg3DD4n5P2R
/5dMp5ezMEDHAX9ussB6rb3zMySDx4LNKge9Po1OSJbAKx3E0RsYL5rYpWOfaPsx
AwvEOwoYxtgXIMekmkH5UlhF3ilOOdDE51R24o7dbASKEB5viiGtZOLxK/Otsu68
WdbKNcJyFiziCSb7Hn4ye/18LpSak5UtRzc/q5R7hnAFeRwjvccTxUQg8GmkEvmW
ERcJ11QDsacOdKg+aA2R/E4e7k2a7UYd06xNE4c4IDdJMHtUUVoQTeR8kG14uziw
pG/9eLbSMIQAujQ9fZYazUFW8aUctIA4d0Lc9i2CvySTgiFD2j5UJVvNdPC6zdZc
KVf373CYyV+M7iMUdSJfvVmLERRgTkJuNV1FlYKeqfy+M1Caiv8evtShLtCLICA1
B4A6Oipbj3s2LygHbFJ/h8CKHY9lwICm+Z1JsLpXrp3buxLG9p1o+yDay0RkOjhp
WDNrFYlfBI58ZdXhOEb9YA0vHSLnxEpxTiAdpHPjuPW78h05PvaJ42/wlHsZzziz
RrmwwBWRBUPe0S6VxACvc3CnMGP1EBxh8ZoxNGgu/Q6jo1F6Zgglaw3yKbAs8eof
GVm0hZvszpPGWY6AOsNivydK1CJCo6dTOkYMXJdt1smn4BLg94hS9ossQsA6clTM
h7oGZRfceYKoMlFhsrGaADDEQ7n8exD4AGyLj3cCoJ2aWx1NzAZQAeXcNo6ADPjz
//NQ4PsZNBB3Y/Nthq5plq8mJm+Pc1qcDq5B/RGstIuoHfWnIZUNTgss8B/1GlRJ
yqy8ou+5usZwGXo5Agqa5vyE3fnNEw1C5Tha7qu++UdShbLFsnysT7MoqlrBSH0Z
onIYoUMOAvoj8jPSHlPF3uvz7XmyfPNF1vmNJo8uY2WpoDYq2hy7TCf7Wmnem4qL
14gAEvRGs6GyDGeMzbEFJ5+L59t3WzzydQF7NI2tx6/50endYaVYqK6gGdMhwecs
vXgG9C0S0KIDKXOzUKQBg3ehN94RIx8MPmpLz6EduVITDHpuxKg0lkGmCqlhVWay
PSCrRH4c93EzV3G1n8Ppd5bneo/Cbb+4Kd6H0QXSsk3kx1rUnnRCsrAdWZs8iCkG
rk7PvF3RCN6VGUW6iexngZKjZsHR21vEMRvX9stG52aY9B2Vu2YzyE4a3YYaH5oz
xBQVjQ5d1Ha2i9cIIzutst72q+pUEQsxlHNX+0hMpTFLlH5BAK9bBCST1dKaT1tI
s/v2IwXYYOSabxXgJwOckSvK2fvJ1uSgyHwj1ur9rYcXf0QvbYNUDkbYBXeKQR7E
MMSrvLUKFxnHTrpfukSKngq7jy/G+kYGl+VJy5nz1E5zldwFzZ+AcrMQ5pRtGIU4
tRkHByHb5oUoTWylf9jTe7Nm8PRTphY0kKwFyBM55pXgQr8fVJnjUGOyECflLGve
5eQXTD8ADf/2QA5WS1Sy8FhzXMtUYpFphYw0+NmoGKnMVVnBfXp7WXHW07+LyvVN
kPBqgntkZ3S6nVo/iLmv5pE5Ez90zm99Nv0CTGVFjrkpch0dWjdqMaUn4chBbEyB
tLqB5vGjCCRFChlrsWEDGX9LdVIHeX/2xrAQKJC/rzOPYQX7zrciNgha7GL08UPu
cXCOjfrPV7vCS81vXR46kUTVW/IgQQyjuq3ucuYDQt2WPAwqUrpNMi4G9iHJPnWy
cvYeUP/JYp4ZKkFWyIUy1V5SyC9mY1s7VyJCOsuYBltW8lutTSp0nNssU6OMQsQF
OCN4R8Ac7JzgsN30P+0xRdyeP0E2ybqTRLVTs/FQvem2E68MSlvdD644NG6CRLLK
SIHjhep0BBdbBWuS9u5Mm+Fgc2DfUvsyw0co5JpY5N2gE4YGdQ541SEdnqA1CTFr
vdgxrIxRcJmiuSIRr296WtTHgzBco5rAo62slI7MO15kWLhe4jbdDHgIghDxdcav
WWu1mQgankgBV13jwddR4+HUM0CR/Rd9EhF2dSRlPDwVIypPx3OWkS4EVJusTTui
rc9d5vywIV6HxcdnWbXJ+hPwLmdtG9eRUTyurN3M9rMFQWezq6lG7+mznCDd9G+u
X/aSjGpp9UYzmJaGmwam4nxZ6WLZgVDtinraoQF87ewiRK9/epYTSFGwyEeBR4h8
0wzoNSj9anrQiGr+mS9nqPgragvKjVdUjHs5eLK5EKpf2Hz123mAQP7R/SzmvcOx
OXjFU+ZaA2v5TZeu4OhyL6eac4YW4sJeUyVHP69B0GWW6JZe8vB0c+rAeRI1U5Xl
rCcuMPPOl1rCzyaqPMrWCeNRCNdsR4JUYHOEoWlCUtxcZIw1NOe4bwzg0KsfAdu4
5Dd+ySHmpZ0+Nm7TaSf5nsNZMsoXBy+7rd9mhLZ1Z5TlFBTsO8L1XZqiJH5wre5V
sztQVl/Rte/Kwn8Auwlnu0HknEYc6fhhkbE0AJihyO77FI2tF/dJboq2RwXffM8u
H1pnefhnAeJTopJWWJHzHjuMpN7haqgUIR5Zradum9S6ZUn9Qp7meas+TifDrFyv
eWK4OieZIn8a94Ozxr3Ok8hwpOsZC4Gn+ZgxsibRezgGb8RUpvQWhQ3lk09MAR5R
H6zBoOmwKeJQYAtyZMaAFFYXm2pGyhmyZum0GTyCQF2EVYt1dWUFC5OBWORcxs3S
wF5QpXD7P4Gm+ymPNoV36aASUnLYqlsWjOc5Fs3Np12PR7MYY9TYfhK/k0bBYkoS
97IebQscqyORhGCSnV7tug/C6IWGonNnUJZGS2yVhsu/FTErklFKAXDJCvE4lSzD
nOkPt/aT68RISFi3r3Rxb49WRQM9bqr63g6CemmlQ0Mv0KzqfPqxWh39/KUEdfLk
n2y/7f/dIXQfXGKzv2IL9wJXQjGnY76ufduTLWhuz1ddCBZ86iC5j+MuZfxPgBdP
s1EVmeawsFDwU85cByEdVhKvEqmI/rWcJBcaxsfDHxoH+v7Blx5LYCuIMoUl+1UW
rbNu01DcrAyIiIxnB+v3AJAT5/eB4BCkVmUDZh3+3eFrzAPUKw2Q0I2mMnyDpCwt
mXkuOd7eYIHzh9j45cT8s0xy8Kcgy1nfy3bliJvaItSpzhIhT8XlZ6qEULx1k9vC
Mv8mfec6fUlZtu7rMqtupCJivAggK0L6cK1cXaeUkfiVAM51Y/OEIYqdmjHmX9RP
GqSs+Avw7ShGBSoYWx99Pnlm12wJQCgIrQ0MaW+fS8frtEMy/Bjbk5fmOBftFja9
TVEtdJSylJ1O/M2bnU/cMd/ja3ah8aYIJMf/gfTs0YkjRS2THnOnYAn5HIrHT+X8
EidEdDVGT+Ih1pfoG2vhywAP1beHhNwgx/6bYJu5WUIYjUQe6kZMV5J6nKICL4I1
jKfdTYDEZTXBiSQjuGnN5yejImvKtNgEpYoiMlnaE6IAut4aqq03ndPeP6lQmBKR
ZmC10s8H2m1nwF+tnolVRqMTA0RKevjvFb4CaaGIIEpJ3c5twzyCz6tb9vpmom8O
wDAyWy2063ZdHePSgYoeF2tomSr1ZdUiJP25gKrwBwIm+i2LBOxLZq/7/QEFnbZO
XcFrzHes2Hx3SG6SH6gSWEA/NmS23bukjpeymW86ULarVqgQZCE01KheNxs4Nlot
guuGDIqy9QAJeyiagSXPCNMJ1BzrPm+AglLuG+Nar0Sc7rAgPeO8BXhs9kU0F9UO
9/m66UPv0Lrsn7OUfhVkp8yu4kr8y7EomVedzzN+89tzevF/fk/rgldHIopYHNIk
DSAvXbUTZLuFzIi0l81E5MDrBP/wsD1oVYiYiJODb2LrQkO+KqytrmyKQOPrelry
09DpAISJCWTjcg8ssEvrLtlJ2YyaZYJjxMnw9XBC3nXxgXn7rbIXoa6I0aOc0Ygr
Urn/RB0/i/sbtNXeF21caSUFUZgjTWnIB7LEznPffMMnqsYkce9FW9ldRtWhwZZ9
sWVEdHgEg/wEkSoOPMMhMiCR6qiq7LLzgGKxt9RkDly+RfpZ3pOEIby/zpOOoAiN
rvtF+r204t1hfstZOjyp1+CN6Zgy0+J5fkHefexAW/QRoX+YFswZPjxeBFy7mhMg
JnSwDVQYhbLalzkdrfoRjff600cfrIn86JSVXpdQBjO/Af2DEIjfNWJu0A6F0P6b
zXE2Q+TQP+52EYxBKjxJLPMvSitwiALloBGrJsWcuKaZ/jvYKpCVvNFLhMatM3qh
uI4qdpqXPE+zluU7m+s3/rTP4kxYjxIMoPJf9LnY9U6/VuNXkXYTrI/eXs8PYTPl
JokaijRxq/KjCIfvKesxiDrCmVYMVa2cpIPD5s9jyfbufDgiYzV88nUUOQ5W0oo/
xyiYRa1GGd9dDViA3ts+m6BYo6trRPkwAa+gNAiN2fozf6HmfSrivZ3SzE/nupe3
/WSRYp8SjaPIeG5z/d9exS8isTFx9gF83LAVAP4qqWxHX3gSFmrwBr6OLpI951Yd
ECm4xMvzkvHPXCtkyZYY4U+zLn0QJ+ZVi++YBxDYMEuALssrzugpVl3m58QqopRi
ZJj6fSgSQoZTCiJGCZuVX4wxj+xL+MrR/k8LAdfOUG/q1MhGXRD4IhnekCcSt4e2
teQNSPBC5jdDoFtzTS6nf0Uvn/a7XcFim922hzI9ShGz5Q5QLPyJUm9gAlKIIoEe
0FzqvR9b/eitKNE61kqlhQ683tFoxxBIADa04wwpCTX5uh+wIwA52+m7Zc8I66CW
5VWOr8hhxpSRH+y30WRHU7UJuMQsdYeDRoNIivvt6Cgrv6HuUUbHzX0NN00WnxvJ
w8vbH5ppsO7brt8XxZllOVJvVIlq+r8qM1dsPnuzUkhOf74PyijNhrFbom/U89DD
ePToM9lGm3BnGVbB7F4Rc00gDUabdRC1Aix8aTkH3nKa0a6TVGEzCWttjGwOIkSZ
IR4j1+stzLbtSS/LgV+2HR+xz+nKuIHIJNy8LUljUANriLfVFnhMmuUXcVNin5Yi
K89buFDAVjpfkEXQnghLnjtiezqou224NuwVklEojZkZ/+Wj6c/dSCa67KXiVPd1
C8WCYrFoUwDDNylIoFEWwjYv3/YyieicQb2dp+IQRqTD/xqz3tgwZ21cuvDoa2MR
FflccQfYRM/hwiLO5VbNbf+tbHRUSaOteKXAsHF94sLimDdfhlEIaQ6bUz8XHV4d
tHdvrU9mp1IO+iXL2lHUh3BKNpiz7kfy+LOrYtprUcGhQTVjM2cYYeHw64TdGcom
8/XEq0pK8FMf6h7/Y+mnvTx8PPQoa5ZSVicwbddbsod9PixribWmpdxs+q1PPqWi
wT7E6mFhpVwVYJxKtrRV36ak/QGUXPRhxVXl9XQp/NHc5h4zwjU9WMID4xgmQLNf
RTdMqZtszZeSaZbfCGXavLJFOL/YTlTA/KIijF65k7ueuiCyJaY6cLfsFKVLmOrx
poulTfQLkkSV4ape1qlg8GqnUNgabT4C4ijtMHsyXZfUNiz5ETIzVzIVxCggCKnE
zqJPnYqpEHZqAAW0QAiufTD7TtLIRTWdSvzRhiEOdFpcor1sCb2BVWTn7SOu8qmW
d2Cztesheq2kcx83063Bu17omkZJhpWYMJ2zUpHujO5H8vBd5LtaOXaLMAOYUx0e
ZJuq63n2f6sVx1f8sS6NqEIhlgMdoRGV2SZX+a3J5dvz92TPiQ5zoh6gW0Iy5T/3
eirVksaKUpIKDwkUSpmdOBtibPSAiU4Ii36H/qZiT459Q3lWBOhSmphDhfYiJpKR
1H/gqhk+pTv4EhHTYrdNz+GvV2xxq0vB3Jl7nM3QRkE87kmYpyZ1dSHNoYPsyDsC
udQgvvv3jVOXUWcJ59NyYgERr0UsiJSzXvIqIwcgVUeBLhroH37b2fj1VVp7N4TZ
ruYYGFe/ClMmZRF8rTvaFBpgi1zJ/9e7a5+22Mv+vrit4ZxMhH8Qdm+XSqZiK5Z4
o07jKTpawemh0okYqwYdLD4NNItB/HrFxx/H7Sk4NauYZqaZtxaC6jP1foFiTv5l
uKlWYvylEm1ZXIYevsthAMkeDcaf3IZzx7gNTy+r5rlCuSsLUaRVDcRPLBvjcRRV
Oos2gNdVZBcG9vhgn6ZV34fXjY4KfMuu8u23/t4+h26a428d/TYueHTBI/Q7/1qN
cMMCBueXyaSmOM+tLl0TsX6+TCpVYpt6JguQR+BH/I6PLoHBimWZs5uXeYyQdltc
zN2u+DK1+PkcKtxOl1oU6Rwx/IZjL86ohrswpMdl1cEF14ZReNcYIN0nzfBnmIMC
/YLf6zsK0zn2VydKy2n17tHZfhppNGQ/PpMaM1iPb5pAROVw/PyofyJcl5A8zyho
AnlH50LVmAmL2+7pgx9TPkohOIpccuX5G3LSIOiZYw6Vfv5S76+jY4Qd1Phb9Tvb
T/eObLUAh5i9wKMgkJ6drPXeHhYLIbyR+xhcTp8RhPvOfKlfsUH8t4g2Go+3wQ1K
dqMVsMKMwdO6FnG+96bK2/O1v8YN+nQ5lQea/NmoNyNxWBTGCBNIfwibv3486KR1
EBrKahCdx5xCT+hmI7+0d+0NxN0x0mjhYRz20Y/v/VPpMeDmSPALjj44SeKS15s6
lx0KzhNgJw+3Q07DUu2YetZYDMQyFZiI6osX4hUM0KLktJezYMnJoIhoe0d+xe5B
pk57x6FsxuxmeL/lZTmFQ4i7oF7XYimQxbjnynAd8+G21XcUuB+AfdlqiLMiiUKL
k6BFJsPv6X1yLHThGPWTpy8Mwoq31oiwZR1nXt9Rw6d6rOxF///F2Egp7G0j/bDn
36GR+9f+gLTQXb0WeySEZU23VxyZyivCg2LpfmQ5+0cL0mPh36bPPO38PH21yW3w
6TjhvbAKWyMkwEhPPlpx2ZeuwGf5ktKG3QbYoLtshQlU95IV8726vpQLwowwGTyg
OFwEHHv8DJwhf2Kdbu2AAZbrrVkxkUbLvR6aEXjHtZd4hjZ8xT2DBw8O72j4NrFJ
GTzDvClbPPiPUsn0Ner/Ny416B4Xf1YM7J4k1jW/i9FHvOFa/SsV6CzDiqxrM2d4
izCvUulKBrfLzWTEOtlFNsLJ8abTqkxSV8xdmd5cB+zriPx/EzCD4GDsAuBNvtE7
JVWST5XQ8GTCacWEz7TY7a7qoWqRJj4UH86NLsKsCuKRWiIDDnDLgZ6PUhWD4MhD
K9KDwmGPrEzFmSxw/uMqHpu9wz1C4res3S5PxUUzeshZb/v1L5/azngjv4yrlejM
NGCH0l5dshlvJ5Z9s032RQOjMYEVS1szdEnrFFF5cH5H28CoKUexox8yUt4rSXr3
3jn/wPNEoAME38EAWEl/Z8m1fSjC5XuXW7wnoumUU05cb52IknFJ1cYWnanfPjLS
yWhWnpYHfy6iMg446qgHzh9V6JdwzXy4Xv4yKXifugXjctKza9EoO98AcVuP7Den
XftfitXQW8v5+dKxiV6nwSyxs9cbd3zRHc4Gh67dUedbQbTbIVP2vGH6D1Y4UVa1
tvc+XmGCw0ZbRGDnAESAZx+vg7hS3kbu460NHpjlkhRNDL16ZOmV7XFqzXn8odEt
sxeXGzbGPhVsRfTTZzlniH2rqUSUM9uGP6wE0YFLDiqyJWoTSr22M/hDu6MdWqS1
dCzvTGJrkvY81N0zGdJR+v2sJh5R57NIt52s3xRvvpe3rbtomRoR7TDmx8IWWfsE
NJ0mOg/QE3VTzZjosy39XwBKf0SQG4T88MWfFtTVFceqjgCJj6yGTxoX0wBCVwxf
nH1st0OP6Ckhr3OOY/qZhSHhGKX+tnBsqLNGJ4SrTkvvB08B0T9zHYeV6LziSF7g
IR4AZCGJvjHBMWyGSb/EZJ6G3bf2y73scfcltsZmw5KyF6hM3in5EIZKcmMIfLZW
hxhwUvSm22mpqdc+tB5iz5gdgsNQgR+xV7EnD76zpCW9Sad+9wBJiyVqbFW/g9Cz
cKvCZszhTJcxZudtVieScbhDpKvpH3R9unCuPmlRdRtzj4r+tl1gRbvFVDd69D3q
BCidc6Dv3N5IdpOezOlDXsJxKj65lLyFahTHTedukASP3ye5PrU4tMmFODi62xH+
HnsY+pjtVlIsrT7rDbrwdo1Cw8GzhtsdqfrnfQyqXo+5WGla1n6V0WwoM6tc1jIi
uze/nbFoYCJx7asDGneQOwz5lezgXcO3o2yMe9pKdAbASYcosRLtPp5t5+UthNrN
BQMMYRR+ky5b+YDMvtp7qCu+B1LEIevzbN2A+0jY+TQm7aeiZN1CNjNzftDqbF0q
ZL+2lVttP9Y4Z840DNCdbjR8eLQeNVtojEiEf3XelL+5reFQeQh7TteiCSIR75Bz
cd3Ag4APj2MAoBo1x9B1MWHHiZbY/pzz/HPH3q9cQjmMQQeHFMJZWkwkM86lilz5
Ns0xqHnkXQaZCyen3CRd7oB0PeBLsjVG0b3gWN5E7tqe1KJm4W0FOBTeTNQqlzqx
f5xPbnORW74WMCxeun9ePAVvI/opsY2fsE2H+EbnifZMBu//zcRl80Q0UJsM2/0Z
NufRb/rGVLy+1drl/do1Q2gz5evzr5qL2Kb+kGupu79sbGWlGuOURUoORecV4tFD
Ka0ZBE+ZjIKnnG/LIcTMdMkizFRoGBENGgTnuORxkpak26NoHJsPcku76jRvEHap
vHfKLSAxi9fhgE/XWyObtmHWUbKJfxG4zj+45u6G/b2PrkTdfBWkEnHf7XwjocSE
K6nw25V2kFpjJUp5v1gXc7uySK9G81WHkZXDmJ38tqfh2lepINIV6s031GBBAYwo
Y4wjnCECfi9PYGIGfr2Ch+PKtVgmCmrVT5cmLAi4qzyY2CWqrvAmLFMoVJ58FJ00
z3SSIKGbPcVDQnWC8uSX1L9C0jghhmmz+8Ofz2UNS6MchGK2ENAIrGH0NQIP7r69
eAM4vuJ1xWDNZvvXwQJF5ox97y1eYbFOCEuAuu21uQKjToRQYAesGs6i2s+ETprq
JJ06rDz0SIhLmNd1Fj9v9CThjiV/8p9bTiJxZ7/dUYqcHYTKWufPsI36zgKIVZoz
h9lJy4xY/WJPNbIRV1HWqZLxVgAdBq/88b6R+5oOob8xCkCJC7cgil9r0OzOCjxY
B3bFE/lN0fDDd9MKkXh5y34FMFi5tw1tm6dzSosk1hmiQOUy9rUyOenO3WUJmKaN
/Bru8wFRaUR9L6tnO1R84PV/wkBm+oWc06XIF+ywBjPFomdT78UrSlhqrrRl68Ft
l9Xr3hgn5s+iopPvbqVt7g6T+96OXhBz6rYj41XpmB+Sq8O1hCIhnVRxush5Sp8k
hQZMPlZ7FjbCX4l9iS9kpJdVEzPJl0ZQKYqBxtkdP2BxhnZqJ6Qj0qDWhoS85ySG
JQAyztpLx26gxM4AjOwy6oL9Ikl7qcWZYHExn6XeZXMHnvvlShzo3iuQyN2xgF7/
BTVg3GkfNXVcqm1VWv2iRzsrnzeCPAczH8zTPV7TapxeV99cuUJh9ZvKC2yOF67i
/FocPEfWMB3NgJpMrX/pGHI9mCoG+cZ4pzlrOihB5sACHvrhdbw1Y1Mz6WJk7xZX
btb5M6bqJJg+ETwZKNzM4MctG8TrasyfLZrD+8igYX9Smp2ih/fAQg9HYLys2sSE
BUgjWtDvG9PgSDSqENlW9cwJXpqysu6zuEe2hHtfCRx2OQY5N34V1XVBhC2AdxHj
mYX2Nusemug/36iKwVw2mELCHyux08mCHZC1PEHAagvtPp/4ZrHopcXGyLEQt0dh
pdbyvBdc5id6eSLtlH8h1rfEQ9pYnljOUnAWmuym1JztJjKJ6B8TYYS+psYIWPrH
99t25L0YdJhVc3uobjVwgY1aNiDtr6VmnY2jmmH5oUOrAYIpdG2dFODpcmel2N4R
nQ1pdsPN2QkMpa4QcU7oZ9+sSst64/gHNFkaTBKjStqZ76L5GQDkwKW89J9NS8OH
nbvNEV/dzcOpI6yIb72ooxgIw1e49c1UnqZXGC45hDnEexooW5xzJa135Pt2RP+k
OcENkeB8tJ/DpLAiUaKvL1/4yqiitLYYQAxiNdjzBI1pynfTZKq5yMV+PPSqlX6u
MgYUe/azV6XF/ye8FtOQTGYBM7CuNAH41KY8vf7o0xGtqmku6VCob9ab0Y9G+aaa
03MCySq4L0DYSqANeApR33mLAeFBcoNxdKXPbAUybjX5jt6rHUzmkojESYWZGxzy
8BsCnHKCXD7Y091fRjYRJ2bNJxRbXgbzUo5gLfFG3OAoXA8lspPDG4Gu3oKojSkg
MgL+E01QqVkpOikSGkqqxRJUxSL5IjHC/+5dqQgYqzt7DMKvBZJiJga7SDCdu67l
M3PFrazhqlepu8TUavwIHVUpAAXI0DFwenMcqkDcQEe06UuvaKV5QIiUrlvVmohK
h2cx9YfimJhxsqPd4moKh3vSamE7jp8IBbeYcX67W+P0s1fEHi7Vdq7uogjGB3Hf
SxfMy639oB55KEinuO1Zrx0NwkH3rZpIP2VZZzuhj6xzswAwx9eeliS68RGlIpLj
pU1pLHdviQXZPHf6upU82Dx9vTCwCkrphfmwCP3a0pySoXj+X6Fm56o87RD2QAX1
Ia3e5VFa/8GRfS8yOdP+IVNeOAJTvcUuQcBczdfCtt684LMP2FP4cbVYNW7AW6FM
NzcH9XB7o9i23IHxbcFTHAKKwq909hiWb73X7/41MwcG+H2PHoAdrAgCywmPfxHv
wclHUutDqDYiSo3k/dwV27GDwAdpVSSrSG6B07BmmGa7aOkUAhMT1Mxk4QWpqsrk
8Fsvbt+FEO3NuFx0zDb8GblC/BO3F+b70ZsBgp2TdO+6UWkdjUCxceF0i3c9FLyy
9c/H0LDUxe5JTtryD7XYM4soiO9ZTyZA4nEhnQANKBJPSe+NZnyE4yGSo6Ypc0c9
cVj8z3U1QGtlqFSGi0JBW0aeYJYM9onELht6Ix3yzK/39fdNtVjKLwZPxjCPz1GK
VdqNf8EsC/XOj22UM01UFkbBuf5bdj6HQv6cDef11eSugiq+axoXYkKNOYO5u3AJ
oPPxDjAJLmQVbgub4i8b4gWC5RNG9JMDcgGI49AFLVI96El4ZgDg1o2XaP5Bfsse
fKlYx8q1kJIOfSBlT+RsSjm6UbAQCdjRcf5+Zz+4+4jX+GTPbki/69hA0jF5Ov2v
/UIEsvj0qVZ1mF5RwZKiaQkZXUMKm79xLkOLRYZ7zjMY1CTldbX80DUB+UF34C9u
1b2yxRRqhb/haqwaJ0pxxofguyysVPM4DB9Kw6RagntnbYf9Of+uBiIUSE7njIMK
MdGIrGNZCle3fc3TLRId5vom9A4CCygCtGEnAE2IEawm1FFf/c9kOkd5PBbrbSKl
vtvmUQB2sB6ORm9UuoYuIBBJMlfg9Z5ODOWgsWXMEXYsqJ3JCzHdaLGwByq1K5/c
5b41oA2gITZoC9PLs01l0POPLAxuE9gZFxyfe4TsT6Cz9qwTyeTh3PIeO2hQFIi8
PmXUk3w4k8HwM3zKCREh6L/9q8WPGdcdSrokvndggKGUpQ48/NNuXhVo9usYJZ+z
jtXIiUUoZLpS/RtmTePe5HGOx53J8emVS9W2yqJF75bEn69F1YDv1P329yjciKgb
Olujw/j3ZTYhg3NCPF+und+dV+TpUwxrLBKuV4xtY3JlxNVDNMcij2ZgEChBPKq9
HVVBTCmMGuX+1vRZg88hO9ybD8HcEkpwe1iO5y5+Wc0X2LHyQxhKYEKRm899WVIY
m49CVWYNKGGUT6Do5/pU+IVMMVtE2WptC4NlLRf/Wow3DKVTn+Cd7mKKolVTu38+
9auTWHQg93xB6ytaub1G12oiH4sx7p93OUQOjn+auHWCx/hL3NhDlmrvy6OcYPyn
rcA/bsyfGD2Q/2+D9j/+ZcHFkv9t4q13r4VZlPYBgyXO1mA573GmAoVHSd+u0dti
Ph8YcokZACKpNYZlrvXI5x7BKteq24WyMc0P11OxKQMAyUFAZ1MC71ZmsgM00H+I
8a3klcdvBLVTd9d+FtbrVjVOHJ8vjyeyzmnCbc2glcau08GZYgWQFjCUJwYVj7tN
AGMeXzi9Kr5TYxI7Lre3DK/+paRPER0ZhZho6D8R+NroQ8Z39EyRzFywhCWVP2Pe
ShPIgCT4WFq5VPwumCR4NUtXMtgTSFozm22aPdX3W6LnH1uZr6kyj0EKycamtxer
kJM7lLqqOFMkKU2l0LrkMLg2YPwaXn7sj0Dsc/SKdooiRVMHz8IzYaxE02IG0+Tc
XirJ8PhVIyEQF6NCGCvUhwi4adBGGD0iAjlU7m8jWFmDF28IZlRhJCoAbDvzWDw5
wFFz3kuUbbtaF1Ik4DIWz5CJae5uqI60Zbbvugm/VjAQv92JKhpiV3uGqHihbRhk
iJx+GMdG3GXG3a0HqjzWB8c7NdZe/nRoLLUaf7MIy8UpzXHunPBiXINabTtRmH3n
SS3LbeQVFeImW3ege/hllVCryEq2dZJQ/vNRqswQWQnYw+L+QI2ta2tZSwEsaLvM
fv0SHxAbxAykp30BDsJdmTNtCIqOCOoHw0B2zT3cy1oV8VKxckHe01eIpq4tu3av
RPo93wFDQxdWK6rTACzyFO1j1ObrCm119GRXDqFmscMAp6/u6sT7fSf8EshUC90T
v5mLlr/joYWP+NDLjnqBQvd8KNR1oI9BA1VdU3xuJe2ZN8E9dLw6ktZ4n75kcqHj
3mNSC/5dz8mxjb4zfj5hHLD1X88piO/LmNftZjWMGBYgzNN/fUEkjwQK0Y8G/EI7
Azsa2M9c7q7t5rv/a5nx2/dTFs2PkwSu/UXDoWt6ji9mVDROVIU9ZFbWNY1ff8Uc
k+dkRFnLu0FTTZc8i6bjOzDcAlw7jAT13jFGuupQF9olKGFwEU9uD+Nq85N5b0m7
uc0QaYVGgvavrtfr9mtsbVeyljwH9DfUuzqOJBaTI/ENCZr/aMcs0ZrDAWGMePqj
1uGI9YPCYSeGgvXBcIFpEq0W7YdB6ZuufTiGRVZUcYD2z09BpXkTEF82KYMFm3YY
8hg3/bSZbRomUViwJFpN88i3OMqvvwXUAbNpkk97N2miKJQjZUPEX/fGBM/QrXUd
qqA1cgSrsS1r2mG/tqEvGRNXb6viNDb45x7HqelrYOu8dZWYan6n3DIH3Z/63wGM
MwcPmVvGpFAc35+ChW6lFq7PA3SJr9ao5qJnlfW8JyNh712Av1P4YJZSKlnVtTTv
CSC30jj525NF1AIa9IHXsMDm+EN5DuOdTftnKa9IL4xBWE2O6HRkVpfAFRU3zM6i
qn0o4B0FDbLrOcc6YR4mYuPXGvANFJ76sFfDRNasjDT1ui3YSU+fEDiJpBNvcewl
TNnZNmP/d7d0E+E7nI1ajRPrAjk/Nu+9fjtmhRnC4SJT/tznFsXul/oNkyJUjkHK
LriR979j0HgeSpDIuQBPO3OqdPS40O+A4NUnXnfrylGvZYq5dLZTsDm465noftba
zrZSobMfd0AwQ8bKoYtk7+HVykCaHqFQx4NvgGHexLSdIpI7jrMukkA2Qv9okkDk
DyQbOwg5/j5oKUwlRv3yMlWkJkAqx9620GYI8uKMYTrOxYooP6ETI+i3uHER7M3F
OaqCiexmifl9yZmo+9RW2Aow6pCCZdV4Ifqx4G5CkVWNRncg7zt00Z/TBvb41cu5
0JrG5NwQyF3RxUGaeRaFyCaLpIsapLQ+YgXu9Z31O9jYvaA0ar6iJPJtFr7BgjY1
6n07mkFvkiiLEtkhOZRYWJCdx+2oDUoVioH4pJtKZhjn2ooQ6vCLxcE575Ym0oLk
orN1MhGhdd7XlzOkl1MyMgD6QutLGxhP9LAVDRV+QTgfJfLp2D7vAcWBCB5OQ/fT
nu9UwZVsx6KUX94MeeIzCrfjl6R+jaYb0NgXQ7LcMb7dCkqSvOQ7tJLJLHP8XUtb
cS+kfHIZ7Z8E+ZdgHYHvltVw6Mt0WxzGbbngsEq5QTRCHfYOxkRRcHqH4aFn7kHe
bzWDU6fxFNi42jzRY3mltT/+IU93FrcBTa9QUTN5YkCAkSKBA3soif+jJHyWPC9Y
AgYLlMpiBgtPmooKTwU1gEFJ3wBCVxsSKICj2e2c4LGcFtlHAXM4vXws9Q1rq7fm
IRv7iE8iuxv5mtgaWfBLWJH3C0v7e0hXAnQZ0EidzCkPNLCXcvecoEcVvEkYHJjI
NTJIZ/7ErNnJmzthmHyVnqCNCpdboinfVYyBPrZ1PvCAXqn9bnWiSS2gxm03XG9O
cLXv8yLEduKcnFh5V0NMdsQloL0xu/LEbXJKRZBQgd46sUGYojlFosRXCuMRHn4e
FyybC5QbLXb8Y1QQIVQXV2hf37Fkbg3Gpyk2lVnvVzWjaoLP23PqxQAgTU0266h4
KXKARcpBXlRuGY+53RrityatnSsWgA6B3m9VU9Vfr+w9jce15moORbYC3BS6K0mz
FDkW8RgRvCxOSWexjYrjv9CmP3dZPAwb8ve8U37u3B4KBRWKzXmkW4OlLTCWxtUL
BDK+7y1rpRL0WmIT/IPsC4bii1pZXDPy4R2Bxe4ei/1Q1ZSs3NKWW6yb9M+wNyx2
ORJP19F1HMblV4MvaF4ENHs0PwxQrf2aBmP3T/dhCNV8dWk+owMup7BhdbKJx+ju
7wfpexRKU2Pvoz2QMnWmnB0/XSsB4mIpXZca7UkGGUw60zjmoAXY7E3bshmLbOLB
NlryB4CKnc/9GYXKPfyCkOpg8X03S1GHw8UYw9ABlSl7Fvm3movpyYRY2aG2GVx4
pg1GAHFizODIEVOc2vwGug==
`protect end_protected