`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 11088 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/9huKRhRMtvnNqb3Z+UU7TahEoHV+T8U3P3ufru7l1O
3DlgtZzb9QxCbOjthp9+wDkjygH0eUfDrEl1ovhZG628TVVFU6ho1d4tuEwHzC7j
b5UyB+2/lsQ04z2Ad6gLkDHTMaWHdbmuhbnqYJJ4q5Jitk6XTqOygRTpXoBd0zgB
JfhOgmQjqlLyLniRX/73b2wcJqvTasEO3g2/p2oF7Q4l/W37OLePsbDoH8qGVgiI
ch1kgUE/FqhDRWgzSecSgq/XWar4+e7IsSan5B8rDIwTvwWG2C9NAQBsS0bKTTyw
8X6JUApcRPR3w8NWLF+tAz6qkTi0OCUk3Tglhm392gF7F08A+Jkw6hb2A1+LgyEm
USF2v276ocqtbw14NPHtuVpV+oYfVtHbhFHETpETt4R55eXT8PPlocwa7eak25SU
Mi6FWo2kgctM7fj170c1z8y6hzTE/AwmslPD51c0ggSlIyfvXOyNTDRzH41Ng/oZ
YVQeo40qvlAvdLCAQniAFtPkq+cb7zrqvqMyPZZdhhgn+UPniEVs4TVsp59WxzAz
kDaJw/HYS2XaaA4CPrLCenJ9PxNEgH6Tzmvu9IPjKEZ4ixoG+ehSILRdqvcsKtef
iGEc/HOZf8E4Hw5nZirjOewYlujhHBYXmAHY0KYXATDcqMbfSESd8PFQ6okkBtgk
ZQ4faeWdXSrY2pHAdiMFxf+K8ZVRPNdwJC7mt8W/YNDndf39IK+7vhZe9Z/CaONc
FYfjp6zMQh8jN5xvsbOVcCkQ/MQmjIA0HlDpYgwebxsFE+8sHEXhOadOy+MkTRIp
i/j/swg8ugQe+zzlDOwNQzlIsBkcRWMmVOD9qv1RRbU7q0OiJ7We/SNgPeQ/gzjm
tbW7rqUTW4f3okcoqbompzUvec9v1Ct45p8r2AH9sJBTtUsbT7bTWuexYalkdtI1
pvQI3ynlSwI4Tnk+TOq2IhxpJnrqY5F1FV91MXzea1fUSnnsesQhOOJOkx+xs7mz
HZvIOYwDrJMHfMOCKruA7/tt1PrIwTglcVtABrog98ZhLqrOZCYDv66yS6OsBnbB
a4LobaZt6VID8S6l/7YNMFX2oRSPeXhVnSIwyFfZIdv2cwofN+9adUXGiSRnOCuB
IRS5gffPpJBcdwSegyH5121uYHVwx0vGYfrmXU2SR/Ahzhm8tBa97+egP2kNAGQ8
tO6Rx9v5o0E8fhYEmQ78cRxcXOStxG6hEUBrv/mr+LvUHAyuEgyC8EZf0+EEAJIJ
cGtmcCzcGu0okAT7Ecyx9/m7luB2JApjn5YEWebe7LmCUSvW+TpHTJHvu6vTYyVW
u3mHXl+MZV8sPt+SaIxZMSsAMmVbBNhVaLGPQIY2+nxJVRgIFq5T6cOeOd/cscp5
o2ghXeMfhGajjJTByOVKYbirkvVIzcxlZg36p5wvUl74K1t4IFa1h+0Kn4b1KUMC
j/rYdowSW+dwB5vBpAdkZQPQayrlAXrEwOfoyeWLJHBEPsX7oWXYWWILeKW8Qv/9
OmDVnDFfmei0ZffzibehztoyXlouLW8ouisYlx3XI6m9rxdLI0cxP1hyEupnXvKF
fhI687ep2CJ6p9PGm2rAEUpMFFM0ieMn9ig9YIXAxTHt41xDxcmw85LsH19komF7
X5aHM/wCJU54Qu23iPGPDWhcHiGVsL00EzZjc7rcBk6f/x+6xlNBSyMrJ2YmqZtr
PNP2ShGhzW9HXPSvPE3ZlC0bkiMJuUXAQt35A8lYT9/9UhbbEbJxmtbsAt0iOwc8
SpDfnSH45J0IxYh1iA3ay5oRvaR93EBPecfg7IlUM6t1qrfO7yT3i9uWjc3k4mCC
vlUWwtXmRoDi0iHhapL76oWwFqOS1KR9Prv4B3nYkNksyHzdzLStGLwGMJN2vGly
2+xOhy9UCGctA6l5lf+kho19W+B3ry6bjzhJYF8uUtzJ4qkHbZ1TgADXVigVMiAb
DGUR+1RAWFgxXaOrSoGZ7Ztsj8ZDMu356Re5pZiSlZ2O3J/Tkg9PYvy/NHwejuGF
xceKVu6LMnloH4RO1dypCBsJxF1uvaRC5AlJlQTn3STqtEfnNwtgYc9izNkPfuox
aUck9OuLwZhuDRx6giBFg/M8KELcHwfShOo1/8GlI8+/lJzo1k4rd20cybZwDxmv
aAgTKVuFSaxGdaUlhuYH9m4I6A73a2rEbI85II3RNgt3Kl+/Q9ClvdGWHQWg32gV
RHXcOm/osjypbDyY1cI6uXUnGISx+5XAYuxBML+034l9Bs5c3cg1GVnmp3F/XpCn
mg6ZnXoGeZwcw0kB8Yu/C9jndNJORMWPhNxzEAd/DpldK7YhUqhh/zAuDMeCjHIr
bJalLQrK8+s3gbYG98kY+PmBQ+PqhhJfJYaiZDW3JReveXWAK/+bD5T5o7DpRLTo
AVm1wqT0Cz+M8bUznzN+l3uJUrCAkPsqMF3aQ2mzqPA+7n8D0sS5yDys7QnNxKbZ
d+1GJsEEeo1T4FfxCCQyMZV1yRmw0gTniMNcytaJfvkq38x31OgfzJGd5Zf8ifUu
1NURADrf+4cMmhZ64/ZaLPcS/dc5xFLq10/r6KdoogfaMiJSfKAMJi2qtp2dVJej
nyQ661Y/GSsi4KM4I/IMzJcuYAnvmTjErodSqMCVSIWQLeIL2Q5OQLKhCJXDxP+B
Xa/y86mggpVw3eXr+1FUI21t9w24+p70vG64pm2cBa6II3nckuVF2G8Llq5Ld3un
wS/W/Lz7Vior+f+9cWNap4NAA01IbM3O+LKsneB5kk1Cbo86zcFgcY6scvopABwC
ulrus7hSjzrArIIQPw96b9LW3m9vvnl/Z9z+tQbpJX6PSIumsl5qh/O6avL5cRxP
tDlYuhYGpU4NBqTk6yEy6k44vdA8125VUJQxfyYv7uhe9c0501PhOICnq5zFAf7U
GdANSFtO6HAOP16IJe8q3QQKIaUSJXuIcakCdhcuCj3KXAwPovcayL9emepJTec3
xcVa6VieQ0pSOji5TftPP0XolqDWaeTKWjeF1sj0BJgBR233FACewOkOgWGMVfQ/
WQKKevPAJbwrxheliOrOUpUGat0HZhQIA47UGpkLGN27dtWcUJD75S83sQ0bjB+o
fw53pQxPT/+54nrGyefUWruhGS+XCtNSqcfa2kQIKoljdjbBRJw4D3DqyqHc4Cm+
4Iv9DjVhKdr8VJTl6OkgKHN1VdDsjypw3gD4cuZd8v3YsoavWoK4BuX0HOyoc/7n
s2fEB1KFwJJ25ENuxaKO2kzFmp1nFTynWZzrCvp5MV/okGAMlI2IxOENDhJYk4E1
cYGmTEaEleY4ji0roqednkZcwLrhBi5zqDSZ14lSDPcafdKnK1zyrquhloYSMzYs
3sP7t3TYaFNhv2bY3ne4vSz/vF6Henf2aD3+zhV8JsAhxCzU617eyo3Zm6Rk3vCW
PVycW24WEeOTWQA93FsaQtRyEpvQmT14PnqdnRGWBgbs2/uGBBLD3IBhpt/uN4/5
dI5zEp/fITjO8RShlDxNMiX7rtOpgwKwqLK6jN4yX89uLrWuZ6GU5EekXE4/70Hk
3W1akAc/me6Oa6iMlA7HKRR9VRSKAs+yd1zvQvX4E4DVvmG3dyRzE3VD3s8eliLx
uHXH2hs/CszyQaDa+Bum8Jn/zVE0xRN5oLl9Rn3zSufGC3xpOVOmCsIBaBQytSem
s9UFVT6Y++mvJUYyRt9NCb4WHmFUvr2QlFsaptGiN/H1aPqQW9s/bBlvrVDXNcw/
rHSP3X1HktwF0qylReq2pviDCfCaLcOWGJm0wbg0o7agx8KhuPLwqKvweSht+Egp
vuhVrFoCoPeR0e91OnBvBT2oehigbzDPOur3PWE/GT8b4XDghXGyi6mmRqdjL2+x
zhHT7XiTegxxXDcPh5M/WBayTKXMfEgSxoS90DxaGQV48wzzotqhm+lPBZgqLc05
TzAO6VmJiTqWKdz/lUGaBTnS3r2moJegi6kNUeSx4FfYeOrEQc7V/2uiB3dpijdu
GzEVCmzH5dSSHqx5sET41oJyFav8KYkcWHgCkJtUbRiKwJqDMk1dyg45bNqi0ZNw
kmP6mB0X0YKE+/pQ00ODivMcapQ5NfDoyLCMhdU+5zKx6S9wcJX7C2QPZgmcIc7E
Vu0ODbmYitnd/+pfoZbHows6vlkFOI8srFOHwnsI6Q11PBi0qXrozIg/ilRcVPc4
tjycJJBP2qGO8QSvCoOiANApo6JrcsscSw8XDJk/J7VDf/f0tw7BrS76pWCzAJin
8N5RJrwi4KJE18Uj/tncn9TkkOkN3D+RXg3qtftsucbL29nW9wLzb3SmpE5PiSHL
bReP62MSN+WE5K19Gtdigt3wF7kWAI248TwE4L795aeng6xbNvoMitGwfpZrSieq
AeS5cy7lg43piptt/6+tccfSgSGjjTnShBT373uooI2WA9p9TGAnKc3ufRYKH7Z5
zk+J0lIIH2zH9uJSyWdvfKqBugRA7DJg9M6T0+KWksmgdFMFYqu6URV3XuYdMg7l
5Msb7/ip6o37TNwKk1NvYTqjkOu/PpxtVF3WDUG7rXV+qCuliES2lPIKsfMbhYfc
xZAZeNfKH1wUCdHONQ5FWhLxQDmtjH0zGW0VLHShp9GJfW02GzmZCPVC6nNJj49L
u0dOoT5u/pt6kjb57jSS7gFe1dfgkjwRcwEy57LwAri3qZ4N3UZpwZXERJTh0HPU
DzEGSzs96xsMXuC80SmT5PTozLazDhPkuHvIM4EVcT9/JqRT8MyefHBxg212htxD
4vSEG0PwYUzwvjaJKfZHBpXijX9ONhwWL/A4dfHd4y8Zxhwt9KH9wy6zhPHOpcsW
kNY2oW1ar0+o4ou5YBfJtE9PujY5Sw7Yehx7j+s/LrPQ5PTNxaG6rmJ6n/WH6tR/
1M1XOPCnbdYFULOatIh0K2Y2pftrafSUv6hNQ/qUIk4H17BbdFNhpiY5v7PUnQeR
uhPIAsTF7hHnoq0eOjhne5xV92naphSKV7l1W5/+JRCLH55N8cZ5tRlxE4Qo66G1
oirre2JM3wtiQGQiHHmOAq+i864LLU6mfxrzfHr08oAaqdwYfCJHCA4MLyU/TAcc
VovK9YROh/J9GoF5bDlrO5Luco0/UjVx9XGM9px3jUaPJiebgXoIAjP3RszgJpQj
230myMxv21WUU814zCviPJJLrl1Je74LV9wwP0OorZ0mh/5f4WVzZCNPs6/rhyzp
dCFrce9N462jAlUvq0gg4cHzkjy4VUAjPN2OCyoO4XVJEJj9vWlGvTTyShpXgTz1
BfcLDuibeFDXwQzeWjlWAwnOsRgKcoMXsp2FOfTvyIHY4MZDttGbb2PaW0Y28Wdw
u2qpa6lU6iyki63txJPcWFsvKBJzsJfQxdyq46bUFrZKY7opuJgN71xAQaDgOaV6
PTiZcSAL8BxkWa4dX4Vsp5/f2pmcJC08iMb11dVC/xpz1u9aVTiC3AXbSx6sufRr
CNabdi3dN+gQl6LpS9cydavkx2QOQZemuVZ8GgN8vEoGkA1d5bOBSw2/8QtWKpEC
YiQWBdv2Vaxi8PpXU8FEa7Z3g9LovnyJX9SfBjD3CJ1DxCJZzPJwS1LflHwXAGMW
AgYbxX/h4xbLjDLe7jpvNir//lsBp8nj/fiR3Iaf8CV+WGxC/vpQt1+bIYo58Aul
G95wjyl/TgL+6wq6nOB8Kc0ezUtWQNJ1nrm6eu894y7jlqcqr4bSe5oMF5QdgSey
+ZxBUlwBGkKT7P53wh/oj40pW+AWDKmuRdkYwYsViQniKdfefspA1dXKKeUzJFp9
GqZ2DUigPhnp9i3Ppz5n+nefcxt1vJbWnE1g+LeazZHwWcLy9ws2WsQjz5iQUfS/
qKzDKUdOwxyTeX8kq5Or2/ZTPs3dbFk2txpw8Et1rcn6rUIfbEQVlaDJTJ+Y9ej2
yYo0kJQfP45BA8ygMWY6iEcZUr8wyGxeb1ianPd5phSZB6oRtR67UVFOdZPtqPm7
qy1DaHp6JsTNW8Eu1lrGzOKY7GvtrFoBzLZZIcQiyBls/Y/rKcPjdr9XcacnIsSd
IGaNdea0HvQ+d169urrIj/8HMynkn3faO0qLVquxDlYyP+4UmeJnoM9VW/2k1HV1
hQh3PvTmLVoQgJzLFbmAUt4zaEvSdxcMPjVw3E/vC/+m6Z24oCfg9XdGr9jzxqkg
adgy37EONmBGc2UZOJ23xA1xsKbZjP//3qlm37Mzk5ra1aXefhTpVqdHdlth2Rng
YHoBW2G98g9exNVV9q60nPqvULlWG/8EyKp7ddsCXEQHJfICG+Y/cQBT0f4pzgs+
PSADIumIv9225zBB17RiPhI8XUlrHLvSh389OwIFNj97b6A/T+SYIyAQeRuHMY2T
WYm0pM/rvzzNDtcA7XsLZmQPmD/AywspCUqUHKlpKJy8DLnQeDLHU0hiNTGrrrQN
l+VP/wnnXU9btTDtmlwTEozNiZEeKtARsYUbAZzlT6ET7LTlhSh2+LEW6qPey9TZ
vLE0vGcJqoBxy/eycbdKtz0WwZbGpZTknOmw1ah47TC7N/+OMgSvR2nH9JuuxWG4
DqkqM2DwJkm5woofZe1z5LVVLD1r2noQ0QbjnaS1ZwDYHb448zoe5aNJLFBOO0Ta
D9+GbywQ4p2uFVYS9iW5uOwKl6JHSZjnyDaYEnFB2tVNqwAcc061pmbMKbMbXxAO
8L9B35VZaBYxpJWAvTLiO1Tn8chLfquOFZp3JZ7nUjndR10+lQtFoyzqiDlHuajV
iW2JeyImJKJr3G7HGCh9KEDb0SqEihX/4vfQHatdenSKKOHeOLc/uRO/Cahzwjnk
WZbHv4ErcPFgLCRO/JziXBY8OwezfDjL3j+LSfIBnPOn3SJ498V2JxRaP35jHmmy
XX6DQ/wuYguiuhskuJIXeFGe377wySv6H04jOncvv0wj7kUb8rJwD+sF4qTI35IS
B5lgEimls5/NSraAjd7u7rHA+fOLzZGhxyGy9HtxP+GtITWePd1jKrqRykcc1D/m
Wp1DPldUZ+dy2xz3lkQ4r6I1j95WbEyc/5nl/cNB9vK14iS0kEr12/bKCb4DNdYW
1dtwcPXsdbTh+Tcz8RaOBZd67vzHx6lc41w41eI/5jiPNOwU+q2zJ6YMxcTgE+I7
iNwiOafzhHj2ZhfV5xqa6IYZromkjch1PPE+NEimZC62eDuDkt6t11zQRTBAZj2C
xCmvQKRLAINRHFynxPnCO8xLNFkkkpmhB9eDbC5OXVYCk6k+aRyTcploqrRzhrjo
rRF5mARJGByq3g8QZYFnxB7jPgtEz1AMCEJvrlUK1fkOEfAKxxBfDUjcB0szAy4F
YrdRbI69CpGWnNStL8TiO0/MDy9n1XXgKcCGGZJnh1yz0hgj1tF0vSEYGxTqazBo
DV+zuZUN/vIPfK09KZIW5518SslCLm7Fd0wX+9o4Q+q3EWbvBrvEE/VitTMpQauf
expPhtipD/XA3Avn7VyxxHNpIwok6AKCy9Oy9BlrizSfrRjAJjaxWJqJt0zepm1c
Mwiyd3oAiZU8iReuJXqzFagQZdsEIjKelVWwnBuSxjUn7J7AxUz3HcSjaOHQGIP1
ELDTYbsJOI3efvO1wMzu3HEVqyXl8avQeBvqLbOp9y0ZsnLTGkhIYCXW+HJQTf+u
2W/GoKCGfNIc3txlB3O3DKEqo8z9G/wXAWX/oZJmoru6Pmt58YPoRscRbI/+Zdj+
gQ/wfF6R5zpkQ/QZdA89+PvPNTFlz2kGg1zjuhDG0C0fSjy6Yu2EzJTryX6Njs+C
wk/FP4FuU3GBaJ6yivmhyjs53xroNNhrJLDgDUnzeEBkrx/2lYkAZOcFdh8ZjVND
1Il5EKORsxJQ1cU9YCzD9bwNtYAYYo2RgfCnWK99LdnHyBlCRJlR1rOrtMxZLgBq
InOiFhuzznM6fl522n2Fpj6wzd3M3h0unow70oj7S0xR0UYaTWHH6qO1JFv7B4OT
gSKzZbgjdbs97k8prFW52+SJ3SjAHWrEzSvbpuWvKPSpOP9uqlgywYMUtp1xBTlg
ETbCBcV4HfyJNxFyjZRtU8SEJ5wU9noj8qZ2zP37om1wImW50N45K5a/UlLuj1sr
wkOQR3Gwu28oJFR8t0AcnRSmNPEM4LC+pdCcHLeGMnldlI0Y2eAUgb7w6C1STnaI
+K0CTa0wMw9ZNuP31iZQNhuZVXQJxQNE8nHmxchUfpsDqtORvcR+rvEeop+411Ie
HSHIcf8Fk48KsAD/R7k4vBqMAlyMsUGhxiZazo8nAMckD1Qv/B7h9dSiIwqmXs2D
9AWcAksMD5PBO8yIpQWG2ObRQCYvfCvyYlI12DCNxPfmfDPrQmYZNN6cw4yoOzpn
0BUSvAWvTbZticpWg66JqB+qj12c30uIGUq0SqMJXPW/DMN85ysM3Ol7wJoknnZk
6XJb2P4eZ9pQU5D9pdakahPtuD+D4vJgQE1EEWpUl6PEMZqeiaa9ow+hF/OT+eTJ
bt+rw0jFzLICVFB0RdChv5bQlyp31ryx5/m94u1dzucbgnb0LGIVY5o5w0lgBomH
IeVXydBvAz4F8x8N054iFKioanwAZdz92OXl3zSyFM2kr5wdotBcJiEzDFmaIdaA
LMc2E2g9yLx/Uq7WQtM60BQoMOkvQ/oFmcLSHg+ntH8skIphKi7BXPwbEnviDQTP
cfaQUZAUj3xY/0qvpWjsVP13UNaCva7n8FgLCeNnPF3zrrQJCkNwSTyiTFA9Mh46
Qr9KOUTbEEsoKOuzZGqaoxCF3O2dAijFQf1AbIpOaMn2NzsN4Iz/ovBRDzrJsYyI
0zsF+lxCaHh9MjtjqUaWlZ22Jhqh6DEWxa0qzP/E3gYHOGsMj7TjeDb72fqJkvWI
IgI3+/QqEV1IWOpjwRnkm3QfY808bSttQhf1JDE70NBz8g4L/UgbO9FAtdh4GiHH
ImyCAPug9BHfzRf/BZjqVoFB9S5BB5A9uXWd1ibwJBtZXTRbXCxHY7EJ/bp898Bk
YFttlzRBCX7KAMlr8HUmbdLf+u2HRQ/9C5SmYkm2woKI9UBgNspPcDZPqStWX+Kj
vMSazQtD4/j/NGyIhvymubu2+yJPoVn7O66LXqkZAAqXfk1WfhAp59RxnaobzLnK
ZADXNLNaerRnrlH10WNcRqnlO0Q9jbsDCr4EuCkrlfxB25B1MAo+qCYqa9iLiBcP
MwLpdiXhmgewjCu+NVAzEEpMxG4GgucmWZfQJlQL3I7e0U3liyyEjx78KatxmAeA
/aFc6vqMkFugIG0jmAHJZN+5S8UNDbHozjUzflS78l9VR99IYZkXs5IilJCWkfxV
QwE60GKYqLqi4VoplqvcACycBT5xYP8/RzKGzIVPbIWyGSXlWArB9QWdg/as1/Pd
ykgrZSsr0fq9oDMgiv722mrifK0IxNsg5JWtP1IvkEz35hMektpVwsc1GZFToFAo
QPGBV894Kxj66TuQgItW6dW5sS69Zhk8e+F3y+Whrwac2Zu6zUuCCz9KD+UwHGn9
VpmaHfnkbn/RomP81VJMq1lybduXBJRn/auzw0MgLXRufhBxqcZ0JMV8JpAQJOhW
GUo30B3TVM4xwLaBizflswuSbHZC9O0QSq3l3BtIVyRjQeqP+AEnzxgo2uW5hSaM
8nZnXNsIvdkbKM8o1m2OR2JP7fxjumBp+B/pBcJRn36qeyWAxgdDB0RTblzjYuac
BMQJCkUfrNN5moN/fcwRNokS+Gh/RSaKA/jBUucC6zgQ3GwGpCJhLXxb1DJthluQ
NtfirWfRKQF2HZLcpuhHy0VaIvvSElWRQ+Q7Fh01/YaUPKGrO/QBwfAyNiSEHGUX
xrbsX8FNn282W02elOALbOFjEZne4lDb///ym39Rrrv4LKrl0WWCE+WDhCv17Ke5
DKsx1e78lWNVSZJdydSjYvVntp/cpflpwNGmsrXPAm4EJ9IBkIbyXSaoy8bgCBgo
rVLEMQ8LvTSViBwjLJHHGVd0ehmgSXKhWRaigMtV+lf+ytIQtD3aQzjv8RAEuCCl
6fANROW1QC58a1qyntQYC+1THxWwaIGKgqxTCUPuERj+p2OIbSKVpTHnrZRJyuNK
U/cWWkjgc5E4373tss67yWzP3Hw7t6giUBmqwRVh5sY2ll1YtNK8x3lOmRB3UchJ
pe3+sdXYVmLpidyy8rEUHCBSqGQFR1Qt9MQkMA/PW4jH1vygVNr9zb+tEMApFDAG
7SBdlwXCBnBRij7yTRByHd9CBnFs859g7KDgAtsg2LyFe7OcrPxqGu1/inkpon8k
eprRFm7vyt5q380ZlHVVHLqKQOVOQAinUUH+aLLJBeh268YB0cIo9oHtfPoFoGuo
NdEV6n465yS7VRa24Xibxw02ncmutQPq7znHaHUEiagBI4uJD/v/uUTynDrgC5k8
YkUKGA6wGbdKIKmB6NR3snV0JjFRkPU1OwR7EoyHKTxfkfDNbc8dZsoKnz2f01L8
47gxHY/f7VvowSmtjMSO8ojx3XgZKVdMLO4t7mVVpCcNmoMLnJqnL0dwzGcLqYfe
orOvUriaU6HgEqLaD5vKwPlcqp3T99Wl71uFtp31eyXOOUKXgYzNii3yeiORUnXj
O7i/SfRtTrvGbL4ewo6s8XP27WHNHUpIIyD7M2Y1n4XB0TAomLIzdk2YNn2FdIVR
xagOkXzvHX+Ieh+NDiyY9NWlhge9H60ShvPxxEUEp/2wakNEM7MJ6j4/0qE7nPss
HUHpm9sTCZKdaNxBKVhBVeMCp3xsvJ1xRoFNamYLTQXWjVBj5BdWa073dVwp/8G1
Rog1hBf7PDOo1lgaJ6aHdWdoSR2BdGcUFyLpgezpjKvmoAhpUm4ylDjfwYYVMgJY
UoFbggFspO8oVhHEFG5xKSpIrYHUZhEGajVCCdG91I0lEBuPE2ezL0U4aGHHmJxb
YcN8h2kkma3MPZROg3g4mbQuvBgUGjG6jgCt33oHwmwtyhBmI1y42qzNo+NeXHx/
e58aN21efgHVhUrlAqXdW9qY9EA73hsLFz6gD/Egeq1N+KpSETiq0bDHixOgC7DF
giRYmfm4STtFrr51Gdx5SWxVN+DDz/l295S8IifZTIljNNF8BSGWMRHgRU2mk47W
+SVHAqmIco3YXd7ursAC57YP25SGiiHpW/eUX1jGh9COgOBtkO3IdItSCT8DbdZY
8JZPVpdAqK13GPtHiN12thL5CLWWR4Y+GzHbtzXvaC5AdYSWiLUWA8lqwYbV2YP4
RSx0eg/+68WwhBEmGIPGBUDTTUyKXrz98WUQAxd6BaeFcLweGOOstPmPtsZNZEuB
Zr/EkWbNvE2ydJLEiT0BGJ4kttBQgPXfXi97fJ1Z1G9QoKIF1GLcIRPZlo9unDlG
jlQkSXCcmE5T7MxboC0vh6U//0l6Kut2/IcOGaz9IBHGa/Hy0orcTjs0njuOU7li
lgq1iN+bPMR5bGWBPWksCwvJAuiOMbo0dXEzK2uCq5R9iNNGgrnukQh5tMHZAKod
KacD2THuqTsNwQ5QF/hkDeISlDmaPzX66ra83/JVzP1ajVbSlIm4hyIw8mhkUaLB
C18DvPTOVNs9ENC+WFHslqdREZy/L6nxAE1pMWZrWlvBGKsKG7qUTZJal/I7wqtj
hCkMgFWtA9g5GU1Oxe2Cai3fG6Nqt72eyxbxNmqULQxb74pGTFLcNw1L/TVp3KSn
jCDhWz+/qMGoBoYgWrWewnnaM/EYNMp0MzCmACfT9SzVawk1oEj3fJBhcxgurXq8
pMwMRXUI1n6AAlrCa44Sa6nJFud6USbuL4My98+GfXs4gg4oEsJnPGH18O35NA3H
g5kzgaC/rrTCqubJ25MNP1AcLtGRqYLEEpeNRetKBiGVdmTZd/AVxvzzVhLeyaCQ
9519zG181DrkQu26AURumATEeXVpEgvyAvkGfC92JiSBiumjoiGXN6pV6XnVMPOE
XnH7WlyzXOgGfFEGEa6+ss4E8eZoUiG1vYtOJiShZnX8qrSKAhPIpTtLf5d0XS1T
q97hpdwHqSLOwaGIjiPswrFfRMEkeVyASj46mF3QAQ+ccuSgAbLMayxuHK3TVugA
5K0nM0r3XT5HPWk7UEK131fdgEnDKfkXr+gWbA2Ziy5iihVwHwEzrVbSdbyU+xJh
x3k2RIIEQueL7lyNYc9pA5xue5g3a8h+DzIC3/Mvoty0h9W2AqYEFMLwGGUhK+u8
MTiHsWmP+Iinx881Dzz/VvmX6eXZy9X3IjKh63lNjq61uINpaQMzRLh+FDalSgqB
YhHi/chsKl42wA38weEGPU4VWNVM2V7mkcIRLzyZC0LDFC68xK8NgRJ+ByzfQQw1
d0Vhh8F0hiRBqfwc1pzDMbIRp0LeaWkJW3cji9WyLTFrdZ4ej7zteGtSa3AvZ9xQ
y3YFnuuJhBH/o4Qteo/rfM937FLqT2ycc4mtBlhDhRYf1bLzL1oXO53/ZdQXsg3F
uzva8kVRhzAV12L2LI49N9C/nuCtIxGUiEgNVSBBF5oNeW9+BNep2u9XEff5AWmj
TXqNA6/hCbRU/8I7gmnZm+A1v2wM0KJqwemNWxYVY195F9qa6ay3DC9NaJe/RiCx
3wiLiVsugL5bL4hm7FawJhb67BQaVMfy6Fzo93yUy6p2bpDjU4+SLtBpLTLMe2Fy
5WHHTroiLYjFE7xrYV3/Nnp3FoEqezlPRqjkM3DHuUEXMkSTqOl6CzMy+uanKHL4
JkO0P//sOSByvmL1eO9vvhtuniabFWFojOp3sgFv7yF6QNeUlu1fjw3YkYVp4uxZ
JnO5YYTUfxY0RNGlXCB2f3R3sE/n/Y8wx93o9fbs1g8g1iiF9cdUV3KxI0xkRaQy
8dqJkKzxAZXEH/cOwoJgnRyhlgH4bEpRn7DbNVcqQ3AiDcoqvueKoXjtz+o3DVyB
tmAmk8BGa/kZ3g7A6mSaWG7C7WgWRV3iebc9PmBqJay6phFIJCKEgBOjvbAa+Tq2
S6XdZocRRsdEPf9yWUbc06Q8j19LvkjqNCCot4A0HrdQcck5PNO7X8thKamoZBIF
LcWNFyX5CikkZ0Lcyo7pVCNcFwR9NrXWj78tR15F7txxR4rG7aUfm6XtgHeHRc2t
nUzh6mp29dAsNwlj4ZdgG+5o0JZvzHUDQca753lTUds+CscT6D5GTNRaYuk6layS
LI31TJ/ictpcd+/wvl2vrcBjWrHxIMWarLjxpIPJ6soIMQq61HFC8VUjM4+0Xu3q
fwbtKJ9v6rqPT9KheAKzvOLC7SFqT7pcNYN5wkYmHDOXNoKq7WETQvk367eb+K4m
xNw3sVeKEaGDTdULGMJxGAv//zIVPJEQdwxWoSH/Em/XaOoS+OXue89d4gec5WRs
9mDoHDkmcU4DovsxHNG9ptGHs3Wn4b4JPaU+1D81mtRHxxXpSkie9lKsreMStPrD
fbNf4jZrS9FNPfogiRWBbAI0L9fkawudq/YOVNllMvvqiHte9hKUEqyXWJkVreDP
CzjBJXHn/xfNsY+S63oEpJ0XeHzUsPrDJd6F5wy2T63LnWlWkHJ3KV6/Ah+ITPig
mO9wFeAWlPnAQ/YgFp60L2AwoM9ueyWKj5eGIUqZNBmsgZ6NuyLKockku5SiRQtH
DCwanHCOFNIOPvLrszSEIJAyuJGMLLk9Ms2jdCJM3J1hsd311Gd9LIgwiLO/iVF6
IM0/qvAff0fKQkV8r/3GdQx1HEJT1r58ZJsmbXsjWbqgrcnfgs69xf18EZM8dKTj
4wgSllmnali89cDNv7KvAx06kxx7lpRTvTVd0s4Z4vmHRlne4e7xowfz7APXjE3R
LBEvyZMYtyycecnGIxLAkmqWE+nMARFJQVc3bGBWEacGuhJoq1P56o9Jg1DiTBWF
B1IKJRbznEkpTw+szQ1dduYAKkboUe+Jm4Iohol4xb84vMEYLjHxQ780zr+4jL5a
Nlxmlo1LUPGvsljwKCmYTn4ZaXzvBOymEYwcBv/jEhxPd/HIjBuQ6WBPSFvTxQaL
p92CfdwA4KHBRn89R8HSU8qbO87Ng/aoefA8/Up5JaIOxQ6dAKdYXSeMerNPPF2C
Kbxc0pGgq3G8lu0axgtNCVdEbO4eeX7GQTOOrs4/kikWtUbZdAzgITQj06NB3eqy
bgRCjUJwfXChLTisROLVM8hovgQsfMX15ichd+4MDFyHmbSNONX6BGR2vTmupxVH
vv59m5cxFi5I1wM4CDKngqTz/+RJkVD0Lokg5wf5XxxSs/I2CFZe9oFzALVBKzjS
Lxm8uPL46iyp4FT/9rWqgZjYTdkgEfOFz2txmfYWIW6/7NCQPRmDKJcmcrLyL2Lr
hWicmo5nUZ2ns4F9u3OJTNMhynyl5eT6Bbhliuc+D8B1zLCZpO0zqRUK1S2eZ6Xu
NmCkSabuoPMtAxvzuTq7YotDPhrdKHWVTT+Ub2qDMkCzpuRIEtfvj43+nGXxIOCC
selIHlGZPYGCHpif6j6W/TnlYUsMtTKLqtZPqahrHnKMct0upX3uWFzTChMwNlEQ
auwRxeAxuFDix6mFaNYGfAIcidnIk0SshLxogGo3CyVkezrKphThcC1xaedGWvy+
bJXewI4VQG7urUypbtkvb5PLg0H4tNFGDuRrOyVH+eJe6Tjp1VPhoKsYrNw8C8dO
QV9Kxms/koeWr4sVi9SO/GUOWpIpsRyeX30kGT/w/XfGItbS0LgR7atrNECQTCXn
Tb2uNWgHQRWzo+e0qeLeiMkM3LVdIsV9kWl9OdjRtLheTjuyboGR2TSeZgAk/j2C
`protect end_protected