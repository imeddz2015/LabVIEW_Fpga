`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 6592 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/59UwEX+aE7FohaWu0/8IpTj7mav863zUNIsgIH2BWb
Abd9opeuBjbGF/waQMI2vMJTwD1ie1YueHc3nSNpEh4OXp8P5ybZFY89uyGz3ztU
W1EsuUnchJoQgbHZ/sLbgtGRgsrAFn+ZoIeGN1d6RAF2wAESJmYP8zw+p00RvjZ5
JxSuSZo4cTLBl0ln+ZbwaXcGNxJnunCqKol9j3geNsIqSpjYWROfheOIYwpGk6MW
Ya0lbm9t/MHwMkxMIe5qnADLvanH0RctUHQ9h0UDPRJzffk8rtTbRVKKuUDfybw0
UMJtGk+CUs4ZwAsqzVwS4Bn2pXEAESLyORl+VWnKsNlCpuGk7Vi7MJ5jiJd9BLFa
ugDzP6QaGDRN9UpmNzTHbeUz5HE1zyxpX7EHXG6FhuXtsnZlOBS8Se4+TFStwqXM
aHg/XI1xS6Iop+3gus9o/KHSXtiAsuXy7Bq5h6v4JO8pWgRUHYK8MP0Baptwh7u1
w3yWC5TuPSWDZ/A+nxTDnoeHZ3mfiJpeBLHsS3vshwjPJBqjV/1xdD0Lnuo8RAIz
qH/l/3/82KvpYj7mfHmll7Z2Hyy9EoUtRaYPOKY3UlPHw72fs/TmF4i4W7HkUelZ
oySjnWT48nO5G+TBXG2YEAu/irPN30EAQfAHlcXYw1oeUhoTPBrJFeyxcOibF4L8
btgwHxuP6BG4rUmlSNxYzPe0iC2tUpRgJhgXp61YRfnWjJcI0RMdvNCYq7kRtR36
97m6CCBFpvTW6GKA2+rO567ttQsNS7k3CUiPMFDPpd280sQ5WfI4s+PvuxnfX4XU
06QIJO++tCOUYs09cduYIprykz4cLEBZPBnyxps+BCkpPX04AnYImht3b2z3fOI/
oTEijrVhWdJF8xZ2LA0ameQZpIbwdNvwC0mj1kdskDfNG1asjMLTnb6suQ8oqZa2
OjMrjztEkJTanpkvtU/f4K7PvXYLjPpLsv3GQNX9qwfpFNv52s5kHD/OUQyqtc6R
Obv69MVgsoUMq9DZZERt/5p7sYE+4hbMvPw7YNBMAZNYrq2/lecaKKikk22gQYkP
GdwuaH4pECqZrsxQ1IfNNZYJZfc4kfY7MXgph09636HsexXJ9R2xTRoTI/ggvzxb
Lu63B92xkPDrfxCxzdBuIIFY1PRKIx5N3jGRDl1ARh7BaePwoSnh/YUtQgTdKZ1N
aw2j8DyChytHQBXgPj6Tqe2eoVysd9CjizUgjQQ5KE0RVL5+cb9D3nIMMzU0XyCx
azvgiqXycJH3Cjqb99bgADT7vgSVB8Ylf/Cwvy7Bhvoq0sqb1mBrrTPjRzq9ORPZ
YkBLmiwo0WR8c2ZKgu1ZydgfHXpSRlxKzEchK95jJB0KjoPXGuYIVHhKKvxCYaX4
OpBrflJpkIl71JYzguNqvOekmp8ZQ4p59sDYXZjYH8wVxyNyCjztB/9DfraXTmIN
TboQuThVVS8YrdFZBeluhqV/SWVZ3du0g/dXD1l/wZkyI0Xuzx0IoaM9UW8J87gA
cttWiEAF59ahRA47ecdEXC62lvh795nccO69czh1YzEPoDyLLGS7i27KJXE6kU4j
1Nm0lmj+lSyIjG52K+nhSnrp0Vp/5R72k0GciFR26wphuq/WkjLV1SnhwPUmNQEb
GcFt+N4UE5Hxg+OosCcXtSf7OSIo/agkBQFioZGiUvs9w5p2bDdChCs3jr+MudMh
oOrwvjPzGsyRg3/gQJg76IUz4FZNHY3B8djem+aHbWLfgppp8oQh62hWkZv0iWtz
gXXRK1GwX0ZUjL1+D0ivM77qs0FR161DzJkkg+6hQ3CHTq1/7zP8JN6eS/Oimz2O
WJL12bFNcUMAWsHgWz9CYc6dZCsFx1+zMdmgI/1TVIuKxp7XG9KThDjY2CF0700r
9yGK1T7lc6VxSIR7aIEfkMvAn5oZ4ns7yRz2gNj3bsh1GzvaZJSRprhe8ci/DKFJ
27Y9OIv/TqwPNjUZ0WWHRqPhK+ospqRYG+l37W8sf9Il3x56oq7FaD8HYQtKSeHE
hyVQrMs/ORNbZIyuscaKbJZSgQVlxttX8aAQejJhbyEVhVRwCF+5Yh3ATJkZzRXw
SlBy8d9wDqjwxzYd6q47I5cIqz2Uc7S0XYLPywJ2T15KZDA5kIAXdux1RFzpwGiG
a1q9Vdun6mptM08tOq6fXyOZr/2NPdf/UJ7/KooEJZV1nsopwCbEIWw9Oo8dixHG
FwwxKKWy4Wk053NTFNNmDUSI6Sn7whpAw4+inbiw1e1zaPFrDG0K5v8SZgoT8p21
d4grQZpo8ZgekVnz13Dus34sUZAZvJiu0lPLof5ScaMsIg9fa14ObarIhXgeEpnN
j9Q0JPmrCVtzWymTt7DAnsLtcRxtZvdYkoR+WnpNx/HZUBOmMdjHNOogSCDzlkWj
adf2gObJ+2F1Mz911L0g95pwXsVjPjVoA2DJYpOhLgiEC1ySdMR1/xqXdBP3PvYC
DHwjBXLexNo06wC5+e+qXYQrSY46FyEWjKmMRLh2G5W9KnHg5sv2eS6u4Jo/qul9
BLlD68wXjVU8WgSfQStk1IV+RA37C9OpH+Y5oYp5bIaQ3XPhmCEWBdYYmOaHfHyx
o+Z4IiFOGUNKeqagtK0xep2sZ8zJUBRKC1HjBabFI+YxGXstrGPFMc1Qs7Ge2bL7
Qg73eDSokwnmkQd0rCXHZND6ZBGqp0CV5+soqQcmnaUJcJRBLXzLNLHRXb4uW1Zi
PFaZbFbCmADkunRMeHct9cY96sYG1jESdoYZ1K42rcKA8llqxl7iM1mPuQLYM4wz
Cqu/cxYDVfMWZBV4TfS/lezkiejk/uO1DcHgeMTPTvHJeis1UGWF0tSpWJCMEG0p
lZL2ICdd/S5FP31q9DehiHbEEkkNSJwqWZBVF9KMTdbnsd6QKhK6MAQg9DrbMwV+
wa9/CIRxhvLuwtVOO0cm+MC1BXlOHgHHNqBuUfOJM5FeMU9Rb3svcQbT9BJzT7ih
E5wSgB551A6HoMoZZ2JZnm9Ve7ybKkYeNEx830Lv3+5FQMz4Djb79+u3ZXwxaDOp
uOWKIOtoARR0CtYTZKgc5unLoka6gwW8F/x0Aok6NmXUWHxwHxAyzFaubZrkt7Gd
YzI3gFDzwbbVpY940JmwHnEXtb9Voh/UoLNdBeADK5/n5snKeYRxdmTotXqyHo91
/EwBSHaCx/GChpmzOuejGJTzuzEN8fhI2PSFyF05xbrcHWpu/f1V/z8h6RwJiWFZ
mn7nBHOmyMPRQA7pBpN+FDRAztGsxmFL8N8y3t0YO5tptMdn18eyYEXBsEena+ii
O0vb8U5IOxfqzk690iVfOBbNv2N6NI/i8zBPUip8jzstIHZ4mtZWg3tWfThlbqdG
0VCu/JWQm5AwtYoiorqG9c3/fW9Rs6XW/twAjF611YvFDzogllJBoUDPKh2z6cY4
pOlW82rnL/tqCxQM2tWvDo766f2h87mNFHUuj/w/ka2TGthxYjJhOid4a4AP48+I
r31RJuCFIeBuksJ7hvv2OxStkxUzSw5RJzTmqwR2CpKvYC2jrHMc7B9Z612yWfsY
iovK4+a0XirWiL33n7GrzYOHSW6WFYENHKt7u2n2byiWYimXnRaSu12gYuAZ3WbJ
Ls7KfD392ffT6eK3BCw5OPq4mE6s+CQF0c60CA0yO8wX845NC6uU9I8GEuEiW6uW
A67Mgf+NLRdKWsARBGo9+4z65umI0L5eyz/ltJfvQ2NFgdX+9X9uWJXuHT4OoyDL
TMsJ6IBs3CuGtVpmwRa3L+xf9Yz5w/MRxIBt9YLcvjsXg+YFKBWItMYy5kPbzxbO
ppF5wa7TPKk/z0s3n5mJtbrfuuQDARHm0YI7pwX5ebzWk4z/za9i/Y0mO/WGW31M
3mgwNL31jMd5bg+c2FSMwSnQQV2q9yn5orJ5PeZB7yN85WN22SsMiGTEKifbHsFZ
MEBqMEtGlQ48mvaf42C9zITW2FKraO2o3YKO/hRBVa4BMWhMWPsLfJaz0ySvvKom
JiPaXhEav26QW/U5/ddgubi3ERAFDgx4BeBc3vjLcC3Hnkishje/9ZSMwk19Qqvv
CqUmvgNK885p89aK+weof9dU3hGpgr27MeaKouGpTyvkSxCYH8IpjnBU/Fv2iAD0
85worQfH2iIuyzVK0I8MPMA7x1cQYJiNBafz/VHc2JgAPloCnuwAFnTFs1ogB/cc
jHKh1ydYnImCp8GYKX9Tzlv4JPURTaJsDO5pB9XH1dRZR60b9kJTLdeQgTBbIGx3
oFaXPtwnImTVDQKUHb9sQ+7gwyuw9TnOZS5y8xJ4l7UTS2UtmhID6P2YXDDVGE6F
tySCKTAdQ0YwCiyV21JfChb3i+hbJq5F6gnvAYtzC/uXSwwEnNRPkPASqX3BcAfN
9/1lW6FYV2krTlRUkMSbkV8p1tpcn5B5HrHqKppsXZs8jP3LlI7lgy76umg4mJYK
63k2f97l6xAX3Scc8IfT0ZNkQEdl2OxlQchmW6ig5MRoo+fc99KCuiGi82duEEXk
f+pBluhabf+8hNZqjX1phYg05USIPGwWKXvG6nQrTiSeWQh5opmlrk2+HScvy8f4
5ARfPLVYZ45pAmMfjePoZEHyKyQiTAlaV7Onx1qFf5c/XIhGwyLeQ+ndW1V+uDBi
lrbpcUe5PLXa1JcsGOU0ruB85T+WipIHZ5+QZGxQ6fb9yYCa5x9x/a54kHPCGxU3
LG9gFWvasUZwys6oBjplHXPrJkoyzGtxZiEbNJyQN4ayvojUwlVo7VwN5MVh3Og9
KVU6CMkPEQCVrMpjbch+D5lfzms9fmL6HfHPChlQLXTt5Ke6489zz51aMSiCA5ul
wh6/r/hQ+PzwPTIRwookV4eCIOxN67i7EzrlFdwj9qX5//T+NDtuXQn2Lta0vxWS
iriFHKeZIifPvMCUgiNrLydGYoeZcI/4F2X6rlAbWGPM0GpWoI0YPXU9CDWNgZ1s
0xN4deMUm7W2L7OIwWFqBGwhsBls7Xgea1d3MGpeDkQ8L+wNM4HCrAmzHPEHqeYL
EGCjcVKAvuAllaYBPwPgtT6TnxD4mZEAPXhz0MO8+SJuE4V6OdIEdM3CFUWr8h4w
1s1UkuRpCTcH87lXC8ej+dAD/QlkelRqB6E1kqEEpq3g2BeS7EN38wXSLpbnDe9d
cxsHvPfzRPcWfTX9+7CAigGyoSfTx0oDTcNwQWyzYdSEc3UWIBMMK4aIrePm8B9w
q6DsQacPUA02t8Z1V3uF2Xsq4C7Pix+WtzS19f4T+6Fho72pASj9R8LKwmBc37kw
dq9L+kxVBXkz+1xipU7+WPMmSB3KZe0Ph7Zhm+emw9aoi0LaUWHeMzq4ps0gQMAx
LUir3efuY9j7TRdDx4PTwS66ia7YQVMilCEHeP6LM5r1p2PqyfHQgPrXMbhJdSeC
Qus5BrHI6ydFL/WAq447wFJOI2IL7ux8uKoPBuzULB3vtI/00YWVZ82Pn3GB9zhh
g/KnxIpkCMJ4EKs+MbRFDFldPfujuxYjLkY0SwLlxDP5/hvKqwjWqQB+EgFdwdSM
xihjtFI3iq3U9WERxVafV7gQtj5RIZMZGw+YTIQJ7Lj+ubEa0ayDUR6ART9vLTO0
M2H7CeOHha1nOUwEDejTR8ATF2H7mD6xeKe/l5c6+3WWLvy+MjZkIjCwPz8oZi7h
1cVaEoUOmvbn/KTD6R8mot1FedDlh+sPHSxWBt4HuGscIO1mmxvX9PJuBcbdaRjF
17Q3fsRpWJYvB31Kycox+WEKXTHxy5Ke3YcMyHfh4tBINrxTeR0BzOGTDp5Dr0Tb
EDZ9wGA6ppv9njlD7krVBQlJZoZXe0G0Aj0Mx6LeLjQsyev/8lykXwfU8NRU8O10
WiBqqHfc9Ihjo2XKQu17gEcz1SjuoYj+HXUcXfqHzFuhR52PkKfieQTQ6qhBU8pp
3lYgNEVAzZK6VUeWd14gs2r+klHAdiYc7ul/e87oMMi/taurI0HUO45K/SXM9/Pc
sYQxTXQXsjDitFVY53MO7Rlztmcf7mpLac0Ew4u6z4MGddK0+rdKc2DsrFdd58LI
nrT/Omsc4Pi/Y+Bp4aLr2SM+ce1v5xynv1skt2uF9x16sYDyoQ0/TpGMcM2DRt/e
rfqwISHY+Bujy6HVz5PoWTvbM5OcSq17eMrL3+6jaRTIJtbub3a/GQv1N/rUdH7n
SA6hy8JujwQwMwcN6asz76rIobaKeyO/XXAZ2sx31NeJcGwqxv2OhT3Vy8nOKjmu
TBFLJjSZGgMtiyCaj/pHxn5fGDf1ePgqkp8DaFvdw+p9P+Rk9HIQlSo37WbzQynY
Jn//ws12kL09j+uKem4n70JaDPVeKZyw9UD2V6LcA8XfPbjrH3r2d4mhtEwa1ORb
vULTZts6xPMOPE8w//CPKrGLECYyhz/rWCbHY8ir+x/Dmc4WxYiy5I4QSaG7E88v
KxJqXukLg30HWiZFBCJIIDVCQDg2+RUwvRbsvzsNpDfK3VP/nieyZs4JNrV8vFjT
xPH2zuYVLgUnGQk3mWnOQD1fgAEGv9MFNahXnDdTxXl/hIBWPLld5pA3C3ZnYogB
pM6Lx3MFhZZKzHrCb8lTQcUH2qj8cGYrrGMreRhloFWUURygn7IOZECovUaupALi
ISX44eoDQPmdHgT5d25rfyYLda08n1Tvcy6KgsnVVn4jLpRJB3KZANaUyCFN6HNg
VYOWmbusB4mo2cDimu78dJh61QT4D2HuERfcKAr9GMon3w+Zs+MotehcqKuRVbP+
zFvDnaXNOPY1a0Qfm7zQTHtcaCQ+NP6ZTRrjXIKX7P97tRs9ADTKmyXmTHJRIk2V
UAyYZVufOCJ+4LeP0s0t5Fq16jh1r6+rWWDNhYnWCNr9NNq6wkdApCJeRZF832JH
56HURduoRSl5QuMRm8xEUcgRAVfc7+1HSvPsvqMUsE2XRIHoRbkm9ttq/LkbhehJ
h+Huf+fhZ/EFz+Vxr6hNnec+WM8S707599wku1qrT35fhoDCG3Q81YMvnQFYeo1h
Y3aVl7U4k2ujbpKVCQHwBLAwCWLy4HRJOFChMLgQQxjduK11SqtC4KxUoG9nbf+O
F2CsRGMhj0LyWTH4trtyIf+y6e0Ng6apCM15S3oF/CBmqf1ZhLvC6HcuUrqaGR+U
10VeiZP1xor/vRDuqhgpgRsXh34vt2P/iP+alzTken3QC16CppxTBfATsa6SlKbY
my6RKXiYIKVEv7PtkmeKbzuyMTYD/kBnYebDuCIB7qUv/meWO35zxST+rNb8N2eV
MdCA4ud6cmoGVMkJ2Dm5bISoAhS0AzgOpD3umaTA4Vhytm4wZ7JzyDtD98CkBnkN
qoA7UKK5IYkEEtzmZBl92760pBJicOCXUpa1oq5npOqXEEto+kVkQRAIGBViJ7cC
sx1vb92uz/pZzEtjBFA38kwmM/P+ut0ZjNkGZ6c+lxr19vQyIio5OQpLxwtZMjIt
TTYruIZm0F88yKKg6Z7Lrz9Ltx0u8oQQ5Mc6poqtbigcOy7tVABNUJaMKZmHEy7n
g+ITnTksBZYJJsNP2oYAg1j8bH6Cpu5ScPrYZ+SBaPdHUmv+NXFE5zzLqbsjFWG2
1IP77uY2Cvt7fAfjeSch3Av/KqVWOSIY39MM5jsDXJYStpG7QLz/QidRh7Vj6nLa
THIpPepAZ3y9aJVCsQwh8Q6fU8eF3jGnB8mey4/rl004QzQ/oxnUpGjzYnHUcfYs
NvIWkdt3/UBMOnlB+g+YNL8BF+U5VgVDvUEKZbwVk5p03WBqPV0ZZgAoJreQd4Ww
fx4aGPO4vK7JwSXT/TfCDXPfUplin0RvKiqWpmLPwpE/RAwipTQqmy7M4wWXcRww
dDDetQt8tT7IESi+pl0Ki6VgknQiRbKs8nxSPHOMa2ZvwjGClSGtF8NYkSq9Cyxw
UuSAWTaFRKWP98HnRKmk2ApqOe7uokE7J6zzdtmbxLUpdU4znJu4GqsIpP2wnLbv
aQ6QbqQQvJ4FValHB4o6V+JIPVVDktwledEqtlwa0VIyco4yTJV7ECKOrepgpzgK
HJCmfdmLjjZBTICn6H7E5B3yM0MimqFP+Mdtu8FfcYo2K+YHk+TEpaQ6zLqBRnkz
gZyLpu0wGreqsZEBFhO4C4DZkMNxMrlGZ/hI404DSJcXPrTNSfziGF3cQHWzy8vB
sDax00K3bSdoUypFAwjq+yTZc9w/nm6KofqjXat4rjs6OnQBkFsnUgy7/mkqBpqF
/k1ugCkwQ5PQUkx03W9cL8TIA9MgE/DxG3fPB5+PC9x6BaDuU448IcCYlmfko+5V
q8hky9ZuZQ3RL1m40PrAmvRx1XIjRdIeQguAHNkB1w0LjeSzCyWXt2OBprZsJM+z
1hmexeNPSD+R2iyPj3NpyuUMzxozCqPd7K7ZhgWuq59Vo+bXq1sU1TEyOmOXEFPG
qxMgOPc1bdHz+j6stXHYNRuT/XzoN20eA0ainO3gpcBH6YhLdtlJV3b+X3jkiHCi
xHHLJi/leYam9we6iRKgBVrZdmnwS/PEtgLIAXAgB9YL1e5U78GxR8O0k5p4qD6D
nyYRCAM7GR9ZOuH2gThZn7UOxjRgKOD9sKMh9G94x54CuWk5a7HTzop3n8uZxexo
0RfNaiplD4M/NUalXKLBGfWCCh9orczMZYCdXYvNEo9uBKYbCn10GcR3p/Ll6BIa
1tol4vOdoSmyA6rIyTrfefe/rLNA6X1zbmTqdtPItEAWs4IczCdaAbdi5v6Ln5Dt
Z0bJTGd99WWl04FbjOl4fA==
`protect end_protected