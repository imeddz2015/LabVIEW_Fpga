`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 45792 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/59UwEX+aE7FohaWu0/8IpTj7mav863zUNIsgIH2BWb
Abd9opeuBjbGF/waQMI2vMJTwD1ie1YueHc3nSNpEh4OXp8P5ybZFY89uyGz3ztU
W1EsuUnchJoQgbHZ/sLbgtGRgsrAFn+ZoIeGN1d6RAF2wAESJmYP8zw+p00RvjZ5
G2ATm2jrAjm+J6bPpiDE30W15wqXnRr25t8XtV2KlSupsNXWXS4u8SIHjUvcCVqj
pUlSZf+hlUBrdNHsONXUdUGfZiAlV6N8ZyQgg8IULf08INNfAG5IvaeN/k0a3XHM
ayDrgyqLprhCjz411nzCLQjNGn6r8Fs+lKeBaucyMW9v6iGpI8tDARpq0Bk/Ry5X
icrtc+haa/yQrOGpBtUFgTDv2RHN0GE8s4cijjM8siQjHxVGa9rQ7F72mxj1LySt
FSN5I8UCMfeXHvuGY0e/HrarGCBJ0cm7FBwJNW0O6fdsfJLrxb/IY02L7R4N2Lr7
Ka4TYdtnNmy9z/3x+zCN5gPFFzX2B7n+2sDrfow7N5vp4J9UINUmqu+sjd09pZp3
twyE4uzOC8ebJb6FF7XS/A2wzpTGqLhVJmkTZCX/TuUgaaH3WTrU1XQN04JKtun7
mHw61XpqtN4azJuMbB7FQknhNHAdR5osIDMcwWnvdTf+U4Pyn09tZpCziLlEm8kD
msoAVoIfMoK9WOsfJy2Q+tCA5xuegABknuovzdLxQuGYtkTwgSN0v/vIU7p9lCPL
SvRAJ7OdvsvgFEaLaRZk+G/yCtlHDhpdJwdaUj5B1HR8VDOrjh9U7Z2CgF4CzLJD
RlkUIaIzLck33+UaHkHQI3ulbk4BQm+4dCkFX81ohJp33jTkykc7Fv/0AZb293Mo
gN6rU08eIhJAkNU4bbt/qPNbZyyGAzjtBF8bYVGczlUISq+m9fF+356Z/81Devb2
60LxhO3zTXFsoKyMYx7s2yAC9p1MGMZBH9Tfe9qgJ3DyqgT4NHskuf7SInn/GFtk
WpT/8fLv2JCcNW+WZlHHoyDD5fwtpajapr+4U/YkCkA2wjDuxwXtOJRHkIG+QSSd
Fgf1p1KG+zohrYUwPD3sZZ9XwrmW5rF3qBS4Txic18iSxxhYfNupBSzjoBLWwGwi
xiA+JQdxHSDT2KzUDW4TfrSMR0Iiju5Tzk0hKrXRZMhPNMPTg6huFv6CN2Smyjoq
X7JAJieQKnp13htlrNLs3noEWNIaOr3OOnJPOn6THnT/0aeBDgncV3SzcpfdlEhP
yr4lzPVyvZUV3JRdL7K+0sQSD+NuwUCSYofw9o4acDt62/3lkdofKWsyk6AZR777
sT1O9OeYIMOQRMBdkBlU3YFn+NEPZJN5QyjUsE1sefKfSDdJMzyqdcowD0cLGZgY
utZRlKRvbtVj1qUf7bZemboLXOwq+ohC5gX5uONWHIm80uuRc+DMR7kk8gtTSUnt
A4atPIPpeJNbR8TRDaZtI12R1kTa/Coxo1b/8KnF0HZSNHSriqn8hF9GNbla587h
dPheosCVJGkr642vp041TWxUHck2Vo6SaAS/ehOuBxHRikDnIDHZmAm/DgcLfOzw
istuLDydxXin57PRRvffOn6E766Ibpnnpaj2KN57pTkAWsOBT5pfwIfnXYW39jVT
IWw6iFWMnvP++oh7GzltU3j+pgicHrzPMGCxkneaCxWoYHMD5G4b9Yvf4cXfaTkc
6lYlG8OXFayjPDckHRC7HPsurs9T1ayxIffqBlQRoNVui5BYNHRCVVDQk+vKoPIv
IWDEoUHuT0Jg8o7LjDEO7AG4UxdiuXMg0QsEJDjMIxzDR81eGL7kOpoKy6zBlFkt
l8tgGw1H7tI/CLkVoxqZ5AWBlcNGmD4/IX1csXqhVOxH+hkeQ8a48u9IvhmdDuEB
rIl94XxtW7I7nD5VOskzjm+RNxGzHv4/LVPv+olm/DsX5MKp13rSt/zoiJetCDrG
CZR6W2SO9Vq8KT3lxzR23wn4wQ/f0sgVNCxWJfGLcqq9mOsoJXiYOyZc5fv1v9Kd
9xXGoftar+AcMHPihtTGZRRQJlfO/eRblqJ89dbxwQz2OzeO4Hhh+e3sdZGwsOeL
ujIusgVtKz55EX3lmgHqWrQB3y4FClQmxGoALVd/dKwWbgPFgQM3QeZbcxQE8qlK
LzrwbZz5M5H8oOvsIPmcRnfA4oLGQ8PZjyPoWgc1UECwTnfaNkljNi46RTWtbr8s
ICZF9qpqEhfPEy5vX2n6+5xz0CJzvzBwX+/mFPpBgpTCrCvHo06R9I3jwLEkUV/E
EbfPIwvHgyBqiUVwN0L5/RptnF6KqLQyvWN+YzoFuLh9XTTD+25rJFs2wjXgngCv
GcG0qxlk/SwzfPiw+zZomMcN4cUI0M8ariK8Q3m48qolrmcGhGJD74RbxJTb0iyo
MU2Lz2MiH1b0TGHe8yiHYIgC0iSe9aWTpKCQohCvhWBDsDNb8nn0Enpxuaa86bDQ
foVmv0saGwTvmH74ijOnzw7lIt0fnE098Euel8MlZX1L0Sf+2kbckQytZthvN1/r
oz8SSPn5h1UXvJtxR0x023uGzlfr4xgXt2o0Rr/N2dybb23W+nMTdSVViggQD0fF
3CWM8tLdGWKgbRlAvb/cddwaI8HFj8NtGjnzL7yvh0SGJ1dq0YyH3xYbB+qRRTw0
Zlbh3kZ2QNVJ8EW/KSM48rfm/Mpp/XPq7c9ZpMwj7RkqK61AINhKdKoqSHEpRdx/
3cDg35NuokwxS/8TFejs7CgY8vi6hYK5IfXjtFHFG70/QV5ns0FotWHl8F9J8zSi
hHuZUzWA3ngY22lu2CzuOEQ7mHSBaCmN6h3ssQYERsny6rEPxy0U5d763Nqj86gC
0pD5X2NX9J7U6KnHIWrk5xrs0wDftgNKr2o7O4zR3lfmp6snvYWZVqsc8r4MRNzp
djTstl/zpsuzO2M8ZdLac6mpVHLgrG5+b5eYuELbn/mypOEhTlMtRXQfbbk4D4x0
5Lfhbda+jynj1E9U0oaLytFKYJ2Dv4pyg9ms1X1rmAMp8UNIGnlfASvQ+YTyL4+p
afgDJ7ixjrkv3T3iLL7waFvCzYIOpi7t7BogU5j3znBfBcFAU37/bheUndcCV20P
5vyUc/q3/DJn4dCDMKrJusakm4y8ispR5kgJowamhj6ZFWaFvrQbv1LoLyr3fZ6f
ETBLc5telp4rFKSR2S+6fDLksaujSePEjRlEGRIUI8WEiYtg++pAAjkSLCiCNG+T
mom3MkJ7eesJnKMQ93DvHyMnCTjDoG+P7hjyoVQPrs45RHrIPUqKrBx4uz+TYkP+
9+CEQPa20QrQW+aP7NKyLLefXpUUJRYOko5HzfDqEOUiIV5f04/1G8vzw+wlv4gk
n0zjcZYC51S/qB4pkKnrcMkg/Ct8qY+uyrFum6unX2aEsi9PWHFGF6xTLT7VJBOh
kd3ff7TadX6Q2AAt/NRdt7hDyVYpZq9QGJPvNfO7531IxbLr39GXSCD4mAwsTJG4
1rzEzup2ThMc87m+vmDJInSPowmRv0m8aj+BoyfJIk8qHaocC33FZOJPNJb40/HZ
wsBb5Ana9OzUlZ7vvcnPXN7Oh/Z9xAFWgS/Ez2efIdrIcV2znlpJU3l9AtPLsaGG
nOEkBnjl+ZAOLrXymScUMC+aRdLHz5L4y40/fmR3wZya2PbMGXlsXZOZgKcEiH8o
o5Nf4oUx47lO9/2EhBnXy1QBRnmHvCxjxcc52+YYjRjujc/IGkPU/UyaUYrH6v+a
L8bMCB45Ta7jrO0DslLouvopIbW6HzLw4+jRprh02s0uBWsGDiogJjYOiogeEP7L
/bcTpBe5mlVelSJDGMx2VMn5wGH3kLs6Ts34ScaV2PyXdZsbbTU5faxachTgDU6C
OWPIxNDsFUwDp5owACDaflNQuu2Eu4De0MMQ/DkApJKG7o7e4BLK8Dhe1LNEwa4J
aRvTBNBmHIWecSv5UXEnY4YennlBs0Rr/1XP2TH3Q6sJxQxnzr+HP7I3BFFxn1eY
MTmyq0IFKeeL6G8Bto8J1BexXJFfCd2yS7VOrfA5tbH6soEceYIDmC8vv+7CW3pb
vCSVIcdaNF9nP6sS2DA1rQH4HshGmn+9RM1Y2a3kW3mocdEXwtMyt4hwVCQP4TsD
0YtjqcpesNGaYaqviTR/294/G5ljXeNL/+j0PoGGD4fQaL/LgQS0lPPTzw/zv+Sk
haOcQUYO7dbg6RABG5H9SL3u4mtAM2ffaGrqzmVbUkj3ByE6zeggE1NFhcBudPfx
RVyw/lQBJks5sBn0/XUqOJDcsaTJyhAIVM6ksKFgh2FwDy+jUDoYSOmqYbXnM7GZ
pXQOwyk5Hb0eLDNJA+LcWa2LRRcjjGXV0rCeAoW8N4rL6YhLqC/Pa3b7qsXaBweJ
ItcdCDeVPj0jeeeDZmyjnAiL6ESc8zvFdrmTcsFlE7/7kFOGkempAjoNbpAuNwSZ
lg7Jy11xQjW+bv3pgmUsQOhLIOFnaUdRwqMyn5EmLp26Xy32V7ZvIdJ+VkyZ/jCI
XSm6fxAwDir7sUPzOMY2gSKPvFUnngXlQJ0OFV7NvQxxqLB7eYJ8M2faNq3EoAR7
4hHMgNNvyzhqfAExAMIF3q5lrur/iOE6Ttm1bvhDF01Rbz0qnik7hTL9BIfEXaA5
vW+Ndu/+Zu2pZIP3kuOe2fucsYPGs6//gi4ZNS5o8UygrUhSWrvP8eFNuy68DULd
VpDR1LY063D+9lgpCknzi10LpFDVPpXkPsQI42MnMi7wTGe+AODkSaeiJ/IASoaY
yBDpWHl8tuiFScaQX6Mdua/CHYN+hYednd30CJJ6JpBAUXfTKVjq4ZEPDXIgkInN
Yk2IP5xYdA64Poyw6xnTWEG0p5+cJj+xOr/muwPL3Pf6i6hvDzu3C7ikS1R5EdM6
A6cIikTOnBfIW3qqB4kNQA6+qsJ0RnKk8KC4V7Fw7B3O28wyT/WMaseGtRsiqBc+
ky+FT00k6pMJ17PpPQUJfSKZp3q0ZQkMpQdRRAu2ROcZyRSACd8txewaZX2RYKC4
pfA0XNDB3HY6PigTOjkO+aZoj0qtm68GXIiSHyiIt/HcUJ9VyvaHEe/SaT/9OWKr
o9a7UoAPPaYCuTzdZug2dG/x8Yfhd0b2DrvPeq+cN2nWHy+MTIXQN0TDJ7IiDDcO
7gGLBiIIpKkmjmI4Q9Ga7SdACx7QQ7wkvfba41UqRP/cJdv1gjqGNrkqMsRENvHu
G++QVa/zfqgXw62hhZ8wCPpJLA4fPQ2jA9yh+l3uBTO1CIOr+wOaE2sVs0p3ZtOs
XE4VGBVMjMVmhhdCOHs7tqRAclBXI5dif5ionyV8vi33p+s9dW419nScosz4l4cy
pr4/aPQ+nA9Cq93IXFB6gjCbp8XkcTXzJuneIdW/sVEIXgampA9vKWSGn/9csT/n
BApq7Mjdew6j2uMYpgoGKz73Jk7GcSmJHQSDtV+BtCMOKEjTcViVifOKgXObrP5C
z+w66E7JlTxJNUcM2wtvSvWEQcfbl2zK7Mleo5ybVwlo22yH08kli8f4BFhqqZ0d
SWpK7a79VZt2RR4/aS5qDsiIL4mqexZAF7hVIrDVRn8U3plz/jo/JpZ7BbL2koi2
WFbdbXLAYJZtvflTxydaliFz4Gpm6kvYrqOOjmbJQEwx8AQIhG2r+hdotsfmwHRC
9ixCoCZsUhJhQH0Vo8xaKMqG0ik+ubjyJnBBWLMdPbGrL6rhV8ZeXbW7Uh9l6eEH
ooohVYxWQIaX99ork/p/YAY+hQwm69HeAGZhpTn26By28iMz1poQThEmdadnv1PQ
5Q9F+WScvzkRuXtD8eM5DdHKkdyqQi1PAgM2cUHmlxwQgfEcBhJ03ruep07bYe4Q
JE1VO9wy4GNG28ByVdREwyZjK7v+E5y0/UXAI+2vnvuK72IbFPt9A79XB2v6/ZlW
/QWG9xfciFXyZrATDKlKNMEeTLmNTw4Etqf4EfsjJenN/h5eyYogqUysqjoG9qie
vNhmqa79wfz9rA6dmRP7PxRN1+MIOVnoOxxBlrcALx6GM/F4uwIq7JuI774N4ZtM
L6JKQDJ5/pH90ZrzD1NpJ4ZRSTRR6dcBvQLx/m/BvNTPL2wKZt++XLgUDL+Oxeks
t7lz3XP5jNTcnCsAYIwA78Mg6IY47d4o7jBpO+7Z6EZFEE8be48krUMFKQlCFbda
ddqpdQhKNYTDekEwilPDoWAczxP88TYbYm+gIPfVtUjN0Bqaz0Jy4TUzguW/bGtO
onuvYReP1WdKN5U3fBjhLzpvR3tIH2iomi/nYbXarvCPNpCEdN3Dpq4Q9PK26Sc2
Y9Ap6IMhDuLVogETyPD+fOiG3kb/acgbBAazI9IXGwtvV7hA79ghaOAkgoS7q4RT
CXrwYsB1lwWCbFG0i2dSEg/txxWjCzKFDdta2T6cDto2QanBtitygspT+aD6hXaV
u33d3RzSDVk8hcSkBovxSFfdt/xQHGLCEv+jE/yVI6xFsL6PVV7Sc3JtuXspM8CR
+g9ihihDlv0IIy/HgV4yzP/U80Y/UWjYWSN2RjvjYGXBXJzIslVQcXDry0sdePh1
WHeHANO9195H2vB/XkJ2gmPCeL3ztw2KvluvMZ7MFeDSnxxIGf8q3oJNPZ1VYxYE
MDH8o0yeqFhjBFkEokwulD08bSDdePuSTeKJGgJlyVbMPLBFAyClfyC4/7CkkXLZ
StAx3XXcbrVOuTrffaK+bmOnSAW06VhKZcSfz86UKK0vjS/1uCPMw9+95OgInq8+
W6O+2iVjFKFiF/f2N/Co9B+m8FNo5WY/nXKj8TQsruVZXvSd/VvY0ZmVSSIv9v8j
fzed5mqpG9vslPost5ki6IX32gJ+G1UyG+xk0YVLbIDvEv/7Q+4G9ZWBk0morQpO
gB0o10RV/q1pY9iSIupQgC0EPFONtZztRjzQzO1N1IP0j42sA7dUV8F1ykS9rE4D
wx1NCnkihh7Gb3U3ySM9OQ+17UEdXf4V3pf9f9ZukT4RBcFSunvJ+WQlXD2vUIxw
A3IoyEvd3jtsTbTiP0NF9Fxy3+OWiBkrPVMLOg0SrL4R4+PpTtZd3o5C7LyyYASy
x6i2JfKB94mfIzDLs/2zjLjBf8wpW5pua2SM15B0l2OdjFPOzk7OmfMhanOUzYyP
fPjzgD1bic7Z+h/WnZmDjIMiY5eIq7V3x9neKl6u5mTrWxm8rmYCzjA8MwchFFY6
G4Ppu6v+BELucSZdJ5zPoKt1dJwqIn6fdb3zwWUvhRk7WTUbpbGzAndCdCtwOeiV
/efCM6VhNLFnv4LThcYDkc8zBDzJ15h8eMuQLd6hJApO160yP8Li9L6hUmHma26F
hNiGajpgfijkqMdHUcUxlEjdoLhb2rIdurkllNixhW0gPmOTDflL7/1y7mQAE4CK
EBn3D0lRCeC0v8AEyVLUCuPNE29ePPuB/3BWf1O76SCVFeU6yPhA5hlTttVIw65P
UCAMUBXnv17KwmlhvrxhH3WgAFZBnjH0SMh0PDcosvRMg003m+kKxlag5ftkr+lo
vww0BhqI7BXoXtrIjMH3+Y1K64O9RxLBUJ4TUwC58a9FqiLf8vrh58s8Tf+xNLLU
5ktZ90B0SpUQxCsutjCYs9gcqQvHAm+ZE19MFbnVqY7TQDWpcBaTRgGg9y67+t5W
QPWavP62FxOcGdJtXqf2ZAdRoFdye1gQrNxs2CCBbgmVnXg4uXlKM8fM28rewwDE
Zi04/KZtRoGtuk9FukXCXFZ2GfYoeNTHGY+eLag69UzPL9m9+8Ow/n2oZU+LSGqd
06wzP3kdCYo9FGaCTH3OhFAvVQpLk6GwYBWIWkUnxmB0AMNsJxGO0VUQhmIzVgAb
pwZFKbcOEvDVOCMaS76lwqpgIpMbOQJo12P8dp1v2Kb0HWu306cuGuozPi8rY3Te
3PVp8E2Fv1gR659FMuk1k7PSnfJ7GyL28rIs47VIW1zs4HWnz6gH0rUbs3IIjsfO
nxtDW1j1mm1GW3aHdjJUg3LhRl4mRyH9Eu7/f2e3rskT0PlTP8WU27cZSJ+MZ0qS
PpUxQSdQXvMXttXUzqAojHHX2JsD58f2uRJLvJyCA5NUJwOY8f9XB1BBmkWcs5Dt
cpSN24woF4PqAh4V2mlGYJgfy4fHMx54JefsxMB75gmFRZPFluOqhOql/EHb3Ooc
IeglVawO6sJdn7huGTeYBzNYbwvn4my8UJtTV2sKJVQm1mgQhiD5ySuUJlkCytqp
EDxSwE8Wrzt0DO6P034nQKBMof0Hz4tRPLz+H0Cwl28VyOrc867XqmWKoKcdBTAT
r7KDjmayD3a/kLxEr7fTEliDldSjrTSO8ioFQZEM2qdRS1BPaP3CfyJSy7W2hKUe
VIBIBvMgbuK2f6a4Pw1udjUELmJPVWAF97BulPPpExCp54Kbk3YReLWFanvmHxgq
kuzFHWoSNAXmSBZCwetOlxyqylGJL7722WONE5O9AJPikdXhxyHfvfr7duHYKbe5
zBuQwIHKOvuh/TQ2HnX1XRAJgNUlcMeE0l/0SxmU7bDHlaIH9lEnOvW5Bu6eDPjY
tjulBd8bhW6/5zB5XZwqGbachnbbgoJt3bDWMf9YYcJlZaQ4HDkx/rEJDM/soUtZ
42vwwtnYk6kPqciuhVKDWrpsO1Zfdj7VpK21hLpTymUwCg/igq5wAZYpOozB6H9A
K4mm05qyutoT2o/xGzR7hAgh0YsrgRGHwVeAfiYS7C6sJdK6YInC35Lkkt5baADe
F22aBzET4PtDJXJnniJuxvPIu1TlMV2Xudo42dhfroqmI3/bXyvaitNRkl25zyg3
dcS0eHDkLz/xhexH7xjdQ7S+EmDK7pOvBPhUdMNNcmOtthKW/COodKbjZqXdjoX7
9Jo74IIsSPmmGn9YTObNNvv3g6WzePKsiSpWaGdbqt++QZKuDImk8SaqxQaX55no
afk1INcaHyw37jFezphC3eHAVKoR7oVApByvDIgumTzrZ14hKcuWx8fQeJjD08T2
kJNwSzbmpP0YwY9TNNyfyM05vbq+LqZHbK36Nlwiq3c8RfZJ6IF6TFz75J1xj0Jr
8PghtgAmIqslk4rwkae7AsFRy5/TUhW8QO7mbcL5W0Sfwxt+Kctw6I19nKJRlN5a
ak3G48AIs5jCyN3trBme/xpc5s/r+XKI4Axas26BuOgal4S1UhDkIxwebR3VtkZf
wrBUMud5KDYwMWrrYmikLC6wcNjNbWrPTnvWV0zgNxp3xNregAgeSPnpzDtk88Y+
fw5aomekHr3sENOI5z1uNDntjGekYaG3w4vlmt6yHVrYQHfBTf+vUM9ZZ3zd2Pip
7hTAo18uhsfAY9OYZoZ7zZzKEevsc9C7blkXgyV8DX8ycenRzN2roP71XuCz/1En
mGt5G9uhi8DUpDbvy7e5SIjzYXlS8H839VboVhe4SILM/N+BQvQFzl0W+/77Jv5W
oK0iGdTiKmgnWxCJxMTWNNd77knVjfJQqaBzQZZo+k1dkgdyUMcrLo95XrPbRZCr
XxjnqGlOBDSHvsni9Nh5N4m/KTOekLhlkPGuzAg5T2Gp0l4nl8SXp7P1CEv3xPMg
gE5hQaEm4AepZSuWSH/5eSg9JYhJ850P2p63DD0QFsV78mkqP/CHUSLhNmmNytEr
MOBY2j/waQFq+3fiEINVvGqzkWBlbFjk4xiInXdGeKEIomx79oaerPipukhL0nm1
6C8BNhpF+3P6MvReuW6MwhuKRBhxHwRtvMkEPtcuGVq2L6/n/mhLVdXhyLv/Gjms
h2quD3ocxX6X/Lw/UV49oftF698/FTz5VKHAFWmX/F1UW+J26mrzE6K4t51N06jJ
uMXkU+FFUqaeJYv00ZKy/lpTAtRAA74nQNIdTGAyvO7QBlfIJTej1mvv7lBOpKPC
qb2DCm4PdjNvSB4CyYe+vzXI3RchD+5TeBfZPzaIjSmDqbj8oey8I2fELqiSoTb2
AtmzpgekvhbezixF/n2uxwQ1F+4JBcEp4XQynJcXEgm04a8NRVmO1A3v5N2l5S+i
AIFmkaG5iZINUi/uKCx+OEsnveoxfJFkbvLFK8D6ajrrk4LC4xZ8ZRRZZwJm1lv8
szs/Rlj5fuEPWbkNw+D1mYimx7WC6tUJq4t0X7Jz8aQ8shoo2ZoRmBxEGt/o4pis
Zr7cVJ6wqlvilk8gyyS+2SJtgadZHMFn3SPyuoehwXDDMqgnpa+jrb+Ee8TAm0Ge
ZUCxi93rr/nZCHx8CCXKIOq6OkzAgyZg49KR90SUGnjQ9mz7GR/gyoBf5t5ecJJK
hyEdanCb9ey1bAjlfRvkOBmW9aEBGHTjO4tYz0tgaizdC3xQ3GnRFAckJ9bspyYZ
Gld6swxXj4p2JzcD+LnWb8RW20XPVlra/FkIIOfRx3Vzr4WHAPFUtkVX6AMEwmGI
/juT1Lk1Kfc0JO2oqeeVUk+5uHHszWrmzQJueVWP7Ss+Op6IZzxeNahXD8UXfncr
e8+ZOnjbqAaOm/426+CfBy31ECTgR0dLHDHkTgXKGKRyjjWVDBoBwz+fsgv41+27
3s4TAE5H1vHj2yPDUSRjtBAL36eNBGz3bDDdlaPERBRS4ir6LqRUz0hgvccvvsW+
eG48MhFKCr2jKESj7xD5fkQzVZgaGsqP9/F0qBGwF64f1QGckKXS4xeU1TH6JzaR
MMyMTL8pQRY0Ohi8faIIyN6YWvip6fOUpvPBRrIxB64ywYmSRCFQGO5RAWeVkC0G
3GfIiX/dopqp/uy9CwNxLamAA0/q57lgMC3cuXHP0ayO9+wCpdzt2Z0C1qaNU6Wn
ikcHTAhDywwwf0a5pVuQ2B07QDn5VG08aSzgOoYBCLtz6Ss0NAgbI3IhbDStkNPq
eczmPXUtL4jdItfU9rAWdIrnZZPE0s/tVKFn6dWYEOZuP/2JJljacghZ9znercAn
ualx4f+9+hlq9aKyqTxh7qmcTWRsTAkjiW19j2Frab+3hNULk/IftvB6c5loZdKT
vw/qFj7XSfolXxuEEZhYfOqqyO/p3dmWZzB17LrkdwOaA1V1j8fqyRLUM9Hkc69Q
KMvqpTqL/QBee/6MhXhpgJSpK4D+sPm/zadMxuqRLLSu4OWUVbE4GBHqKhSQ/V3l
7dRceX/ZyXE2JzCF8f3vwRqPnnlTzS+jrFwYvXPT50axKqYhY0ogFG/ZJAj0FBEw
sp2jPGbko9IcNs6WrZuvl5L/sH/p2/+X6bPVdbYjeV0hEySTsVkM1vDeJH4dRWV2
IRdaDBMRLTsOlI6PiRc2uormbpLyaGLnAURi3sCOKUuSSq46rAXJrRwGQ/QYYtpZ
Gd7VWnfvrftSkm0F1XRZAO5b3Ch9U62PiCYrxkmxFNM+U9JVXbWo9be9ugSI7FlT
Uab96cwjvS9vT1oteLN5FfADrRRIHMJ/QBOZF0dXFkgKKs3SbBznPvlTdQgWc8l2
REfXDh6tK0tiW5RePuvjU0BJeNfaUNXA0e+k0y9hdd6WBrz7H/A2T9W6wqt30Pb1
qcxDOoRYh7thdzbWP5Acez1t9yS5wTEoKoIAPN8UnxI2WteFYnqDVuksMJtEYHsr
kDiMCGKtNyWza335Zm9+aq6/1aH7lWTWWVCO8w8+zPlqWSdcdz3JPgbgALqPf2tV
oYvEsE0NOkCfukh5ltGxJe1M2tgmbQCkKYYj3sVlTF9YN5TtdU2fYrIEJFGmwsH4
jexYJ5MW9mJmLhfS+PnH0+kZzos8VuguG/XSp7c5bu3BpSL5tgaGz8m3mAfpoNU9
FQN1yUBizPVeKIQAviOR7omNS0i010eawn9vtdJ9YDJJRtty5olKnMEQ7gBh/Yb3
IkJip4CDAcxaC3hzi75AKM76sYnpoEK4vKVk6JXHIDJ5dM+VQla9cOEmFEV6BfsG
LW/7R3lERn84wa3wTYkq/2SlxfAFSVX9kwSNMdHc5eRZpR2v2TLDnZpJ/jBfsenb
f0EvsAiLrnCaqNjPv+B+KkCSy2+x1PCFQV5MebbjpecL96W9kaij4HhExJmulSHL
BSWk89zo4tuqva+45/JbMFL1FWfFBx/pks7zEqysqfMHr/rraczdkuNu/NbxjVz4
gvlAQjWg//kOnYBiiIZjYIIdjrI01ljCh77WFEGJzjkcELtoa5G4/1D6/RxESgQz
Fu947CDYK8gCbZmeoO5YC0gHlYlwHw5uoEje8CpRzNMfUec9vKUUGtKNvpnkdUC+
N5Gi+VQYDvnYr9QQzEbzeuOey2J6phxa/S1bCaJZ5NajvHh0NDvTNNq/3vTpIIZX
rEqATnTCwi6tAW4BQ1r/l88vd40KZT2g+bc2hEcKt31BxL9cjQ7fhLFLdfY+xFwS
c7hGwb3MjkXoMUiL5IWuWes0LJuYI4GUNkaMW6vgU68ttgKEn/s372KLxuo4RiNh
a/72pkTaGnU8qaPrMzkb2bUGWaFI18SDxAEMb6PpYtAXCH0qRp5uI4Bu4FXIevJO
TdGxPn1IiuuWke004gB1kprNepk5SOlGLbVeFqpaeN6fnmMaIeMGXswcvlenaaOt
jp8R3iFk1aBc7S/wm9CY8WVMxS7Uf9uGsOinDbXhDoWLxfZXCOKUMQEJIIlGIh34
+IGO3iaMCGlUD9oHq0+AW9svhSS/h1zWy1JotJP6uaBelxvBD1J5xfuTOJq5XVMc
e+uwumxACDedhbx3d7u5MvME3+i8RDmrk7lbL2zlAMEzvQ0zBj5ZZcsXKAKiDMFx
iapBEAVkNoRzISY1uVQdWK3+YTvo0YN7+csI1LFWNv+okJhn7ntlYmGcosEM0TWk
U3DangSNYls2iiA9yVXsbwN92jrPWrg0QiRhFrPbnnRz/FJUIawQ/eIXqXB6Qoof
XqLM4gtHB8ChNXOCCwSWTtqn6KtceN0CX3dmCzjzg3IfAW7bcc+sGu3bn7MrMHVs
qgTqO/dx6Mb9YKrcwBVt6HsH00+zylFba720H6gc7bTzuoXUpkHpnNnGDubiwKzT
ijYgk1PBnSzyMYeBAMUAm0DrU9mh1UBgrJ7nD0/7WqfiNQQwRY+jxiWAh9cbNstd
UUdIfpqNuNp9MHO+eEIbK8lF6fdI955Uz8sPoS6EGM00DEZQxeS3iPsTaUVITIf9
ZgeWQoSSNYwBeWFASpyypmLMYogf9lI4/1hTNam/6PwhLNGRubK4Q6UkPGWfRvx5
zNzC4A4zAMdvSYfT+890YEPLhKTRu/o2uiPtCfWC0qlHGKgLunG1oMrlJuWG9SNW
TFxfgAf9WAYWIWWtTp5VdTCJnaDybdN7D6LEevpRylq2ZIOyg5R2nKU80bcYqTgu
NOgDeDaFYMtQf0m586y7sU8rvvpv6uepb5v7BhG/jdz9AfDWsehFfmC1LTx+UZd2
vvCEwWu4/Ml5LKPXa1v0nAih2u+LsqeXALG4TCNb8GrilBUdGaE3B7MDOK/9HGFj
HQPEPy5RSZGpHZV3a2vCiJf/Af3c4qCmk6qBGMNogCSfsGu07frMdkBnMzw3+Oxr
wn8Q70MhDTJmf8AfvZqmpHhdX7VrGShQ/EN87YSCqaQ+wdDWO4MfxtqCXN2DSYGi
DWOhYFG80r0VmsisGozPp9JByhmVCypjrhI8LH6Nxx871ufUZhmDcR1lpeE6s99G
6lfIl8gAUfAXjxoixBvVKd4TzpQzIvhwLDaL0r9IchdP7yzKLnEXYRJ11L7H+p9c
wHauc3PyYRECiiWlQhX8VV8z3NxKnZ9apq27J/qcirjNlVbzdrg7dfILn07OfgDM
AsguGZRrQqOHpf9BuuBcPX6LKXzOWxH2AgRJ12d1VzLlwZGbZ8xXzPMOFRYgofQN
1AoEhaCq2+v0PQLkYWrkwK8M0U1EDS1dVk/j8DuvIDF9NlPKlGDO55yMvz+dOtyh
HGDI3y6bIYdq/Tf/K++z+7cF3O72o0bb0363JkJDjOQ9021GXAJQc9NzMLvwn+nS
kcj5y9wofPVaIFMlDn2cZwnw8kfrY4vGjCEpng/4+RPDdLLgN2d6IvFuLtP998VF
cH7w2mFhal+yIORl7KiS0T4DCw1QB1iNG1Bk/k7iBJbTSe4DYn68lfGijN+EPR9l
uYY2KYSfYoR2VfbUl3T8+M6x6eEqu3DwyRlYiqNanIublaDuAbGyAPmV1coRXdBa
M0IcbbCICNrYOSrhF6OcUozRFx2u7TazXjAB22LxNh0UAqYlgBvwXCDHNBd4XAyM
TNxkOhOKPbgloUUb45RebP4nCLHTf5wgtaSClvyFTuR1RTdoVClaG4QQ2svLgWz7
xoZIKVRLqqDJnhY+uA1sbf0ogpusKkeZpT4RNGCkTxdm1PavKMhN6Ml22ty/ijta
233p3I4GO085tw3PZHpWP8Fnfy/uV+oSckJpwnW/hd/Tq3F4rVVkwEkq3Gc+qAGt
Jcgu8k5rnRXDlL8zHUrQONvaXnw7UKeux6QBHef81Ao6hCQNy+YZL7nnGA9gHjve
qKFf8AZxGm/em/Pa37Wt4Nz40ifW44DErrr1MO2Os1/evukGD/PJ8blLdQo9/2uy
OxRgZkmJ7SiCu+5J4e0+UY/H7WEINj5H6MTp/DrYCptL86Ne2pcq/pcxiVrTRW90
MuWkPJYGgZZZZbu17eHsSwlJLoipTcDMWK8ZEQ2xVhbsssGYfWaWfC2s4r5kyN8N
AxoeDJTvOjAEGEsYH31wHa1Ig/H8o3JIKsD1Fe0VpM6EjrBtuFM5hmIgkpPX7O3y
RrcG3y4biyTjhFihrS8Qint+QgwEvUs6JgN9PvWiIibhrJdAz3H+00fqGkTYuVWw
MQwaXd2TbxbdrOIDquRQZFaAzWuD42qzCMiktuVxEURS7a/O8/IFZN6o8DQUdTCV
i4udzgaBcfSvNv4Fo03oibuMmP96LDpPlWDf+nhCQjyBuyxIzSqgvnd2a6stLgrJ
rzB8MvDuhbHZEPMXB0VxxruRwDafQcKVLQlYLxXR4xTq5NvfZgleC1KU2e/du5+k
5pT8hJcSgax3VTBC2yHMZhq2xJaK1FRMNKQbgYB+vwC/r14x0zsNi2AVfvd3/Q1F
mdBNQewE9NOckZKTvvOIhv08/XXqpZhwPokdo6KwcWLBbNWL2nYb5wEukz6JjAvk
cYmO28OH92IM4bQeuw+9aSpZgSgYhVNyAMsUzPaSP0Vejl6zLuh3evIA2RTzL8Ch
KVYzMDzxRwPYz+TLKLJkoQIB+whsxce2tDPtbWaSw4esgoqObm6CFKbsvrBSXZgi
nXBC9w6gXraKqgj+dP943NYXpViLUj2vZ4DZIrO7xc550+vbQAs7M019oJBZNhD5
3EPAGk8vjraY/AwYmVdUfzYgaEdq1+Mb+LJVQqPx06c0EqcmTa1ChjLrf/5FejeK
XVZiSyz9EepmgAppBUO6e2/h5GnGQdlUyM+fKQxbgtYvRGebygQcQbsKQ6JLBh8O
H/riH0CYhqnEubnoPatNzFnTph481WV6txfjlV1aSWwB+HXFD5MiY/YQd71L3uD8
J2RFCC+C70qzNsixGkSsb5b/uzTAvbefsySsjLCKLxaeXmZgNumd/BOpfo5bwfDj
jmnpT5aXRSFDWZ6Ar49H6BSYqn5KKHMN9cxZl30+gtEhH+xGKyTwmhFs6jUcMGDD
tZ1y2+B98Y0VABtuMfPOWv+9LkPmfCHNDlFY2upoA3W9mPC0mns9o/K1JigIRmYY
PoIpgbYNJjpbYyFcQmtFxpWs2tySQCeJtULwfuwp1hs5Gdef51zLoQvPgc8kq1Sv
UAqENnQuskZ8Id/fXb5wXomB+8vbWW+H03Gbn5W1uaXNmHiP3tbfhF2LFJnxvy4c
Oe54jYPw3FoiKT2S3k/3t7+7Em4dxv1KbeGmoWaSOOb14xRJD5UoV016q5YEpN6U
B6EX4pQlUNIqhCISUxJoZMZtyKc63ySTqXFUOerbx1qW+7207i0yz5TVxPZboFES
/N7WnmxAQlTUOrXUmVblkq8RDlyzuJr4nuWVJ+WqpPa4sb+NxOgreL1XMARQFImp
R3QKpUOZoKrJKB1Km8V3rJUx6PLw3KBKITAP88hn5yGnd0exw6ADwo6GomUqJ/om
4a+ywSTJnDLt0e+XwZ4jeFEBGo1eglHeS675rDKlmQ8I0A9oi4iUWbD02e12DQ0P
jWOfQSIDNciu0VJsNj5LjlPvJJIz3CJfxzi8JORbQxt0XN0kGBrsCEGwKE+nIQg3
BFmR/4EogI3MABNdI2DJ/2Ks2QaRpmzKeucZyE0IabSyTKYOT3JJ4VGRFwpcDc5L
PFeVKIfAy4GlIXi+KqBh3gn3U6z08U44wMryypT9nSHbxhNMwwHaOeZwXMTWSaZw
NKYU4CNh0puJ920B4SnkR50SZyoALoTSW1SS5WFcV4rIlN7kBUUvZ0JD9ADEuPFM
ZN/z5sYW2I+57kmORMR8WKEO3CWg2TF2wPfVVo65n98an785X9mk/pV0Z9XzOv0M
8NLDm0/eR01vDwznOip6Eg6dtSXagO7Uy3PYRcT82ao0BsS5Etnd489mPFPIJK/b
TdYTySyfFxxdEAt3DH0e5NMLarBHFh2s0T2dRIRj5KKhKBor/hbzeRycGgX9Ij1H
YEaoGlpH7O7R2+nUky8wjJ5aWZmraSm5ibe0DTSUTyDWT1w6KKvbF857QzVV8ZYX
1opsn5ZzmVwZOXgqndeKn/+jknlowBbi9yqzw9QAVLw2aSPIIGc4/3UmSbOtDu7Q
tOHDDAwEue9LkMEDCDZIKM0qXT2D6aAKKR2zyR1WVm3ZQQTMPpwmRcrDfeE3xI8U
Na/jRx0pOlUPrSaTc+TlbpfrrGTQshpokFzqTDF7ikRt/ZsidJDhOmUWoesJiENY
Y6ICNZRrCdfwaKuFqO8NqscPjhU/b27JZmnmYf9O4Yab+sKBNkWe5dgc/wFOL+ka
esoAcWxpm45+noRGiwvyu3i6igqRGgJamX19ndq7ho9D5cAZVCj/3rybqzrSrwvf
Vbsag+V4qM40nTITadtUh8PKRwo3CZ3UMcQOSMeREKGyeS8/Ba+Lr13QLb2qMMWe
FWv2WLknLmgorLH/pZFmD+am7MiRNCu/Zunne60Cwia5uujtsrlPPQUCUWlGuDWd
ysY/UqXgaTxhNfFzRL6zX+VvVL8xXoFb6Kpw7yFD7iQfHQOj9sjAYNmYETvY3rG3
LEfwufapKMpDldVtQEkKimxyX6PXbD5zeWx5N3EZurWU1fOv5ppJaS/iJ+cbLYtp
yWnYIY2Dwn6Bd6ZKaF/ZsFeI4CplFj5gUmszrb0uf5fOqtq/ZF4V4arGkiMs2XAY
brrFjaFbVprUeXzP5Jm5byTCUFd5oMjWvFDTwB15Z86kjF+HG+y6cuBlpMxGUqlM
DVbVVX5eRbspSXQDuae/euCcyNYidsZUcFd9J+hZOIFsuXLFDZazKbQKIL4ximXG
h9y/nD5+dtMzpsip6cior6DBMn1BG/10AM1eRBkzd8HlIYSOfnPh6bzCWwnapgdU
3KVdAMMtmSzMU5i0vi5+aX/74O++ztPQOXu0jW/9oabZ6Ka7tK745aYTOIspYmui
TSJqA2mZZeg626euslp9g+pOssxRyvpf3bCbjfmddR9ifzJzDpraTv3UBhQ2oOe4
hSGHSVaPDpTeaGv7wdno5RkTK5P+Qjyn5Ysb/gooLyayHvjWAYEoqpXjigIpDAvK
dFNjDF1oIGte93Ls8cpdawu0qqDzY84ZVb5q+SXY1GrtDvS3wacVQ4jYqFN1lUCs
ofn+6YC9ORgJpO2ZaHfBNRsL3J5Nihk9pOThyzotG5NiMv8BQ4s13BEIHfdDzQ7g
6yhAiGG7veiQ68pcslu9vAAsF/fFW/zu5nJA2fcmuZMdp91G0IJKovQ8RcZqzSXq
lYRQofAOZOxDuZhZWjWgIl+NI7HPzkb8+Ofw+UuZiUAsUW/6ey9Phbemy7tMPFfy
WBeyEGsHeBr+0nZnbOyJZ08kY5IvJF9ukNUtlsjNMgRsnMYShKoPq4veE2AJ5Lqx
bf0fOFsLSc/Fe63zSrHB1nG2wSCcCZwGxZ4kADHgwEe1TbNC1IFpBo/b2CEE0fFc
YI7rQjOKsi/N6rDgsYjtToEnEtji0R3/5frjOlL1zJwL0SB1rDrju2EntYi00UYq
zQYtNGG7OxGI87Xzs2bFqpDTZoD+LxYGR1pgUnjLFgv85hQDDOk76I71nCMCDg9q
xfw8+WZWhpL6JZJgT/yRTs95CsU0OTAVa0l1/1Gov8diKlm8SDSXhXTalbNnSvLK
Lk+dk7NZCtjkXGIAIHi+xxxmtlzznKMWQV0dVulZgDPoKDW8jBSTzBvpeKEKQxv/
xjq70xa+yJ+03yc2m/9bkfxxqB7XGI2Zbv+uupdR1/qKw337grk3X7sLIgldZz5U
1xKBf//wag6A3a0Wzzs4sn1JsYLUqbm24TjZ7huRJExMOkMC34y9ZRmHRK2Q6V4i
t14iP2niL15jbwYSC4kncfk4CzFG7hP8098tgCbePvT0JE+6fDa+tkDMn5uM7CvN
9WvmM2WtwTVNdqgewrr3Knz8jqkCotue3PdbGJMj9W96ofkOz6AHp2t3j3nI/r2g
K3q9T5u9xqW738yKgkeMZ94eRyWHeogE9N7H7g1tAE2Lxo+PQ4zmehco2k89FH+3
yjbAXAywtvqGbBePG7Ls5gBa20hxZivIAP9AeMReUHxo/7vMsAP3iWHxD3YgFTJU
Jjai2fhnyxjcknZAt1/zJGuWgp2Fs3mNMDChyF1yKlcpVwex399OnU1FJiUktZ+t
7KNHtsDv42N+Vxe76Pb9JkotLvo9FJh7KADcL9AyLduL/TQ85f1OOtglb/PMIKjj
nI+3ug3ETkrcsmBA7ljJn1HePBFRhCUu4lN9pd4xPrKCVVEHjGDo3wn3NE6exTpx
O97JPSZbTOld+UatB+ec6+k59kFPMLIPcNgcMI/hLusO1mah3IqPOSGDIEU90PGq
J3hW20j9jiI34wAibOi1EHt5awBugqxU/L3kK7CONYt735CCVt6PtPKrtaV9CUV8
PIw5qI04GPYEZD755ib20qf2ECH7UT3CDMkK8RbjSJPw1WccOPe1te+kX68u/ADe
qyxL2w7HFJTWMCDrO7ovzvrYNRMGSgXLiAZuw5TbbwOAmZ1B9WukuXXgsJovGZt4
kok95/r9Dte50xfWwcmAeGldy6FgnK17gQjkGRGqdiE+iMNfdBM3By8C+9PTV/Mg
ZuehjP8cVSUi1azYh5h5X12IJT6qECh35etNVam+78paruLGDMRGsAaRJnoJd9vS
0WVNrUmZjuyf+gIAdPflkIgu/rhGK5bLOLztPhNKzCJZ9UGc4omK1UtKy+4bwYOr
VaXf+MFW4qL+602gw0tX7HJKegMmFYzHwlmUyAixBvguls9JhR/Zrs2Ozuh+zD1b
tk17fobIQE2OALOmTH/OK2qIAZiWTbLfxAT6/R5u8XQjNAKtngckk9kokAEsXru3
Qb+HVqGdBawHd93+C/9cf0e/uy1s53Sd7lmcWLO9agU4OPFJW8In0mnxCyq6jehU
ZwUxBCVPQgcTZynCA7BHYrVibShp2TwqRQu4mjHFMeSYifxC/QH7zN2Xf64+vOEi
MQp1mFEvokDbBF+F4kZRMQpj08RoMb7LsYdqKh+LaZforJTkmeFNGm3V2/0wh0ih
OgxCoHuuvCKwZKKJhKzsrnzKdS9Sn4yls1raXpNUceK75j7LC/+sThiEMH18O9XZ
GrlL63fvoWwrstuxm9AdNm/T6G4y73AcP6rM/DC/212MVjauX9qpRmjCz1WE4vzM
h9VGOnrDDXicRXOH9lUTYg1+VS7p7pRQySHxnkSgsxSiKcE7RfGhLCK77WOUE6JJ
dzWA+g40loCJqAkCvJvTgSEyKZuLKD79HBzZB5MLyopSCoFah9ThnJHlwd7bY8iy
FUN9UO3DFjVQkyT0ytGzBTjuBhC7k7IF7Mf2mT+61m38KjPk4UcP6dULuTbOBlE1
5x1sPtqHQFtpQvAPfHSnfYp/HrJd8DDHWoj/oBWNuLHhn7ZFU4f5cXvUcFK0Imj3
bEpqb2IKVZh5o1VUojMIp2Mdxi4gagTzIrHDSL86GeZPZ6nUjYhDenk/J9Ajs/8D
vZxijnKGzd78CnYxrOJk13CvCaiGTCWcRigiGTlo1oGQrsGmcfYIyVTCLUZ6GCGd
8H8BHn/+/X+6CYds4WMHR6b2BF5SWk8DS+DDb4ZN5jl4nzhwKfRA9UDVrSEsFTFx
5miI2ESYwpVFAJiLXR8BCy5h//0SBu9wcVzFZHDQStbo23qWknTK+obOKR2QzkSo
P/sFZHNBz7Q2/w+0ffjbAbA90mWN+qDC75FXV43VSz5Qr3dIoE6MEZqv9kGBxFCn
955A8w1K5h40JnEp4y1gzaJVYnIN7QN6c046ZFfSkV3dTORjI8tkTIKQfLz3nv9B
7RNLOplvq7+nLA+sSjXepUkgzv3O8s6PAR2noCAwyubdLEv0gDZjozcAxnvFf6L9
QcISz8Cdy/DI3cDnGwDRw0QlSNnIhWV/7CWm5ypdXPhYcSdq8FsxehlNDEYcNzQZ
8QiCp7t6qml50htxmc5syPRCJFL3O7hP0FqHdlA3eLEvSZjJDbUKoNryXyFRkFnG
b7Pdfk5W9giUamj3G9MzE4xKOkl8LPMtJMzEWDkEEfg2cLntOTQWPYtO6la4g4d/
oVXSK3FgC5AuOU0lWZFj1bVAfRTSn3CZ9uf0WToB2J2Nse00qtLAKzln1028aPoC
ljZf3Cis/pUzqsDWZn4ddHWWg8Pn6hzP6A1tHIaSUg9JESiVact6synoS0Pfl5gx
SnMF6JY4lbXz6KaUGtpeHzgcaANZSH4bSlhNdIFf0OaKQMoW0NrS0v8gnkrqW7qG
yiuYBXAPRPOuF5izhvh5159jcyjLyQmU5zCMZgiFd6ew0IS172vlFd4VRGmVY+yR
wxBHGW21R8Z/DnKcFUa7SoHtzjYglRCqLtL7+xBzMmMzdtP+NjU5dygpoggtBO4N
u55hd/AD7uy3KPCrdOz5dlSF+gQHXU3+I3XC1z13AJWbvYC5kOFPXRPc7kJienxm
9PhKZ1oqzn7LOT15BezT9j8mfyYtGEKEMbJKqntTs2ZRS9RkI0FEl95PJSW0Wpx5
qfKcFex0kkSAcB/WUg4w+1lTyMLevnt+4lixPu5Euafi9xB/BGnzZOiVAGTMskih
dQVPivKBxS9Ngjxziase8X2C1hRaI/54x5fIkevldIZFXfF6SU+47KblUsYxrwl6
iwgpaRG5wYozscuTqivB8WGVUbLiUTHy/rgvHdJshfbenVMEV0GTiTe9byyqXm68
WmHzhMVq4+Ail1AE/p9WtX/kxDqVb3dXaqGgi/gFKug+y4D6tGYLFCRT8iYG4cD5
IlFfbpck/lIxZVAg0g5rcnYapelmbsrPiLUF8RyqJDKdSofQt3jRcdyidq1BpMmi
3JHkSuEBjOKY+esqGiJCyH8vesZBJJ7mE1dLRU9wBsV2iOXq447yFOxcKtv1Ed2I
5XPUIK4UOMc8T3WiR1uxvV5K1K0loBJb74KFOy/vTEVyYTw/KgQhTD5eZIDlZT7r
SjwTokhwA6shxHvSTbJVh+LpztslqIQT3UaWA0epEbeld64dSkMen1AiDszqsnIQ
Mlwnfi8hVrgFsZjIUkV+PkdOQVY58/0XMsoM09XLh0GT3Xto9NfiyOHVSrhay+O1
HOtFjdzWdHWuV3tLtQLpHTixMSV46gaDmFw9q20fO4vNLNPmecK3AYfI4EvZGoSv
/FIlaLdemYYJCiEyF8CwdzeQvX2agxiplGZKBNjYMB5G+w7ssi5jcQluWM7apszh
H0pKaNJ9x2H5MguJpHiE5HBuLLxtjODCTWmAM4G5rzLmcdSULfrbWNmaLlbiFMBT
swnPUXQ1EbeBQ/6ShR0wXGHx+lm+J8S0UtQhfa07voeNOqh5UP/gzzCWlPH7n/mB
bbzo0xJW5EstNaN6X9GZDLoqXsMCY//K2Bfnlo2iLATxT47b7ZP7rX0MuWxFl+W+
gFYS8Eap5V/btqDMz9x1Q3/lo8uaWnTJpS7TEQK44bQsTghHDcBqkiRBy68uzJTw
n5W7DrYRaOTjt1IUhxCaqJVSl5VnsFuFUlM7HyGf64AmOjmsQRCYco1T1F3dYYDU
FBrHHWSSvf2VHl/MCcfh4Hr3ZOY2sksOZh1JXu9PhFrQ1XmZHsQHEAIcv5rfhQWz
8/lG+xPTZWcEQFQhsr0RzPXlg8vl/ooCasjdEZfT8lPfdptU94CqRmPS6YS5Pe4Q
2E30/zZFTAe6Agz9zex5z0hPz7YcABO17QHne2Rc/ZCL5kd2apxTdGcBIwifKp/3
u1Rc0dC69LRH12J39LM0J/YA4E9NPGi4zusHfheQ074GDcyDZsatmVwsHiLmTNoV
xQGD6ezITxrvXO7mKCGKOr58//3XzwrGHXQXYvcimvki7FzNly0JasRPd0oJeT/m
JYd89YgN45T2f8EmiKE/ygF0TwjQfuEVwFpNrKw1BEWip2ng5awKFHrmOs7MA7IX
6C2dg8lWDMkvEkrhGueBseZcl0aWxdmnikLHVDy3NOZYpbsWokHyTtdRL7c8q7ao
5SqttsK9vz6hkCfJ25tgHpwwJS9LWhNbd6T2Plre/X44lKWC7ERR7+jK1CQVMnEj
xjvppr6urrowG+13BPCCCOy3bsJbj2xJkwLZrGWa87CRAJh8Ei2h4v+NMYb4UGx2
hPfPOTk4AY7sUN1apgL3PQEP2o/Dzm5dkWkCQzWF9CEOtv4tiBUUW1zbfETvdouG
5HiB2ZxaHrH72Qd7I+o+1HxJ9+dCrjWdGPY8IiWCbYPTzu9U5Dyeu6YBnT8DFKjB
J9IZ8h/kL+VfdGlKfiJJOey29/NUhYOTmKHiUsvdYe7rMEsMGsXcsiijs3SzWuXM
pvEHN5+yljk8pUtGKo/oIQ/5wEDIRr+sLj44MMBS/oByU9jaF0a8Mu8m3jnNabvp
kvK3F3XOMWykqUUIu/jPtMQ01fclqLJ0ptpqcIgleytlvLZTCV1/YRDMEyYmZ6OA
jjoW/lN1oNFaRX3WWBRADR8Rl4EYaxIVQp2IKhflg3aUZWRgM4aZQBKCVEjAGzMu
vG6UDek1idJTCXL2ob8CgRymC+unj/SnEeJjR2LnVADPHRVnWCdKxlClgY77tqTR
ptoDw51GYf7eK3A+86saI9GK9z+790EwxeQtkAH9BK4VwMqXSzGeGOwLiN4BmvL2
P0Y8JIJzdnh3d1mtVjcYUCKruLw3Rogo4PrCIy5i8zJwRnEbDwoAtREK/O/2h2Rb
5ySUwr1gvePohAmxYv3rErCHpkHPrmhAXEUT6SDgUh5sXpRj7G8XsUyIDLYGg+3I
my1MNQP29XIZjX3D1rrsuwIFnzwu/q+8AUYGEjhQguOSN9sKWi+xA0TeGPYeyxmq
isVgugSJVdRy0QAONSQ1hnxBclbJto3YNoEfR294dS7T6txj6ynBuD3sOX9tgG4m
IM9lRd6qdI9vGoZaI5TjarCEbvFwloJ5P9xIxrtXRiNg129ylfPg+G0oVwaT6gZy
jvMQyw+5PFgvHmCXnfN10fqIwzxV6jLWw8gbOcCaK1yRrHJe6/y4UYOntc+63QUy
xGdP4kYrDvwF+aI3bITAAZPfC+qRnXnPMUDik6p64LqVO1ppbk1t9eVWlcq+iHcX
AhXwdaxxPUDM0aL3aKEV8Yje5W/HYJKjPrMMNrX2V3LyVrosdMoPvzvKIpvtudNP
R1f90rXBK0tqlx2v3PcmDFrpAYDusmi2/D2JTcOGWdxnJkl3uyYov5bgSHtRkWcw
plK/PU4hr1nxmZ7B2Q9Mpfyt6B0vC54KBQxJNjV4Gsjjiw35nPFULbVEq3IIl3IG
BPw1bpfELNDZS2+OQEDABHJAKW3l8JMPi5NXVDV2Ut9mxF/OIgiS/a0ZydaCGnsS
PJ4pJmcoLyWSxWPuw7er4oqBrD8r4VDJRikH5P4GpL3y7k5AYX+85LQRMZHCxDA9
/5zQLiJNfeOBEEHq+5rPca3GhhyVAn13v/Fch/9MY+XACR1vUtqQ6eENy8lCEjKS
9aQXv69/jRaTMwxw74yby/APA2UeK6KcXuwYieyNnDCd22S6cZkcQI2WRBJVMFT0
pRyQHTLNgxAIYWp31Q681avrY7BLACZugm/8+udWXI23eNchUtBmswd1p+1l8Pqo
ya1lBu9y3EyPl7zjOvF4n6S9hv6eSfnxFJIDWxPhnM25udf2XYPLbWA9WtJVKXO/
E89ojYFCTcTLpNM5+invaKTMOYqJyVfxZebDkJFEJanZtXZ0TNwmBGGZZpY+C9V2
aK39yDesmpQRi6qQVE+zM8PI0PYon0yBrIytvXlSlUrKqH6FIPT7omGcu3wvJZv9
gs+v9PTN8PQJ1V6mNy8x5tC2AkenwexDHl7pQlWNrT7S+svrRRak6XLmLvBNGzCL
BQGfpza2kZ/4+L/hitydhCo/wMPgzZQC5vnOZf/wpDVj0u69Hs0dMI82JW77LzKb
f3Otrhkxcli1x5DA4lO/QmFJgDCWcs2P7ZVAnguPcA7ai97ivSqLPfDxWkKbcTfA
EE89wtJXhM9K8KIgxshzR1/eXQRJ39z2rnlJTxrh+824mNKfjYH5Jqa+OvPo7dOV
tjA3UY/K3+pIKGA5eQp9GsrhxnlWvEFx/rK4PZOY5u0QgArh2cw/DVkz4yAEz7jV
6bRwZmSgBCA9U4WK/QCtBvBPFALBqlKnBaISGkOGNyX6NVxOLfYtHjyHfD/OX4Mm
tGKI1t4BZWp/HFiLcdhEqNP/3T6JmQLvl36/OTo8mGf9472jlCfio4SFPFeA4/0w
CwRSl7GzH8kyKZfpXusROla4zZmSBUVGEQQsVX2sVw4QAwR0aWn8foJEovOmdMRb
lojjIpYO44EFOm5dscV0h74FVCsD8iEC3qd13a8tJVjADu3p4MVsCCgtr3+h8QMP
run8b1MJqLDjjjg4ptI5UJcL6tIDHxMa9ynFvguoC7+HZJP9n/zHkkJsqIDPses9
FEObEi+TdRq5dqJH4OyHqgAc035lkT+wGvgNXBImJnD9pjVcuKdQ7KU4I0IY2s+V
YoBniFz4xoZA183ZvZPlFFTu7mSq+5/8oM6wfKFPC0MyFY1VIo5DCF4UJYox18jc
MW/aBKPwfV9MI2USHzSgTPmxN8jLbYmoeL71vxP+C/+yazA81UJrfjO/nt7o8t4V
wLmIxpN/8cxyk6xKymsTJ3f39jrmmS9Ekfag0/Hr3aWG+Mf/CxwEfarlbSKycJeW
hFGi9wSe2XCs5uaZ7bEyPIbQvm7d844utnqkbxw/iYOaoIDrqNv31wnAfy6uh4an
Y1+1R9mdWGqEDXERRjutfEtDSHgpYG7x4zJuxhbFLXY+07WjEroYxNRmwBsRgfAV
PIN9icgk39CvIfN1RrcbMbM5xcPdJYBUsIxOByNw30CBHS7UeubQH7exKmhGZ41T
0YSN0L4Jbg3ZJd+mUEprylPBH7KxuWPSPBLHC3k+6gxJ2mMycIydHwSrHPypyWdf
XaQ/ET9uWX7YyLuWtfG1xuOIgszqXOUNT5u8CKnu49xV8sb16kQOSOicJbprGvh6
WilW4rd2cQ3dYR6nK8s3oEloRae9+uJkwJZDEo/trUcrmPdn9OiRAxDXypdTTaFU
XZjTVVZypKVYj2zi3EiuAsccCcaCXdfsdpKY1rjDt5R32sznrzdn1h0vgIYnf0AC
g854J7RKWXNgnAfG83HhUnST8D7JcDiHxC1s6JbyM4eKuBOkGTxkJE3GAzQd2hnS
HGJqsWbB+ZGUc2Rkj+YHTdgz0LeztwOkVMpfQoIgvtf7SOwzn7Zua2trSEoRy1Ui
tOOEcfgnGZKWk67d9TquVCdLx4LbCRRkbdg5xIRl0Z2llVjj8xHFH3EkSlCucUda
MNSurE3uEuS1NGox9apNSFtdSExGsshPfTEFlUNK9Uj58Izkb45kpI254ViuyiL3
htpSUsUida15vCnTRu46iUql2CBzsq08uK8ohZ8gwbYw+0ZQYHdOa1mPtD9/CviT
uxgqepL0vVQMjtNMw3oV0ObJn8mkf/RgT92vErb4aavyIAB20QLilg2wcEJYynZx
5N2U7GBFtTp4sQ4ZLPB+vKvpXHv0cRaryZnVy2Lwv3jg2iRVlM7qGnbktKvFn4cz
1FZA1XKCAHCS09r01nlFv8A1XfinrwNPDSh79ehTuwjS7NhQMPAV7usk9e5WAX91
U0MzXGYOV5IlF5R2u2NZ4eyX/a2nEN8oMz9pcua3sUrx4uyIXFF0DtGK1B7pcH2u
apor4C3iq6H07bKkBk/GpRp48QGhwJj96nFvI5xdQYblrr91DiK2W0cH3Zusgzfz
7W6ZwG4SpAWC+wLntb8NujOqWLOgrwHNq5alF6gUrdRpIySHpn+tbpCdC/xpbrcz
+52QNNTbIfF/LjE4lWTplAOyuK+S+/XS27e6zCILECh8lzh0hZi+XCR1W5Sl3Xgl
ujQlV5RRM/07b67IMwu4p8VU8E3N5iYv6FZXU/+4SKy9dyvwkjG+NGsi5yPtuHsj
8bt2/ANmD07OMEELD0JyBvNpMXfWKqr8AftAoS3XnvJ4hm22QzsgMprE9ULQbXm4
NK9ykPc/BDSmSu49fc4CNrAq57VkysWSis4eBWJtl2PI6QBxuWBF2bXYTtPTJaJb
nRCeyWTsv5QXYyVr964dXvGAyZ7Syqp6qhM2Wb0jYD8SL9K/U/aZlukHCCMJCINL
G52hKEmzaeZyAJGrs/ZhVUnZlZ1VhJcz2APMITzS6W7+GrKkAGppJsgIqJ1jrnL6
qdVHERu5dywxOBlVlfK3xf5Z/Idak33rORiTI+PXKR/pQtETO+YTUjmwnG7BNd65
BNg9seudhYpuNEu34iEOaxa6YVOGd/azGMFUSpW3ced35CP+qWnNSiRjoBDa5t3+
RszmyNMepLEigk/YOtUkMthtGY0Y1Vw5kyMh22zgkdfTBm7nF8Diq25FLCGOjHKR
JAu2tn4yOFKQ43wNJsVAWonlrdDtFGOFapjHt0Ad051wSZCGKgCgzJvYuopYWgI0
3GBZjGxMFRbako7C/RMDW2AM/EDfNt8Yt+p+Vx1+j/Yu5l7mhtiyrsV08IdUeYfH
NAGWv7owP43cEWTllisCn2TYgYwaQCfRA4UKeqBLRlbThAR1bkRQXhI7Xf3WOt1T
uISc8E91Dc8kB2ZlgDtGiTATTHVNJpaf/FWH/bLgkYCk+GiK/NlMQUjWyq/cHODW
QMYE5/giidEsQg+eiS1hpfu9yFSd06569VdXqBJr31wzyujLFBXqjq0bKeUb/l94
V0t42Wlqo7qaRav9j5OcU3zekPaHAAsudBPwbcUZifx012iNX8uZX7lITbC5ODnH
oZm2VlmSiCGmZxGfQUTj2rKkzvkKtbwAdFbNe4eyRd0ibE8SZ4qaDyGrhiphXqVa
qn8t5caJNj//Its7t4wcWX1x+p42pzA6jjJWoPEJe3Anj1LsVWf7BJjRpTvsCOvq
cDpX5bxq0+0W7SVBdWfccVzYHIzDUmSjURLY25nzbm1p7suWx/RSv2tl3kpyoJ7b
ni04ZMQ3ij2ARJDTU8nvb3OHvBh4MVLr35xmuW3QfiopGbnYa5ze/mqp2BOEacK6
HzN9AUJWZulDVVJIjj7VZYuFKwxeDtdMwJnY1Zogrn242Dw9IDzmIjGf9xJ4PPRl
c6+gVWCJcFUyU+DnO2hugJlEaBQoOoH8YYOY594WXAtVgNcFHMIeWJ+RQu7n2Nnb
nMbENLQH1dLwvcmPqubdZE+GvbHCnHKpK68VvcsqAPMLEJZkqGJHrLHnxcBtUeYy
g2l+I8f0S98P3PrHceJpRO2iXOvwCzGKHAjKq0booGtzEV2i3tTh7PwyyTZagKuW
vdXy02dOmg+gfdeNod+rgoMh2fX3oguMuTecHzWRE68JxOJk64FHKFX2Fp3s5qpm
M1ubUQAAt7pr79ukTKbXYr8bJd6cnvzpexHFqXOOU8lL/N1E+dpREKnRSZIBm3N2
aV4CVujLTMh3ltlONj4qo4eLkPUWe50QmyAZjeUElpbw/2i/KLKnTOsVzwcNMM7k
m+pALf4cNIq3Eax8SHj225HD2eXrhdGr8edg6hmbY7xgzIT2yU/4Wc2YLY2iAJyf
tTReGesP7IQ/sOt44Lm8/D3yabU3tAxwIdSN/OcVb/ZsfyQ/yZRhVBHsYMSFti1u
oZbl9bxhZ18oI03UnP1ySF/NB97IUlPHuKMqrX1Pm5EPbudtKS2kfxICJ7ae03Qb
xNAX80/I/Ctc4nm2KD+J+eIIRkCf7DHRzYYIFUITUR3IVv6fB639aV+0+OCzND9y
PqWWYdshZOzTo6RtvLPsRid0xFeels0SUsFUT2zRgi/IWNCXRaUdSUDsIWDXbyMr
IWZc/HwlVNnW8a7iLrvCC7CGxRtUy9xKZj2Gyr9qRsBNinkvcxAXbzf/tiApYOwl
vJdMlZWIJCAc8CPwK0lgbTsL/e1Ro6y/CBzDf14/l0ySdYcW/W7AUOu2D8Ugi9Y3
vpGSm/umpwJSQz5YLgslxhVfziaJtK1fmJMjhzW4mDutynT/JLTae2ZeyTUCSESu
c7g0IFe0VSah049Q/7yDSP8RubCkWMq3hSG7rW1lwTB1iqcsiQhtyKCvwVP/J0D+
XkKILXXea3q1dJN5ADLfhO+RRTMsExV+Mn32H+HuxDt1EzTq/BqbcyvbojndFF+o
S8XBNx+W3W0/w7TLNJYR8M7V/16+A66yEO8aLU/fYgGmK+tigHV+B4Dbp85p6/W/
q8qM0+laipUz/kKWgh1S7IP18L82jMZeqC9QG+QQ35lfy8hdPyZieDn4T4da0M5S
k4JYYvB8DUPNX1khOuk/lQ3/xrkXFt1NnLz4LixYqSn3I2M4xrkM8x3nK+C8QZ3a
QqFiwZO+7hOtjizJojXoQavgt45tVKArKauL076ykFDasjU1Pg8I28jK6deBG8GR
11SXEzgaBSHoV9YWHHCLll3z9xlotMeNea9mkUpp9tfKdb+UXjy5RL7ElSVXVYAr
yKHCyiBSuQxk5ygMwUNkdYotPa/MYfM7z/iEQG5CGfJpqYSBuCWPr9ztFcWVleAk
VHzt6wvXIrf3PqsFHQ5OZNocqJfiabsADFSnjxOo39Y9bdiBcGIcf9oSdQt8tiCI
nsvSb7vux0bc1CtLwIa8NS1mTOEGWUYBOSxrk1OesdEDyOWYtmO8ZBq/KxjY6bLy
mtTaKCr+eU7RV+pCvT6j8rk9nUT9dL4d4oTcfo9G1ND25AdWsF9EpLAVqxAA5OMK
LGq+GGYkpcvRNE+HTFczEIR0kgtQ8dmzdxOD/y/BiSST/JHj1Rh5EseqViOMS+sx
zuGx26/g54/wXOnZ0yecyvYsXJdAZRBo1OCmKCfVxvZFHNhgLcKx1lIplBmHCzX5
R8uwxAN8E9puTlGincklZgS4uqFEjiC7hhblGJnfDpxKhqE0/X4Q1pEQGYqknMXw
Y6raE5MqSVBIdM8/E6A1U2/fwhUQ0CP5iJZs0eW/VTfiBwUlC/BhS2vQXeT6Kily
hSEAtl3SeCq3gtxIZzkChDHA6b/D6F+1vfs6tZz9QyJb9QdNkgWW5N8m02y3z8g0
pyDmRVbPuWJ25/NuAkeNPXIpkkYZ25LNZlGraQcuI5a1z6GdTtIWnIAcOrbIWoet
DHbJjPuC6fDw4y2AloRcEzaUeMiN1fbZQp3yO+s4w5Vcpi8bkSZV0J85e1a20Y/t
bbTRo88x+Dc04d6Y/5dVBr9NzefSfNAMzOtpuWAHOHy6MJK6MAH9dBFgX1AdIO0M
DMBN4XprTWHV5o/bKNseK0IW2yi3jQ14KYcFumLRisEBPaWPBd1P3ara3kFAw9BM
QBI05RLtzEJaj8VX1vU1ZdCU9Sd/WvfaCULOuWarcSrIvYfZW1ZRwaMjwkwmkMR/
eOgJHWrNm4lVbeexdSDZ8qSnjrIMyzfAVW5uuYcd7wJiYg6ilyB+RxaL5fIiCAiX
gPiv2dyyJR39thuNuRClQMd9gCLFBr13y+gqbfTGFUBT5rBaP9VLTCW4gfPgje4r
HzlMq41kvDucJ3byNxiJHseu6YQs+D9AmZLLVsa32Bhl6h9Zj/e5xrvreIQPeVAz
EgndrhT4puw6y68Uc0RIha2pBuRjjPUl+2zcLQVK+PaI9DfXXOpQjoTlLlJHehuI
0jbK+i8RpWhqr0CzuWp9OmoLs4/CRyewHLRTVIVeiEIWuwJ/q0ZfH4IcgNShP56f
vaJTCeOnh4C64MsHm5bHa3bBYlDDKOsg2Xu2UuRYTPGTlfEyXkGfLGmZDEXxJFTH
80+aFvkAaRXZgLbzNtq7YoZL+7HFwbheX6pFbIgwI3On1hVxtHXt+JLOcw30aIHp
6/2hnliegosNIxlezSs67F9r7M3Oor3voXy3afVm4UcM+kPs0JTAlHZnPfXzj2Yl
fZoHeFAo92mOQgdTqtc8fLC6jQ6U9KlXzhe22QgXDWxbYP1M4gdYjSM/mZrfH7E3
dcAKKWxIgNCL6SYtZ28WBYnU8QO8ZKGT9fDv7DncJp+6Im5BK6NG+gB2iyzHNcUY
vyhjAvPKDeZadztkpA0I9BQjOYd9a+n8h9E8KbOt30esGr3P//OcEYwit+YeeXnj
o9iz8Deqfww5scsWc/DoFTkuDZVgSDHSRdAGursv9g7aWq+BDzLR23JtnDutEMND
umnPk/dmnXYM0q+tbcBdl5DZaJeVMLeRnR6TZ2FRmu1pahvxwI2IwmTLXYLJmmmH
w9h0QZB0wXP4uz2ocYxAaenynV8blbRHIk92SCOoa9VG+tQCE2oShWRGnrzYbMXz
dj/v5Bb61SOidYpCRWWttMqVUtDJkjUpDkYoWfpcZmAfh5zJ/cXJ50aqkdCs0q99
abc0peOF7lRBBYbF3CIo5te6L/ER2vJwyt0SD5miEgyJguY0FB0ErG9HTfbGBtI7
0KBRvrI43oiHD/UG340Sh1ltS5xl+GGdusgC9HA+OzW3nQQ+pVQtHvZph1tnzFbs
79gIE0YHuZBGP4vZxpVbw9U0rMqf4+tc/df+DeOYyux4VuIBf4dvD34n9Je+GGXN
qeZg1JZu0VZupy2dfsTXcMqKvxjvHoJiMn6oxWfc8aB7HVBGp1vXVlMW4GEX5Vwq
aEWKQ6iIzVz/GB0DW9RqiQFRDJLtB1LAHO0OSGg8LyVjzWAqsJMoXgfYbrL+Qx/A
U6wEW8/pyBqkCIEZDGAzvWsXdotuZY4NSIxb4jMOvEK26mQ4976fYBJTOuSLRmHX
vGpNSb+W+hc6U2Q2VS0TpXv9N4/8FZXvy1Wj+KQ9cqJoobHUxF/HfxtnTBFl/9W+
QUj2vdF3nLRHVHEZwnGN6in2Nv/B0Q39ZvZWASvenmFqHHad2diPfqz5t3af1GlS
28CNXtY+8VfNa76beFBpDGSt3TMIxIgK9yw9N603pHOnq7MU6btVir0TQGmhf5Db
0sfdIpmAJDsVbB7q9/WLNbmUKvLcnosjjmKOU+pJ8FcdmNFtlT1Xo8MOmp7KCFwq
K8Nk7FZKV7n3ZkuLHUJzFMy3Iwment6UTnHl+JwNe7hpFBJWLkonFm2Finkm5rgr
XI5BXTQ01OsAWKGLx8f6OtYlJAkgpZg8m6Ncl7+A7zwjeNYifGimS8MKZ7YJagh1
jmLP6QLKCFRBF3qg9ygCO/5fWjKbLIAn3+TvsSKs4WkbLFFhWOVjbiE2vgqJI6I1
E2fAT04rf/kqlziwX9bqJDIfKIqvZjdFH80E7xaYXBhZRVCi7jr36A1Yy6ES0vmp
4RZcsc2F1GxiQVYVH2+JcF2ALAm9w/fMO5Nt7AkBEZHNYUDUPXU2NPZZdTlxQC9M
tnEKXkU0NpJItAGLbHpcrlmCkRjjwHz3GGyHLniAu6xHHtzqx0Ir5RE27IqlkOy+
GIRWItTPgcYDQa4oOg+pThXfogp7BMeKNlD3g8dhqB5pQYjA6gdwenaq2XxmUDbq
1X0kFQPvMKZNfphIlYUF+rn492W+ZubgZ0m3wEa5lR8rY7eeFbgBlJTZxwk3HrLR
hP04YHXWSMoQ597hwJpM+RV54N4V3bmiYqaLLXY94EhAbVjQmC+/vDdQoDt125ba
+/b/iqhH1xjwNrtqmMAss0cSasF8cgod40vA3KfVULKF3MQm1jN/o/ziYXBghjzC
++rGjHh14tTNWk3vQ61ZQAFrjfk0J5LYRT8YaNZYqycKdIJ+osV42/7tnKsh7xRe
NjeVyofn9smO3q2hxsWFx4Y3LV+1EIu8RQ+T/XIZAZd0mQhazTxSHXM4FJ8RC1qI
8cvRtoWsUEHAqBieHu9eLqdOfhnMF/w529tQpSx1dIDctpSS0sluQbUZ63ziX/MC
XUGxRsUaDUsnCTfwugE+LDMTWmIIgJsHIRyzuvQzwWbVvf2DKVrB/hQC1KKqXU9u
pUEz1+Gg3LiI8h7cBH80BuQLqSV2Lxg2iGEf2n/bgS2yslt4c3pXfoeQnnYcupTE
Boizuw+IbpGOY76FMKA91//fq0zJdRRyot7OhnkLzX/XPazNNg1OuG4hToLxJq+N
NxhicrLH/qjQ93VZxXFh0NfWeSgITLqVCHwTWpgGZbZ4SoDiyfM9JsRx9V4AOC4P
FIG6bZL45Zn4QRhHr6XzrDb51YRDD23bEmQQ/12+sTVW8o9l3HiF6fXYV8K0clTY
tZpkyF0Wdi/ia8p0KennQy/lNI/7a18WuT0mIYlhSSeCho9JqcDA/bNqGqPZhNLf
3lh4pXzthgpiAQPCZMWAS4EaKtUZU1F1idbFBnMHmPF6WbmDN1pWR/F6+KUoxjBO
lPD6rGxFOmOlkW6F5yYM6ebhCLy0NLc3wZZqAeLmGFup5qbbRoTPJah2zG9me251
kohNb1+QTTSgfFMMe8SRzKmdQy8LJgiKa+ijaEY4jQaeuasc7O/peEM6kTHfp+dJ
DfEpXe4gpGzrMRVIbyFQOMVEEIl5F91vaLtQ1heGV7fz/J/S1MR4VgWnhTAGLnYR
krsXm6jjdSLnatTprIrtjz79/jDWuarNKRGj3TEYszHf9iUbsh6YSnECTuYG1gf6
pkpuF2RXmFIQlZXlfsObCHX0/gjD8WyZzRwfH8zadivoLdMQEBuEIsHi3vXyB+ia
UN4qH8BCgAJHt6ubc4glOysV4n9B7IEBbDtRzwENSFbynbnggVrWyj4K+kUxgKFf
Qx+YlTk57PpLDHoKv/2kHmPwC6Fqe0bc2Hbu5Kd+mCP+DGwTyfk3tweKfOYySyD7
JpJZwiRxtSooTLZ/QDQpffnYdq4RefC9tYi0bVPOUo9rD1DRKTOlguzNPoCit7IZ
SW38rVlriN/WSwUPBt+xazgPB/RN/i+aPxYs1FQh2PV+P3gp+Q9+4wNwO7bSxSFQ
O9DCjdqV/+hwk8V/D7G3514MavkstI7DWklvvN+6yAYyMu4pKG/kQsjRA7BNQ9/i
yThUi/H2CBQwGhnJy/YfMjIWa5coj/uht6KXK2/Ukc8i3Or+YwB1ZkXbhVxJBXCT
TN3V6t6n5cE+R5zppScwLLUA/Ayu288Xk+jGNdOoxXokFuabGZmG5C2O5jwF2H+7
8zOb7FfozN8kmhmy9wY6AduKnOX5jkM5ylatmzNZnLxNumb3ptourYsVlE6x9a8s
WKIXoIvL2gfOJNYQ6AXY6k9MHQibEaWHmoU0yyshjofmM3/mRhPMiYrOFs3Jq9C5
713WK55VQ/PyNW+sz7IP7nBjRJNBLNrcK3XtuW355QVM/2eqLKm+fGAZ/Y6fKtPa
G8y9oRDgl8SO/5f5Nq7Ukkxz4qaxc0UN7MoN9KPyrm3kOddPGnH8/7IqdxXr5++J
cHybT6jHaLceCwTJKDP5x0PCZIsgE3lnIvp9Uu5OAxIH+v7YelROdm1SQygPvePM
38NPzYn1EG72PXnKdmfk/HKm6Mf4K3+Y86OE1X7gaJPWe80pzTemDQXwwImh4tRJ
Ssluwz94g9ORDtvhfvNOFW4HnXzrnFTGRtR6IamUQ3pPtOckWwHdkMuV9Tw+dvDO
A+h7ffiIvVCfVRy0XGOZ3mMdaCkDVTQtZmrzTZYLFghpmZpqaG5stWdR+UtHccGQ
OrEytjoXVs4/dzUf0ydk2t3buhjNWS3m29I/oNerUuQGgOAtAZGWlSdC27a6lPag
kprRmd2u0Ew49g0xavcknhgE19B1FMc8eWOpgu/BnIdWIR7YQpL1Ps3f4A55CLlb
O9g0V3lxR1Rq1j3YXRMA0mUMl0Ijwpj7pS++Ns+U/ySV6MsBgYzyIAc6zqnAVqb/
HXUdzuCmxq7UezFdkCi+On6EIKrCCNUQ46/CjHCceAa+tqP2QTY1XUOIw3M+MdEb
63HH4rj1WzumzOYvKdK8QInxhEk9H5LOfjkmy9QuVL3uIaFUPT3R8kUjzntP4nIB
mScnfs07WkZmcf6XJ99ubsXCFUNa36pRzwv0E5ZnNmK/Nxk+xhv5ZQAJ3kwDFYJe
b+faamiC+5/6rLiCeigNHqAXclCQCOYbVYVww71LWRxKiT+XPZTKUzair8r55ppa
Q3x0pb8PnJOPyHlQi7fdH7ZOIACYuyrafVQL1olU8Okb9jaFS0OpeG0ruXSgkWpJ
iQR67OHd8OCwJdHooSlk7whWT/R0K2IBCQvhUv7ai4r+ueu8WKYeAoI6oTlwrUNP
VJEm/WKUwDXefAmdZwozUizGBIJul14YfIyZmdhMMLz8sBrH7YH6OG1Om8HNjqKZ
F71Wh9Ts9JSMDsah94ZNmln3lLFlYYwmkoVPtfYyanaQqiFZe7S6R4MAqeKVrjlO
HBcpPqMCdnrJ1BMS0L5FVy2dYLV8Rlds2WIy5GFBDrMW8WKohVHB1FFHrZYyXjEc
Gj6MDvbQXSgyfwRc8xUExx8pCMSAIwcczsKGw0YpwY4Jhjn0lrUUZrOSwyP0nsuc
ieYhNZEh+c30/1gZRqEoWyAultl7tcZtPCGAKqtPaGKxs+za5sFUMjpvdQlP1+pL
x6ge+jgITPPuSq/eAlwZeIXj+oZGVXqpn3A7GZUsURP8dJhSVTdE7TxybUeFT2hq
ZdYDoNaT7oCDZ/Glt8FclIfIeEOCpRTMcd1EEWMk4p+0O7007neSMeam4UgEs9uA
aMmsluTuSbljnGXlsQqsaW8MLR2tASJLNrsMb//JklkQjd9EX1JrPR6fcokefsLm
3/7+u+8QVTw/JRaCGNjLHaV6zWJpHSwBWsuELsOlCWUaEZYN6whw+AoZUE27/VAW
P9cpJZ9wEpBWGvEyZSs1EAyo3BJBCFpviWyV2fuOg+Pn9eAXkmPLUOKw7F6w7+t8
ZpXpa2CtsxoWr027jy6hQWJBfnUp0ODI8UDBNz+n1808eo2zDDjNAPqFNYwe6KiL
vBXW9p3N8ohBc6r0Lb+3sKIbpt3P+3wL9/N4WQnmLvY6beleQeMyRDUtVDWZlQm7
KzwxaDiUJoq5+2HvV16dg9gta3+UlbDhQt5bTySkY91gQK9iMcjOyyUTPjnLt9YO
HChdMqWv8aiIDgokRuJ4JZQ7HTQM+FjtM1+++GNSGMLIlq+OoGPugRlpQnd2YA97
S5PHOVYBNB/AIS14OsvzxWwso9xLL7c6HFfbjteq9dnLz3htbqm7SZYMrfFbvMPz
CIu2VyVpUTy9LZtqdMvrWyOKkwWOfJyv4fd5oIATyjQ96jp2NvdQl3jscJGn55Vm
TU5CIVCZ64a+AmXSrsYh9k01segNGbXzV51E2UeWA9pRitbVvtBvz0GTn3bCegP6
cE5/eVHdSqCixtORtgL+10bbrVLs11+ZxJdQCJjjUnz+krs9xbhVMIovd7EnB06h
MbjP8eyrB6t4Z31JOOSrU9uAYoZuXsvecKkVEU9S+4EA5rfQrP7xjoSGHdAzxTbp
TrGOJ7xKdhhElJmFo6URo8BmPpN4krDnUNBRM33zzR+FMMIKiFtiUp08DzlaKIcX
KC8MZVtnnBiuqe2N5EBuKySDRAiqppb/4eUaHYAIx2RcWiWmPMeyci4+J/K1zZ2r
w33FENkwyYGSx7wwjHgrncXCrgEdlfWDsp78QNV9Pfd70+rRcr1VVc+XCDcgjp5K
KJo9k26nfA2yMFoqVseAabDQ4cjCrStCqU+iimTBfQT6VwxSLknD+yl+bOZ+ZbGK
eZ6pmWiTd1966iWyhSGNsIOqb/EFqlsj/4bKrxveU8lxtGpEhD+lFJTmsERh+/g6
RUffaZ499zE+2O1u0dEAhfpI5ACyWuFZ61xxOyIx7UO7x/UX+gxEw8K/lMAv75PP
dyFRdhrYNbrnZN0a3ul8qgJjtSyHkjtJ50nIA4SOONKk1vymEaKCt/b+ZpvRp1yy
rJi8oh+QoLjhVNe1QKn/ZNhSeJ+zfocwArafehcZclmWyMDHG1cVBFjKSqF1CAJh
ls5ZiSQKVRq0rRmS1CJyDk7ReH8DpADvWEF7rIkAT6oEfxs/nDU85u4l+uIVsMTG
pIEY6IncKm5I6yTvcPrjDYjhi2VaaBHfa8GoLAHH3mC7WPUrSY3wQ1cGTvBzwgOd
Sq0est1KEY7NG1ztCMf8rhGA/MHX21W4q4zPgJsUSEDMsV/h8y8z1Gj3tOAX6gs3
71aUkmTEipGsVr2RqlW0np0Se3r3tAoji2b3/Y9KI1FJGcMhOLc5eFSeZQ31ULpj
sQtRBRpmib6YgBVwss9yFAjlO/z1j3hVyXMrTHV/7SMb1V5Mq8/1kE5QDkEByGTp
Dh8dmzjaZi6mZK6oMkwFpRCTMaCS+i3oJxJKGCo1yc8iCrQ1X6S6fmpVRyW5r+9L
nbXMBkZigCTC+xRRQ6YZuEXZ64uzJKpGpztX+7pV4gVmWijMyNhO5Kn+VJ/TR9wb
aQ8NFuJCx97Hmqk3qqPBvKY+LRAblCVXiXDiKKD3LVX8+rlKwwf3i7/yXyFGchMN
YNkbw+yFPEOZ/YGYoVccIQAqc2tdOMMWTqxiwcMrjZfN4gkPy51HCPdESj+nwQZi
xz9Uw5rcpKTJp87jFntzqL8cTpuNkaH62Pwt9wxFw8eaFXqKnVO47nBHfBkEtpen
4wG9UJGWPiuCwGlX3u+xObxVlvX2HpKpoqrrrEhrgFjngAeQ5QAGNqYdTFcJmDEq
FyhA38QON9/nKdss7gxODsGxyrafOCBeM6vC/tXnueRiExzgBH6Bco8BD8RGKWJd
Q/t2KOmkDL9xLsJVU9v8RYyRW3dhhNpkhvvn7Zhve/5PQ+5GcNmQFX9bKqr4Stns
Z+KwOYoG0rZlir3Xah+TN1VT5w9qBLEscbwuJ2Kg/aTmKJ5/Wvr7sGn3G6x5J8Ui
FeAgGBQx0cEKURPzmO3BfR8EGvYDC50tgOj6tNtX3jiZOo20VEecBZUq8WDBpv1W
6+5nkuIBE+ZY8786K/QyrlAD09DsQzVfkAIM5Amym4aZ1Bzv3ZjZU78GEa4Yb50P
IPf+G7iocLhSGqbuXehzSCVveLKbnRLApCgf/DZWwnrMOZtJPKBs0f8fZW/kGHKc
KwPodkAbPT8DC95TYRZlqYYFrCf5XzW67P69s2/uBJmhdn8b0aOXJaoQZDQ8ZEdR
v6v5ay2t4XOcb3iLS3atSx3pxMtX6oAtFU9too9xqelnc9/ZcqC5QPK72D0EFjhd
CQd0tthpvkz2n+4Ac9kIduByOrsIDCo87ax2cysQ+VJz4rE7V3uvbNqGrHm7kxes
5I7VzfuEZjdCwTUrEcNwrTYJn2ubFOSa7iv7qSH/EH1LNkxhlwJq4QEa9sKRJdm4
4Lsk9WUn0IphJyGbSrQFa8hVnsiJq1yhVeArP8O6O6ApFz1hSLe9CRdEVXNbpodT
jCLllVxWCPsl1ov2+Pm/G2UkJlcPhWGX5jUKDk8Oc3AQdKLUE0tNpj1Y2v/0VOfq
Hyieo2vPQKSwoVsZPj+t1MkWpjq9RML3SOXMZzhJTDHOk7eE4vXIOBdlFH+5k5P0
e9mVjtsgvTsPM+vE1aIqoiSBmUCkWIqtSJmaxiKeP/o3J2m8BQ1+M7qQgbKqaZGu
Ke5GIOUIonNwGS6OKHVLs8curYLjGyy/HvbE69M6Qi5aODrZpLHOV5BBXSzWXkBE
G9TYVYBJrCuOCZRoZpjDOUzXiMyH11TTMr8/jKyV7w2nOhnTYPk1Nwvk8FwXxTzM
0fCstt4vu4+J6dUNp95sY6IU24uFRFtzmtkeFU/ffJHvuWyoy+qqFWb3d7ApCjUz
6dcT+3vsPv4A0XpuyIgGhTUkPeQJajjy/F8er8CH4dUab4adI5zJfjXR77PUEKxe
bjxcdZsK44LMtEUAA43M1mb5hwMLE330pNFpG53K6lu6GAFUT14ldIIK5+ll03QE
tySVJY0dZiA1eTAOZoCpJKGCCsDNgVpMEUy7F5yvHV/36IXXTgTkc2ihI+JIMX/D
BDg5paTUL10gLbUKWIrYMwZqD44qcFpQOMKKCVmIu4digl53awBCHWaVh6sYZK6O
VEA20/ifdjCKPAlRt+18vVo43dYGZLIS9k9WKpvdnUx6LWGHRLssHscnyB1r1mTu
HKgftLPm2KCzUFso1bPPVRWzTJa5FU9QOdNJAlw2GajN5oqAFyEYpfJqpPfA7atz
E+xfJR4mXxNRf4u5QzW1DHJngY4lB/l6+/TSqtOsfMEb2Js1ixOzQnAr0yw1GdG2
IXLPxYeNQScGWJVtsPBdL5z9g6QmAVcAm0EL0Rul45a+HeUAfUt0ocHLmEHa+HXb
YCra6YdbRFi7x1zDCHgGZU8TRs9ts62gH3UiTG0pwQRaAWxwH3Ae8e3lyjw/nxyy
qjGznQwE27Z0zZ0xUy+hXtUFwUPpd6LRPZfkMr5YEIHeEAI+Zu63ZDC3648wkZAH
Ve2bE5/RAprywxCw7AMbapDX5gMu5/gsXhoftL/tPvNcliOMky2Jtbfyz8415JHK
XlRiyT5MRwcdgMurPMkhCF2YgL/2QzBQrQJvMtgeEZETdNVcL1r/WO4UhtUXwzyK
NtxoA+MpArryP+ye94XyDqJaL4yMkkdw1dPrBagzz0sRi0CyuKOKPF5YMZvURHur
00mRSwt+auwi+DMmivTCdsDSY51y4m2Wb6zDEpInzg6Mi4Ie4gx3tM7af/T10Dpg
wB7GcGq5HBERYK8rMx4XRuSsybRGyVtpJUwLpFlPMfx+P0t2vT0I6igGGLywoV41
fAmjb+ieqkcvD0w3TBlHTnW3pmRbPITrO5O8d45RNC3eSEDSXIWhE/NytqGWoiIP
YHoXxnDAulc2ti/gVfNUSwy8Q2KoWJtdzN7k0GEXCGOvx/nCS1fBy9mArRLfvHts
Q3278PeAwVqw0XQvW6DwUwuVPJtZVdLxGSZgmDrADtW8+jK3UG5I5RrIYydeDgg6
1hTw4+jhWYy9RzDFuZYkpHhU8BnTp7o4GqfXEyc8wo1RJ9GysD8ObIkBbXBZy+j6
VU9CnEjJGdFrSlYgEvaHKwYtj1yuRuHcJ0ph974dT9riXoGklKd6zEHt5Ga0OXdW
KmDul2jnrqbWwn2UWNTxr4Xjxh9axFaLRhi0DQtIflA/eemeHkk34shMFRG22YJf
iiHzH/I7/WakPxulK6/QlK69tocnCnJRYqnlt6zDOFjb9E+4c7iLb9oF/60cD9cb
uD3uvoJVTrcT3hSMOiv9VuoWJ8Og6qTSJ9ZBp0StIfyWC5HGD8OValEUmDOg95cO
tel2hudP7SgdK5VvUYkGwKH6pcVuwFm0QgQnlpreKwpe6K3Wwz5uSAlPXQ77vYQW
AzX91T3JrjlN3TXf6B643nv2U08qlNBr9upczHMX9naLPHZW/ozSXeWSJXaeys5s
EDPrjMYmxtrG+Ma3uv/b315o/vkup2t1UVNr4MGulUgo2ZB+lJDYFDCpZnBFh/Ip
223fb7tu490Rd025uzs3OYdUvKstox7gEz/qssu31ha58cOzchkjw+mKQz3EtOsw
2Eh3SSbABP/8zeqKgIE1BO6O96TjfnOMRlzutHq2Tjti8BsqEpPdiTSRpeScnbeG
QDbEs5q8XsSEDtBrliKe/CofoglTnbYWl9MtpL/HS/AmNterjgdvsrCd6hoxD4ua
e9oiRXkyNtQ7TsnVaaUMMYkWWvhfoFp+T5RP0Kz9yyy+jKG7bSYX41ymBbY1GPF1
gPGH5ShQyk72CmtYNlbXYpov/EkgSMJP5d2xbkdNnzuxqRYGVP6gQq06FP2lmHqn
IqYcqO/m9gAZ9SmcULXW4W5+nK4M16zNKTCE5zxcM+46DmzZxQ9sy/KKrbT/65f+
JI4+5gObZf/jrLys2oiBfrEiWQhr4X8CArhDFqavYH99/nh3IiO92KdXKQ8q3Z+y
l8M0HYClol08YIgX29vdRk60OZHxeQbm7fDA8PHrNgvnRMKK8uMwGk+CfXzViNZV
1lOk1MZJvQIJaAJUTNeqPhQmX2NVtGf4TXnNEVcVqhhc+MbqDxYXdMrUR5UY7qZM
Zow6a9N+8RT9SjZleigUBRMBmP3Al46Tgyv+w1smth/sD2uDq4xRAs3uSJEJumaL
qBl0UZg6SjqKMXGs1rwmgBIj69YU5PyDP3pKEq/wzIRlesDf9z2SkMxW2jM4ZRqa
OY2oGVmpM3jIpGGMO5xCZ4DnCxMPRJ2sfB/Sje34DbYXGjlRTv3mExdG8QvARWxs
Ze7RC07XXN/BdVoxMGbNHyQ6b0+qiVWLHX4sl0oDK7CUzmQZjY3WdhNBBODJPUB5
uuXaY9msoI83v6FdgTrrwnyAJ9MMR4UFxnHpyRLC//FVc+4lz8OUGNjeB/GFARrU
uL3DdUjfNfQlfHhmBB58SSdql+TE0KUgKqPaIs+eErKSlsVDe3ao2/QQav9tOGfM
yG19oBA0SQv09VEDHm9o3P8X5N8ZPE5sXHlDahdJdB/eKMHt1jW/EEiJ7DFWNj9f
IA6s/b5W5XcuhW2QYw80H+nQBlk9wVqLKNxo8wciKXnMTqoYgYhNYdLj6gkLWaNt
edUwv3ziWo/d5fmhrwyzU8j75r2Qa893gbrI5vqPb2y0U0onBSW8xzUmY0qmBa9c
77UHeuRl9Nm634PQBm6tcuNp15vZVxPTxmp+yE779jBTUrHAW5Uo48iaMKEDSI/c
2s3H1TVkLGeFN8yVYJkVApGYHzT6zHbPBZhioEryCbjapgrO5PDNq1UtVhpzwhdi
68+Yv9tEATWb+o1ts3eRv6dkJYEIzVaY7lNj9ItQEUsHeexolxnL71wD4nZpVz/p
/ap/RlWRg8YLtKzcM6Hd//O1FM+quYOaFTctn8GSEU2mUouRbji7DmSv4DEYv5BQ
jO8NAnhf38b96PzWzPSVk0Kcv5NQ/y5uTv8B0Bn+G+UbsTx4wi0KqAjQRitHuHV3
INXGGLMy643/F966d5nokyYX4D+tqJbr3BqF6rOZzOc0umK8+zTcVwU9TI15pxLe
2v/ktX1noh8Ygo3eaIfNzeY2sraHHsjKlD3IbznxfWZVd9pyIfBv0uSLxy9erUUQ
p2ZeDUBz5rvwWjnIlnphyI4vt9SV6Up5ptMMIMlaDMYEesHA9kJAgP6B1IMey/3Y
+AcrZHEQ0fZNjTfNIOArtnrCjLxSIBfxUgi3T4y6o7RjwDWBN5lalKtci4cW1kRj
VR6xQBT6UAzMUOYyW4r6fJrYQNH7eAkyJZhl4zy/aEQidhzdGfHvTpfApJJSdry7
pGUptXCfGxsAoJ+Bc73UuNK6fFolvPziAQDwXu4lsoWPsS1Q777vNnuglyP1omrC
06SgPCman+uD+4ku40dg3sxoNF8CCFLjWb3Khrk/tmYR+31H9hXV+8DyF1zfn7Et
fka+pw2qNqKf5oPyRlFse9gFsIjWCmjdx7C8vP2O2Hb2NbfkGifX2DTwVyfOu1B8
PBSvjYJmyTu1CMF35Styjan8BABiHBeHOP5PZNe15/OniNsmFYQnUccaplHPxHED
pCbUzhpaGslF0sTVkuHdBGUowyPtk7rrmZZmrISn0ZdtTLkXYng1rOQwm4ZDUKsb
w+/2rM/M7OM0GNMk4GWGszfj2g76SgLifQIMMu8XmHcSysyqsB6fSA8KjzIDENuf
6isGwolMzpBe1x9+X2ILSFliNv45812ojVkpu7VHZu1zpezhEKIjEn6nzRr83zbK
iel4K7rCad9iDn6+n9uf6qiApsU62ZkGoG29+Ey83AqmSpOUOANJyTSoN/7Vcxud
XUN1weBKrgHF8OAv23gu9N2zDSK8r1dbEV75ZPpqrGnqcFzRI3sCuwuKjnMSMpVE
8Zc44TvBvgeEftSoTpZDRlylSqhAPJOBiND8mN1svRq4ng2IK7X54wF5k3DLIhDP
MmQH3EOHeQpndaDTFyU8O9fQSnLmXhKsPS3rq2l/tuM5KLKVhXmrmMyDWHM+fBfy
mSmdEey9YNwCEUm9R2K3ONhViXljlJihGU4bswWuRsR/1WIrx2iVqzwssJrgkQEg
EiHA+JLl/BVpANrPIT1k9QL1Js1vB1f2lECNZfVZXOiEd1PqHz6NzNQLjzIM/NqR
rS8b6GdTfsP4mKkdy3ls330v+E8J0RtnlIAwOqubkO82g9ilaprKCTxhPArOwl1u
viHuTI4gskBB53b7UNvJ930iwSBo7CXZ4oJwgtZYWIVi0DU5IPHJxRGcuO24TnZ8
Y0l49FzLkBzJIWxCYGz/naiR4JdaGSj/cu6j+1rkeMBZb9W15wTc9CIcD5p6Hfd5
20Gx0RylmK153BAW0P28Jum8wZzrxzB9cekXiVpXbxEZLsL3lMg1iU4A8rND0Ixh
Z7BGkXbewijPfWrtyw9W58OBt0vUaUrXeh/UimnZt7io0z4eJdVV7NO9uHkrc3/0
h9lwQ0cF5iLSYR5Qh6mKSCewGUrcoWUzY5b+AoLhligHeZ1gjUH1cqc1HkHRLa33
xrsg6zPtC1igFc5RfjYaFXSKVpF2CEiD5j/+aDUBy2rNADBHyILOwl2hwBp6MZ9y
QAaJLeBKzi4+DCm6UAskdC7qR67y5ttyFxOmKN7I4g/a7Mh4HE+xbSHptRJt19EZ
DCu6fKr3tlctIixljqQyU7gsKS4/50tENwHaRkHrPVDa9WLP9XrvyRy5L+Sy4wPQ
dX57PTwOTpB8A7mVQyVxu7vsZXHoRRCILulR2+UwfIrb9YnaaM//mpJ1T6E8b8wv
T+Oh4un0cOkIpJtqysR+xEu+xZCv7eS2i6KQYy9fiYIt1JjR8ta1qM86n5rgANlK
oCjln59+7zjLi/yufxOB8Jh37wQvSmVWG6lsBxWhOVtVj4GAQzWdgMLK+4GvRheO
pQFYxWfltBCQWPzMZQjP9t2kd+TB7Wwd8438UNCVP8T1ufqPbnK/alFjWJxvWDtd
h0Et5vspm7aoeSGtmLIEiNflxx792DIZehLKWsBVQV5TGhYnLbZmU0RU70FCVIBK
GSvm4MzC6z/Mm7kGXoS7MUnim4ZqyJzpaVARSphVUkprcq6hIvaTCrYr42A3FRkE
xBVC0yuGOwWOvFfffMZpnsGh3LIuE4m1x5S5JjtCqTrNfuD6s5wRXGu7n0ssoHdy
r929gPzcvHuuvDz9IDISePGtliUcVaeXJ6bAw/0Yj//ABXLjz5dshsFT+pe+7Nb5
VE4WeB4pisq/4zT8zameorfHium380QdX2eLCacVgQOEFus/q/Sp7TiwXx215TBG
Vm6gNywd0ztgxefhm73z9/VGGUAHYxudUHKorlTx9jjDVVTZa1HmTIXO/zkhm8vN
DaL3tuvDpEHHjeeDiHiLm1olSEGbybxdyRO8fVmZAAaxIB480ak5l7huoHNKAj43
Olgn3uwxEkEei0kYBCVuhmbPdJ2dGHC6xc++qctwkdz/11eKdjhiYzQaF2ItrsWn
t+UaiD12id7JcLN/JZ844Ngp/LNEYHT7fWC3BB7EYXgPHQzIfd9DEJYQlTDMUuoA
34rsKeuGEIad56KLPXQog82BaTJ2kQRLyAX39QVK/gGV8OjRKIl9BO2HxPg8k5Wr
pdC6r6EgUmWZFHlSohK1sXwLcw8mrlK0Xl7PzjaEKuRhWK/pHDmkzRngQTPToDg0
6jNqz4ZoCbdg1kZoCd0WP0uNuz16bgueixU1BZrkYZl09EhYAAGb6pOzSfL1wTYw
/5eXxroc16sZPrwTZUnU4FGeaT3acPB/pG/9sbX5V2uxbPNWppQJOuYzuhctMrTH
lmhNAu1GCm9i0vyGfXyEVmnm9QpSdhQd403vVni1cBDjxCF84IoHj0VJBJcit6T7
JeA62rG97b8jizeUs9lr4fgss2mihzDdDsfp/RHkB+ngMHOzcDR3TulCMpSDQJC4
uUfOU5sgcfrLseTi8dp58xQ5u6Oa5KAkT3GpsXS/0uoyCz5/hodZlEhz4YD3XuUh
cGto/qfvJSif0MkK0DX/D6f1av+ueIAqiUGHJHHFDHv7yxOt600Rr29P3kcX66ys
ndGp7s9+vWUrl5Qt+HPGoDAl/KXiioRoakDRMPnvrPCBlSrXdXlOgufqsEPUnZLO
1lOkauID1b5cxRpkWspQU8Ht2IBG1ONq0nUXyY2H6GzNFAEskoftCbU5R9FQu8P7
RsCEZA1D1gruymvZnths/K9goTenQqgieOm1Nv26cZk4FzZuXK+krFWk2RB7asVb
qi0GaWva2fDRoEdi5gpYU7fkL3muO9JIEE8k8ZcsOu4CA3zECLTK8mONH9KR+CbG
5INWLUS3B2L2hcs8C0L5SBg6/TgziSSHmJYcWr410p9H8HcfwxjKF3q2yhTEi875
ivx5Rurwdb7hs6r02zqx270rMQMha97hN319TRikiLOjJqAKbIreJ5FoLKLLoXYg
5ywXgiHN9C1V2qJ7tdAJO3aYSXCzqetKdaHq/G/k2yrF1Sb5oacmVXE5jEWQEd7I
CIyGtoVnZTbhFKj33Nxys6DZKZZ7++r8tUUu7dFFlitmapdd2+ORaQKRgd0zPEjI
Ga0U5MB4dQ9nHkz58+DF7RS9wHqibuJ1X435AlWVoNwTgUys4GBIwYpFKXRFho4i
cuiVda22RqZvkzgxfO5tkaWbzge4o/M0wAniqfBeIVIiCeGpADv+OSV5nkZwmy3x
mNSCfG6zPz6DrZBmz9zlvsuTZ0wHsbFDwjQa2wwvm5MieqiiQxeB6g2nTWbrlA1E
2RpH3jYUVan9v3+eKds4y+ERyxbHY/IVBHRJbOUQXGqrxqbDwAuR0q6ciItmO47o
5xB0vQEAP8/KmpG4eidzVO3OLFz1Xno81m9Jtz02IVY/kSLpVRHTe8+xLO3DUVV6
eGsJawwaDWGyuvLeYReVMloDq4A8wOZqAMX4mGmvF31go+uNpV7MFghFV+IQZbnF
8UwWt9S3k4eX/wOChCxKeTVTw6wOxceOqMcfs1ri4x3EnmuAD9bF3QMBZRzlWciF
ln+ojVYdCk6mWmjSugO2C2/AI3tYxiPxEF58x7fLlrD4z6eTDxD/DF6PNT069WhD
9NebGhH2LsL7Uk2OwqWQFasTpbXytIHctVCrUknVEuIN+96CtUGmB2iFGRV6Y0Q4
aclZWYiY26COx/Dvox72U0MtAvXa/jf5I2jIaJ7s0XHn5kf733kKGej5pohyP5k4
Ft32ecbCdIfvByVvJLxFo7v/wPiI6yFCYDCr4XdmH5aUaFp5/LeVkf/eyRjT3KID
XJYeYuxapFI1elFOTML7qz/suEwORsYG2WKSZ7wU3aAWKXu0s6QzR3AlwTWZxNS6
uDSJkvlx+BMrc/j1gXLxU8uVAK3VqMe6svNLiN+Yu5P1cEB05be/PyIAnPJm179B
W/YkDVhwrGxfv0DNnovtkPSrHQJWIjbgseKXotH9eW9In8C5kCalaRV1KeoGhO1U
ekMfEBd0pEg2SA4PE1i5tvZvtBajNHCyaC91QMcXDwO1gU8HLwompNZcwq4fksE/
ykpzF5oJhexTkFVNReCgEPRNxJqBbuVnGEXtL2dnB9Omp40aA1cuZTigvY9LNGBR
weoYnbc138CJdIB3pXfpH9vr6xSExEPbtHnxDvDn23epNM0UfEaDt2ra8XqUs8EM
XTzxSWFbBZDZR4A8eH22GLqhsEf5e7ayrPrRy4XuUokwQqqWXpxXEvd5ah5kXUQp
WlxCRRnHqitLGMbTeIzlx+GImAFu0UkuSQ64l3cpffCfgmfKtLkxKCpdgNef9v4W
TOeSQNwp45UVHujdqGUBHO3EMUjBezsEhNgCgp5RjOzxi0lbwXM0n6U03ceB43a9
FkrR6SSK18d2Vh6oIEnsLgREPFqPO1AAKoBRiszYs74vt3zJneMopmHdQpzt4dQe
pI4XylN+uoLebOE/FjkFx7Ix0mSRe1voWNlur1PZmZr91sso4/9c4CUoKOw/7qv5
MNX66euO7DN2S2tdXLIm4pZE0H4Jckt8XprU46xwl8VZheUHVEakkp7g1YQe+FhM
Qvv/WoZSP8wqAMfagiXXqfXI4D3C6nMeLJgtFPVJ8Z/qn+f1AYWlPgB3iomL0XL7
uWUUcWiJKSMKckbGfOoaS3X6sc5WVVojIM+98lU50SjyqRKI/ImWkD6DogEuoD3I
IFT7CK6KNcxNlwnVjMMHp3ebrvsxNKJ/anaVFNjgpE+pQOR+Z/xE3sV1xSXl8xFs
NTsTlU3eZTPwMa7lUMH+fDO2HLPz3t7rmDuIUoF9MW4xqnDr1e1+opthUAToaR85
Zd5Zv1zHbb6edegg9PSioo5vKhsI5+fimwo+AOAHimjafnbPJp5P5KmXHcVNrmdU
IGdGN6C5GjA1sGVRj/WHHIVmNoE0F1OS9Ij/of7cNcAWW4dm884O6BGXuhiqMXRC
utMexasSTQOWE1PmHwn/mzTG7+kg67b9aPlZCPuKarMTqcdbDupK90KzyF83qBOX
12lss6OPfN14jNkbvVkbaw3LNCKnLVS3n5ODsBedsQ3A9WmMuUvyG04WjowLxxn0
Pi1diaV80cxniovsqFHlO4PQpErG8X6DL6iVCMpLRmYYqUKqZTtxWBDX10BQqyiH
ITqgW2LzowgutVjsDfrxjA1zeq1DbbweoRyCeyypJMKXT76Thj6ITT56aZKvtI4Q
zypj9pfPERYJ4dx8a4oyJXVjVVWfuJIMutCQBCjaFSGpzpMBGIgrpi/jo/EpCeLx
sWj24IpgIyjnZzAlXVTcUkp3s/U9JkIhAPuEqz6todhqBKqGfVUeMjov16vc3LF5
Ay9gDiQ8Kmu8FrRxuX8H/IvPYVlyNuOVLvkICL2Y/ytjX1aQDq5BHo/4Yv2++x3t
6E11lTFCfbHk6zB+zCMIDsRBCtXA5o3wbvYwDUFJb6OIvbAEwerP/kXl7yPUQG5R
OLjE5OVlJa6c786XS7MjsMqCOcMp9yo/PtKouwC8cyLu2Fll9yctnWA163Pcr5Z5
A6qGs3e7AYmoRWXrY5yxOdwDWeD3oi3uJ+/LjoRWAe0pJlY/WZGnF7A+qHIoEoy5
fdjBTOFUolQ1Cxv8Ai39iXCcYydP4q1sxaub1kSHXM8WiFMjhyTNk7XgFTV6l5ZO
mJ92AU0EVqBkKgOwVU/TQjhcSahYgebeq09EIQ13D3DAeykyKdJLbCM05LRWuIU9
5c4V/xf370CORLxshaSVC5ASYC4JysClTSPdqI/ioL1EI5CV41Tvopbrz+85JQA7
kyLUB6vw6i7S46deK9mggyxrnWZ093VtRrSoPD9fGZZpBrYB0KSY1FsK3mPStqjd
Jc8nSPZKi7qpSucR6KpM6iBeFIUF+gp4gyOkAIVoPlNDPuz4xqYnAJXViQNK/L79
ykXcfKyQnu1M8LVqrgcDkenYWyekvazJ7tNSbXLghE3Wgum5zNn4SBbILafjPmak
KgoVt2dDoJp7e6g0ix1YThnduQi+Lza3qmgdaTfx7qJsgYoqIIoERTjeT8+EVZPR
GqLViCiLuOkDMMLvjmvbcpFwcDMBROgKURNx1733z+3V+4Di/WgqQRILzaonNbBc
X3gXXBCITFqYH74kjmZd5yTmw2nRTTtEdwIHCt6IqDnvw97/ANwKZd1+ouGBr2mY
LnjC+nBMnLUAy4k3YqGifRjOzYQMhpCrmevDqqd6otg7A3/B0V/KR3o2NKuqss+D
W2xtf6EgaMkUB0Qxwdst+8Tj6uWNffkBrnn3hyO+tutT0kUivBu1b34b7Y83spZg
NmgoKqFdIsdkpKXZXtVAVoJrfL/wuhsFYhQ9LpWM1KRZTTMo6EO3ffpqa7S20Imc
9cCp17WXbljKsyknm4nCmqKhVph6pSA9MUTqfmENlkYhTJK+0wiRsd2WPgZLGZzR
oaQJbS2wX4nza/G2cssK2BdFu4I1p0fC9N+02X/ct7uA/OkJe+kK9/oQgqcL+yyy
2NhOX4THsf2jYEDFyQKTpnV+KEl3R6qlZU5+8SAHtFB8cJu65bsq87TQXJuMUxHq
J4ALqgeSo4mwYO6ZVn8toHxOIaJYlErdhPHZAfNJOAnO+cVGUpc4Xhypsm27cQ8+
RwaFtEYKC98QrPmx/Ellk/yvGHARgvlZPEcXYQfE/F1QJj+G9ry/V8DErhTcRQCo
t3TB+QaeJROQHYX0HpTmOPK3hH4fFaLd9PJEfo086U9RFscwYiUFayK4LDgP1OeS
kn4SiGAYDoOWaEK6oEqywv0m7wZyGjexJeqoE/HKnBRt3Y7zzoNZrsVn/+lrOQY7
FZRJ8UBlwM2tFfYq5G813qnE/6jRydL3cGEglcOM55agsc5aHeOaCjVyBOiA9+2Q
vUaXs6yIgfzVwGIqD9oDz5WgPUDK7NgW8pYHyewUyVruuCiW9YF7b+wa6TthZEtX
Q41GRTZJBTtVJQiN0AWeXS1LyyFHN6zKTTdS11YDvnERgeQarF7DUq7AB75sqhis
HyhZ5QJ79Lv88ppzCPH+p5NH/WjZXSuPV1uIWBaBucdHlwFwDHrpPgRYzgDowF1n
lodMFbmePydMjkd53YjveCJwporc3mSeKurgDU8zCw0PRoSuyjtUgLPjIy/+c+v5
aa7emuaOgmYSwSqOW76DkYQ+9COM9P6YR6Utfb/A3BFb5kkmDM9XYVtVqosjxDQW
Rc/pa7+eqDvELE/Vkmi344rwjPyz8XWEbftHTTgmztknDnz1gU++QczFb0L5/7S+
J/bx6jiXyN6ZC/ZyiU5CkASIe7mhHg2Mr23rIWunoR9VqYui0sOSSis9LXGICxZ5
e2TsqwQiu8yTVm9D3vgT1OzwCifGSKWX9UL08auaAIzKC5zFhpVDpqZ6SmsDIqE8
f2sDyrv3N9I8yyye/GdLUXEMxywj2KgMTLqWQHPMN72oWDBHU4natt9KuoIgH+I/
u6u073RZgGJ9hppqg/qyZh7Jv5NfJwy4qANzHW0Cpiumw84ZlTxGqx5pucfb3x5Q
9elGJZCVvezrHtbQBXrhvwJffSi1JUPCmrwRqltgjOqNsg0LLuxo4zmJlylK6uXU
bmwXe+pKUnMxTrtEbjQ/lglGAupjm/ahgg0kpkqUNJTNWFofHiciIRwFDbflrYUX
3OT9hSPS1Dmnrn8G/LY7Clmezor6PRLx6cJYZkcL12MB8jdlTzvPJv2l7gGkD8Yj
WwP9COEbTcROvJT3SgaFTgwZDPy88bnkZKNgY6qtwkrYzCxWaXt2ZboHvgbQUsjE
6ofClymu9etuEMR7u72/RgVwxkLeiE3AbY1Atxwi7RYTj9Unfhwl/6Cq28pQwRxK
e/Gltvi7AKfA5QI1yiMfiRC4UCyPAaRkAnufsAF5AkZ69N+jLaptpi0kY5YP8/Qn
79X7m3hoSwAEEl9NP2WdkXEBDlxYZTgS760+9sczckZiiKDKMg7fFYlAMMzo4MQ2
EmD9R2sax2p1WGPlnYxH+cJyR4V8OKL4DEFC1aO5zkrtD0zonFCki5BCXs393i0s
ahC4BGzT6QV+Y7y7lp1gbSknmrFtp67cUFcllkkV/gS9RpaTmCmvKZ/08jLq20GK
yywc7EuRZlpGEnopH52PckF3U2Cy9opxtDAuJ7sRPy2evcYaUfmDpMQAwgaZMKaG
aWCWadjhh72nHc19rwlcb5MlRqyjyjygtCGLxmmi0tzYnFEAoPzbMpjjjZuf6hQi
28CsLRjAeUl3pgbqKjFt5Y6MuwCGYIWLqcEuAOj9D5ZVIuhz9uzdNbXLHGyii8Wx
t/h8e2omWEscy4SC9bEitJ5RswSlBiTPhmO+RtnAEjfFVMutEh9zGkHIyWc7IJHj
jkTNlBrj30q6vb/Ny5U4J4ucq5SRPCympYynYTzQ3yEH/GSoiceer+aVhBn1fMTb
43UX6IA4d6UyBSfUdy9a6oVMYcMBMKIC3yITx+DujSLdzuIOy/G2B4AiRVEO5qbZ
bEouzS+c4xEVcOqeXuz0VuLyZhw/8Nwu5E1+jGKz1kl2x/yDexou/cx3G+Kagr2I
laIkf+kA5WVdrRQ4K/L4ucAvk7TEdcguRd9+zdDVqCiiDmOb1wWxn1eAAV04NLbI
ToJpHA3KPkJ+Fp5mBClIQeoUxO0urWgLqvFsTEbdX+T5thtdtOgxKCJDYC/fa4DP
gykR3p2wrlcKyGG1w87ekcNLlgCUmofpLGFOB/xdGHWOrYI3CBNV0VHFUeFQm1Ro
G50RdLzDLn+psIEEf5lDIR7s+d2F+g0PfddtBL/Y0h5FGjFs42AQHw36rD8YUOV3
jZRD2fF/B4xD89rCW8sa+GqdK5C7jS9mPmoZjpoPyjGRK+gif+S9oJ9to1DPSd8x
0sM783/S8F5Hgbr0oKsHyYhUTYDN/JpEaqbKMOuqf6gVR1Rz7oXvxzufMxzKUVOG
o4hnDR+ym/hnzVq6p0XwMQwaCb3lGQztk0n/rOuqKeJdeucsI7zGx+lGSKaoH/M4
FbdFEm4+7jpZBcgeFS3yhrK77hlP5XipT/ptivJWDf0mOzk4Ksi7e4R3p3XzG722
/0zqxBeqWtOuqUBrEWblUo9kkh7lXUn9l0qSRVx+0+4xpePiPBI2r9HMX6bqf0uV
BcNW/ip0KznEtzqCDgFLoMvIehBE0r5322CnixJmP1MpiL8LQmm+s8RbYpOplPHh
XXigvyx8Gqwnyc7TIFYDXza2Vh7kjbCTS4hXV4X4527r/nI/beD5xDcosDWxwW6S
j4XeunS68ytYqybjCld3AEqHnLiB7Jv6ZbyKP2EQ9nz8KH42+4bbWdLI7iZe5jTC
Wfa7CitF0QEoRTFHDpsSZXbYovRm8B+JkOdcjDhiEy0XSJmr6lIeUy84iG+343Au
ysXFV65+p59T0CebTYUMGJ09xHXWkR1tPaahrxZ0yE57asnK9lmOS+Yty5ydW4Ry
yh/rRWzPCXtRxpdEkLd062YG/+j4NoEa89xFCcSmB+GWOidXMC7ykvX/IhOEy3H1
arwFhe+0vyW/sDvqhRMS1iJ3ZPfYCtlmFJSNrskM7f+zxsrRZcMzREcWlnmZ2p3E
o5VuqqDtLNvNRPkGFWIebkGfj1Lo+b+p/dxWFGvLX/T121MVLOwwD/K5GXZhYtDR
JlBhoC7mCE841Up7tCIQ4jD+18qP4aZKdX0cpq2sdvU846nMJjwGMIoN6FWvXCm/
KPpg//4um4cmQ58wKvH2OWLjcLkxdohWiT6nTdYrDWXk6rUwZNs2Z0yY9ElWAXGJ
t6VCgf7KPnfUXkA2aGANp2+cgxpnoZlwyYBQVnhsr/hF1hSas//xVO27IJWtktcj
hOc58ryIwDVSX8xZwjTj1PKQST4rMN86lE8UHZ2L4FCv2aWGLkI5bjKmGvcYTThh
8U07am0CRWS32ucWm2D1H+iUSkjn4VvGWl0XnprJX7d28DH9lelF7RIIvTRaQFMW
q4nr7NlkYICxKE48ymNEzqDRXSDKrCiUgwfKQnmnCxzIeBAFwu6ENLHdF3zrJwVH
XVlZh97ETn2D2Pbq+FQRYH+l2PO+cpCUcj5mRSR+n143iWEqfcZEZDJ79zFqMe+e
S4B739qf6g24uGKeDKYGEihzzpdaJgEo4K/pRAo/On7YNk6Aro/AxWSFdOAWdUJZ
5S/Ml6Uyz5srcJ8MiWk9ZitgxYT9VAMsiQf986YsUssGJCRlxB5RAdrqf2pPf+U9
zyF6HlILg+kmFZtL0ifNl8AhgsTuQYU+H9SZ2OOd94l6l808PMpNGWlNI48T7i5u
JPqs8LA4LXTW2o3DJHTlCo2HzPusyKpdHrM27qtAI3gRiEU/J84x5n7CcqU3q+oA
EePr3wLdCMSOORgU8j+7yHL+A+e/RfpPtIeAh3GZ0UIOKwOrq2DtN6jrD9oCQXsh
Hc2DnR3MgROprG0jqY6pldlKm8wbiMatOGw9gwpGD7gHlDhBxUv5Gd/0Vk+7KEls
fyThdpYNY+KLWwImM6SN/gdmiHw/47HZ0kmGGj1uadH9WW/8jVctvDQbq3cmIVoG
RIeH7ncSIHOpte+i/698oM85BbAVlHN8va6gB4jUpIOuemIill0T6JFrC+w7eZib
vR6DCSS183AEERwPf2QhG6iIAbYsHzwSehPbTVrXmA8leasNEdi4hewi5tqxwDhk
aldihzDAv0BnuuuzHheX0sNoK7bJLfzr5HpWsN6cUNoCDweqrl6QJC7o8Ag6TUnw
SFiRCXawIrWF35ZaHQiEXWFphK17h2zg3MkF67TFBVGzSK64tXt2TBIN+cyBCrUA
Dmq0GIeevOMzJL69iqB6tFl5yCWjzC37pDM+VgCH22b2jl4cWQOMJs4v3RaG3u/M
KNLyVu1pDX3dVeqfgIZ+WLtYAM63vFXC+Xb+9t+wvjRPgIpb/ZLy+C+objm+xQs8
SdsTeqc+n/A/18xPcXNPk4il4+UwxFN7etmTmyw4R2+2RnJ7oqa4jgsUVjnchCfb
6y+gxAf5yEQ/o++OKEgF+yMDgEDH3NMD/bjIQ1U5mMogNXF2nkvMX9Rtobiozg7R
uzkRybk76Zay3yTAi1N67X6SKOLc8XNCLLVQrJ8ESgiwSR8Bacx43lV9QOLm34xK
5KerhslHGoW2Rkjd248IqVGkHSWd2m6neWFrVmFzCVqM0bHdrHBAUWFWLWqTVq69
SOL8Tnovv1tHTKCcZdHbM2rRUwaKIkVVCgKuN76sULgex6UDMyxb+HRwTpJv7P81
TS7H12yQU2y33SqOfDU4WGS5TplWTdPcL/5F5Kv2EZG8N4lDBTymcO8hzq5llEwy
hHUTBm4/Wdd+jG1/AB8i+y+M+bSwRuzFvApdHaVdLUotm1kujTgPPQwl8/TD7dOz
dH0EYW8Rr/5pR6744rGcpeHZVNxKpe/kAC6ohhtP34K2MPlnxQ87+F37TjmqGDBg
m3xje77s5XMpy2uKNIhLjts5ftnf6JwTLzkQAlzA8XRUo9ueUbNltT/suB85LLjh
3uXkNeko442fCuZ/ubTJb2KUOCsW2LvrtWm8rPdI+AEP4lJ3sUfkTxrOq09pdGdG
1cOmdh4l4b7jkUeMLVk7EC2jxe+UPREHCsqozeiwmqVqNN6X3SOHGI5851MjB0IR
/qGQtZH4vy/pZpyLuyWqZ3hUsXOBUBZypyJ+U1Da89aA20YjJ7zbPSiFr0B055r9
N+DgLtPAJblyZzKbBTru+SJMS3RkzTD0vH72CI3I7mOW10BUgU0d73yinwvwKglR
7o5Fddd+rDcFnYLQzeoQmvAtbBICvyQSOf411pp+NtRogTiwXkBji2jZ0Hxw/YoO
g4hO4Ux//qH3A7BkyztJOX02MFR6ooOSkQa3dmAiAJQ7vQ9MphM067fUtDwupyEV
or4x+DiiHhRK60tCmt3KpbFVF9PgXFJOqlQGazIXaIdCRR98R2pXrI/WKkQQkIp/
udNr7Lr8ueCwlpeG0LAM520xRHC3iNw/oXVGUg0Oo+/u2A0uUBYNCRQkcBvq+jiA
EHoubb5CbFUT6DF9X2iCOkvbAJRczU1UbYPW06zwIRckpeTebULVtlssuDMOEfGq
ixu5zGOx0uIzIW7hjg+kjp0Yq3cDxA/iwKGrtJWM+rvhsH3/KNdMxwgFOFn5YyhO
r5o+Dsrl2zeX1OEhpG+B//HbdWIdm8EFg4TDq0JJ4dCKDPM6izDBTy+SqJafp2po
zm3Lzf0eP8zcxSnHNWt0Mkb9vzRDy+/Ltrtbp/RdLIogqow1/MGPofMIXZWzP/ZO
gxnWrjz9qQ3URPZDVVjJ5EGWPdkC1J1TwlCWnAGMKV4Pq+2VxIFOBYD1IGphleqx
R7sewbnBzdgjND1H5lp6n5e7W/SLWbnqe6Bp8KUEIpoy+jJc4Qwf7uNhXnISwtd4
Yg04pbS0C7cVt2/B9mqD3alzUO/Cmz8glQI91MKLFeu+A7oZgKWemUY+3EkYEa7P
FdojVpKzF1IM648r76hq7u1gHXuWKXwGvCVbsF5MRAX01SMQZbidEdq6PYa0jEOf
jnAltTirZ7e5ZMGK3xnO9N/+I0XT0zp2JtQIaoEQRkYuz+GfpoLIfwKZ3FzCTjo7
SbWIZwswZF4h5Nv0FY0hQ7SS0e+um4f8bayZUSgKbvkOQAjsjew1pCLAiCAs+6r7
BTmmJGR/dPTowBMK0L9SwUkZTtN1kcZzhXDfIYP7+iUKE0r7WSkXEQnsVhp++lg0
hCCJPjScJTp/4LFpfx02APetb3//onerkL5ZBQH1Vcv0N74LCkvj/AaYx0ObEZcT
rakDG5bV8JGAWt/ouBlPufOJnmjhJ6RMU7CRAMtSW7hwK14cR4JrIbli0AZy5gIE
5JbCwKDdz9NEPaFFKPhNvnylBzdErsL2XDzY70o64LRr+vWMFM/Y1R3TViTje1f+
K2mwjuhZ0vJJSQN81vEdiXAHJzWyMvqOXrDvkbuyDA0R2TdtFvuox/VOm3go21Io
idBUZ9SF/pO39O27/gb+z8PrLSPAIKrsHrw5MrJU94LZTtgHhZlmlb5I1TF8DLdA
3U+LpZWv/CzN/uCt51wq3RT1D3FoQaZQ1rr0Vpa9A6UD7pqnYNV8j+eI/PwSWov9
4lWmhZQBNZ3+uhbonG6Xz5jXkDxU83TAUmOIoIOnIRz3+wsL+m7tsWsZh/t+p4He
EyiDLfEWWJKPC8IjzsjcjC0rjH7M1PuJiyWRiuXKF4tRWIL1OfRmJEliME5VgNwR
gLyRQnA3o9ohcC5BeTvTVBwxmBBmggSoRDniDtAPP6zqbg/uNqyM5Fp4Py8aPt4J
EOjDG6iR10/sa/xceSoJFInGGaUDzZyVcYUULCPKku4zZF35IkZ9tVErm9x3fGXu
pKXX0QYA9gYme0Fyjj5A0y0YF3YpLxaKJvuo04vtTNf1CJXpg1TZjPvMOO4DyOND
9i7E4UjAheLU78kdBei9M+a07hjL+SpYTZeWgAOaIQEa3yCduA4503OVfvrV3B1G
99+2jg6pYhXjP2EbXVpvpta36R2CEBGHG7sBDkcMpydhA8KL9891F+0xPahbviyB
Z/0N+Sy3TNZORUfiLpOhkpMiOCVPQ5U0NCerRUHk6+iF9PEL9i+TXDMQY0EfpiBn
Uv1jnKz20mzT2ZbPRIzM0/I1TaweHVErj4HYSbNIccFrYom8284x33FqK7Q37Q4r
ElKv0EseD50rgsxVFSNl95ibA4q7/21nE7aFzN30TO2JzWR0dMCYIv5EvZ2hGtcD
nlJCTOe3dRVt7K8b/5SFjwpl92XrPxQyaV4uVLRuYvyy3J4dmgpGBJx98C7qgxjB
x6eymCIKaGpt9uiNPjJn2pq9/4/LZrcy8NTNXSe/ZUG8UwclY1+ZDFKjNLXaR/fR
rov/5v9FZUUsTzFxKRxbafeNP/9LEtrr3Zpu45r+5zDdgfAmsDJRtMgEFKFrypP1
clKtJmInN3dlldZWhUmgFQRTcDgRBL+9+G1V7+gfJSU+EtBh1M2NqnyjjBvnfvRJ
ytT7xesfHRXcNOWjRPIftXHrkuxyTys+lyH6OIAh1Jf1y9gz6aJbSPCmLEBBSoto
XeGFCIqNCNuJ8BpyVaQPnapFi6boaqQTHTQQb7PMK/87ZUtLY4SZl0pF4dc9AkQ/
tV+MVuGkw01pv99BoN1xFVvnuXQeoykzoODwGl2DyiLp5vymhlE1BKXGbnyqH9oa
B9JA2EpMUx8D9Bha68DLEyx1S4G1zHVU/LR/LPd5JXW9nihNpo3sZqfnUyLJLoty
JZJZvj5MOVdJUIBQdbXoC7fOPL4vxoSOZI5R/iFKUMrUB0XDFCfQ5v7IXjtf1alj
U8N4fiG18YMqcd/qM2s2fLuG8R6Hh1dl1BoJUVfsW9uixR/d3K6rj/VyjvTz2hd6
QTyonkF3FWZBp2GHNCZxuCxBPq+TywHGlyhpH/iIRnH3gFdWGLVNFxA9isTUbA4Y
RT05dYoZn0IMzOsJSWkYa/+kd8v7EdcD0K2Q3Ep9VatVZzS/l3idvmY+aEGsTWQ9
QtiChSstIDsW9nQ0Oy1ay0ebti/Vra3fpWFAiH+xf4xIFElxePCLLzWULzaAKl1Z
zVD9v2vYyVMjwmGhcUFwyi1ipnH/ZBg4CIB+aA8EHsdtsWDMV9jvZMcipbryIKVY
vIEaHp6tOcjV3ZJ3zMotWhpUsHSKdsziy9QG/RqeqZXbEJRY6qlMepxudNmxZiyR
AbJZaeePxRa5Jd9dfXCuKt/w9iN/vvIdNtYUPuD8LM2FhPc7t8/9sHgxMd1OYAn0
hvhOGKvZjnW+qzftVqEHzhVbxjD31nxOrSAaimO60TmePUN4SlrWgUxSzX2eeJr8
eOgn3btqiwktExjmRzBK2vICCy9ng19fY5c+tQtgiANeXqvDrmKtAjyrZzfZ45BK
dQE+LVChi/tkB4nhKPDAvudQNDRyJs8NjVjJ1+GmfBFpMT6dskFI5NYiQgU1v05f
Rco7LYiYh4xRGkcmilCkoyTAHxOszUsjefVgwBXSJC44FhpVYFSmq3IEfde4AXgC
QfvbTYlknfyo6e5pUfHmuocoORL58ZNyBprvJu0mF0cVwkk1Nr4JvV3TuoSmxGf3
5Yh9aQe69w1RIICREhO3tmOUasVSc0MdsdZQitRG5yBSx5msQ/v9WWlIjl8GjC+U
HGqZWXqLPlVfIgZcKFV4qRXkyg5yK1NJqfCz/i1fFiqnW/fzRhcRPT6WRqZrEcwd
Z3MZPDgoamdGz8uY463nl1m77jw7Ds9ltJty8E0HbMLZGxsaqODmNo2zq1HwzrM7
aAuSjYV9MTnz8czspN+47ASYZfA5bUesu9okROqdR7LysXKyiATz7gIlJjQitktt
1DeBgvvRaeekLzMDCrCuEAekYhDSNRGrkearNlMcHeWzO+gS1koAAsfpSqmlJdQg
wTWDRF8rhzsQUp1CpfV2yHqxVgHuTcCYtRXfH0I1H76+adaZtChnSMNaRp9ryK7B
txCQXhKWkhsuUbwXAmzWVIvSUKVPGTSRc7v5k6pT56TH7PB/WyW7yh+TkgUzNoS1
zjSt/mX3oQtlTa8Dqr5r/uU9FXDZavvKvQnGuZEnFwE7OBQZ/6VJCl5MCuso0N7k
kKzBIK39ynKBu/ng4O+rqD3QQyRPsZVtFQyGlYZVHMDe9RZ864VVX7t23sxCs6+T
icaKdBp40cBAUQA/zKMHC8D20WS9DPdFULT9DRIt13YSkmV9Xrl1kHL430F0yDu0
INduZoVAD5UnCVwRU/R9/LxkUzuimvvepk+0Ms3nzBNH55wCnUT45Bdv62T4fKfd
rrOpAQ8rwcUWGzOpnK9/KdBLOgts0yz9euHRooPaVle/RiashbdKnZQs43Ue2W1T
ac5nqPmcRA91uIam8frOAh2Jo/E6L2BaTBmbfaNdBojZStUu4Qv1ynQT/exUU+vi
LhKyI2aKDkvZOkuHqVtF7qF/yolPHE2Lx4UCemdvNjuIsyuUhy0xp+XaYIUZDPTU
afOBsGntWWUKI5HljGh/4jAakSH/X071DHILCjvJ/s58E22thLZhedtaNb/muP8y
AzfQuqOgfrwyTdVjcSBQuesMUpBGn6SJJxNahnGnyh7a9m/YlNmat5arMrdxXfDu
yyGqjkT7oHYdTK1+MPQCCqBNW71Lrs5r4wdaOw6XGoZQv74Bo9LpRZ6B7dxR4kmm
F9xJr6VHPwe+iIwcPnSy9KEm2qi8BlNDMgYdTrVnOMkRM6Kd49BowlrPusi6Nvfp
pVRb6mpC/ww1LpGfZB61MaYd19YEHgRKeOZLX2b3/wERt3NasXHN+WDEwg9SnKHo
TAspfgILA0AD8/MvipTWN52ilRrjSAv53RGUvHaQff/6XugBL7c3n53SpA9xI/BR
hIQv7D/plkiuSspqfyhPZpOrQR4WsJNP+N8fqTs3schulsStnxeedVLLjSH3jrNT
9dX+DrJnjEEe9Ehc4cbLxES4Fot3DGNUMF+9YgYEm2C14CsQeFabdUrGFfbj4yI7
xcUI2KAGNBRrjhYV3oYa0kIti/7VsxIa5j9DAEEfGPYrHXzbIr1HFnCoxnRlmxO3
HcFierwVxGW7tyG9acdNEbEwZJf/OFuPkwz8YPocBdSwnJgydiprZd0KR3g3Fyw/
lI5kAOirTZdxPEONtpfkD87DL4JC12avlR7NQotkuVdByX6KO2MITS5gDLdKlbcn
ww4GNU5uOkktDHNucAeNJQWgIVQCrsbYYV/dewaVO1lwT400xL2wDCPI8mbAY50n
lxaf8ae4F3gqkFroIQZPhcny8BBGbTqBaqLm6CL+eSo+E6QU5WoiBexXWmCWtjGl
cfFwUZM2VDnYF2CVtQBUCqYIzpKubXsZQ5ecdgbS6QDSeOr17pDwdZD43peCc2Tg
0XlRZEfH0aCCjKuDXxOeSZT/skB7CYYYq5Z2iabExV2vFufo7CkYKIgJYu3wLMEE
wZF8zcWUGN1/iv9wcaphvAFsiczHchv3hOxmaX26BuB6vniJWIb9mDHrTS5vIs+1
DbnmuBw6mjZEMFPqKz1Rt4qBKzH+K26uqKF8QMdqTd8yTbla1mB+RjAmSxtui6BX
wx60uKt7bn2nT7z2jo6PoFN2cb+xvMWdwtSAW8bTzQqujHlNgn4F/SWyEP9iyDuJ
2PcIiMvci91ciO/U+qwzi+xQEkA/8M9gF297xDBsxoUWqjwwiVlMKWqTS3DO3s6x
zEfiDHlGqap9Biw30cEimLI25VsmBbTb4syIzqO4XsdcSIdp6oFJNTHZ411nqe/x
Fww1LShWQN9VnOXjbgXpMFk05AEUyj4v81gfODRvVY4dUmYpQza1pInsJC1cuUcL
vhNMK+HpamKo9M1QTNOxEborYaimlQ9eu2Gk12ES3zSb4pgDLZBl0CW6ZZBblY8J
W8Acfs+AWofkA2ByU5bGfJOpaYWK3iiOdnfbCkDFBUiDs42hQwkPC0wa4zmD/cSN
95MjkyaSEiq/trFeTC+6kPWX3/rC8gv0/7PzLFrathgkUcmSakYQtZ/DtwwEZXjV
/SYeqTRJQRwqWzI0SrBtz0CD0dockKnaZQtzSs/V8bo5Jnbx7Hl4Hiu6GUbZpVzq
LXuDo1q51IR8Ak9kLfwqdR6sqNAiUW6lRD2LLNqk7ZX13RxKm+6E6P+5GwQMdKDx
d/KVg5o4lcxrhUKLTeDNxSnHjC1zPGQ9Z3uC8hPsmjTiZVi5afQmE/BQEWCRZFon
FvPyOc03xaZEMm909Xip8ZoLxL9ZtvkQ1zWRIdO6POyzEtb7FJLeTbrqBKl0HaLO
PjD1imy/CrfOdbs+MvlzJD3aGNq96kyIz5oeE9SaeagzzCIhc9qZTZ2j7lsePB9u
5Bxo/Ti5O6NZo0+wsgmm1pAHlV8DhBGhF7EGVcK/TIRdItcA9ITdfbuSZu1YaFNX
2lCBMU1OsJcruc1vo+Rg1ChHiSwN6+uK3t58tgepF1kHwP7DdSp5NVZIGNGyyTiE
28PQYE9TSWCnvsFy6WorxbH5RvFpNm2+Y7dZeV8RhHy5SRUNK9hFbwB7nGKBBFF7
xSm2nDEbCmnTqH8AToNEXc+zLmLJhfWW1S36otxTWn9RXrBmVOJOUFHS+X+LCUKO
TLFs1bbf4Vh/pOr03+Ipvmvq/u830/F32AadDfGsEOtPa9gWJaSB3m1z8Lmvj5va
wCO4KYKLkmbeuFaxaIZ5HUxw/aOzxvg3SiJXkM6TcwD4LRx59tboATTXn2UtvA4G
4yORKXNmcEUNAoikKunh/WFR+RQl0feLSr900ueX3049fcqOL45fi1fFr30mQqGe
qQIbA3yxyzwALoh34x70+V+WmyIqfpTx/pJ8x0XT7Pvynwo3mQpeRLBw4sWKp7K4
G7wMxyBnhrt2VAwqWEZJvplRvG+GTZd0BDVSTZmCphVcGVxmZ6/97bnoyuoYTstf
EgDb9H3u5yRKHlUAr5AY+AiwvqSytyX3btqBGnYbVZcfqYGYOuMCImqyQJro4uUG
CFRpUFJv4vWYhuRGiWadg5sHuNLoTLAXIXucObR3aQ6XCBNRLbsBoQ7K1kuY9Eg6
5s55quVyKdyOc+D+ywHEK9bvsMD2XJpwWmai5PcXrBC/QxFuLSJuNQwaoYhY+WdR
xXpvzJ90tEGoU/hd3m7FRp+B5wDtYoTHDbF8JWF0WPgcR15IH7p/oSfLOesSaY1c
hf92HsNFg7IQcPPFcy7SIMq6YsaYwVsRoEwzztAQ0ApEBkuY/idbOHwW5ukO+XcH
r/5/r8FreLunH6f94MOVXQ2tU6/Fiec9J+NiWsi8Iw/ds3nxdfQqNT85m01N/WMY
s+TxuY/8gp+WdQBpVEWgSR594QzsfdEKQWK0DcP1PuI3DXYr8TTk+SKh/zBKb53X
zPt3o3FU8Xk5kqCLsHvs6Q0Jf6eK4XSlIEMdLDXeCzbTBBRMxz4vAWpjCjUraXzw
JTEW8fLgw6OJZEDBeB8YLiTwWQs1Mgo5wUW0Au9r6zFEdlf3naz+SNElsHZ4jEaJ
Czls9tgKXOj6fD9TGY2MqufY6dD+iL3Kkp9bus1+nHVIMYXjF3LCoIz92otgkrBt
/PyqnoTViIfN3JeSJTem2dVF28CywntrrqwpnyL4jeT1D0oS98Sap+af3WCxuwv3
TvpvUosGsy8sSWny5Bh0BrSCyqVLIcXifMB4/FM7kA2NJ0Rb5nlY/NJupawMPOpj
r2sPhoB5sMSXoPtkvsEodAIww1zV65GaJ8rKmMmDlWF86YxRtrsBYO4qlVf5GsI7
`protect end_protected