`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 2656 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/9huKRhRMtvnNqb3Z+UU7TahEoHV+T8U3P3ufru7l1O
3DlgtZzb9QxCbOjthp9+wDkjygH0eUfDrEl1ovhZG63IoSHBtF4u5nbYCqlrY/Y4
Hm2YmiRZSRWNFDkqJLfABSjr+vva8EXymGGlj77TIlZGwMMypcENf8GyFLAc78fo
RMHpVuexAqpDdbxGId3t7OOEu5yIomnnJeVgDXS/Ro2+DtyW4lRklKivB84x70Kj
O2DJy0otsIvGg1FzQb0V+SHIw3yVjpmXJ+R+PBW7LPX3vR2W3a8E7IehZVg4Q5b0
su2TPD2gdQGu83ikaF3bNPu66IYJnCp9CRmFXQcaRPixKhpZC8nuSiA3ThHtnIRT
NR3/onwYA6OFBRq+1RWq4+BVZdWuWyBCptbGkfyhyeYZ0cNi/stYNiKQuNzLgP0V
WDwJUNTiPVqk5BRASCh2AiHMEU8kyTAu8u4ISjnOGX/QBbc7GS73AamVXnTzyS4/
prmrioSLLhM0eDyfyuxJ3O+9VqCA3HwCG+xdR/ZU2BKTt1zVR06F8yyutqZNFOz3
Sowo5wLZesfaJkmj0CBVSXnLTw1NQUG6EO44uiE30DjqiLEzRtEHYYtgYJItEqU1
YueAXPwCHE/c4NWjFAqOyXGCsvKaTz76QLuCXwLt0AXB7WxAz1XocxLngDmo+NxB
tC6mrqFRnDPCTL5AHIj2DFiV74MMMmZeTR/BRiFH1Q2/z2thLfXbVnt3QlgDE35F
VbXmKE5ZsEuoegkQORbzCM9uHQvDXKJ2vNYQdex2wm3jMarDmqssnl2ZdJ5/HGQG
pNxJZYSQmOT37oH72FZv3bs90+tAYZRk+Py406YPLFzS7bk1IaW2bj60ssoIMNoK
7ixtjUddjB3OY5PGpwTvqMbddYSwnXrprAasCQyQ87v9ydFn0DiCurT2rMv0wvGf
qmWwRxA9OVXuHfCbCPpUp7stgmlz9n7mQ6Gmz1Df71ckaODbIoaEh/Ecuo9dsRiw
beNMf1XbrQFmYygbZxxqpILRKFJ7ASMUUCT70RoQc8CPEpxLX+5dRrMmx00+a7Hz
7mXU4jxnEoJUlD0Cl/4DbtFvXxCjBVrjT+Oy1cfpR3fv7j/bm2yBAENCquJ8Q+YH
PgvIUW6Mgm1Xoj/eTAc3nMd2Ez92df5VBPH0BkEZnUWi8xYVZ4Dvmx+JbqVkFFFC
UQcU9NXMbJWZaR1d1YUjshTmXNOXLzCZOZroOI+KNaytTwSaBXS80DaWvyBuPJPL
p65910J6rT78iDcBsWU6k2aj/kmm0aAu1IO/p0RSgo14MXy/GMNuBmPcVEh7qRlE
8RrnTjQLNYrLFdMK8a7Uod61K7fYdjpaxAd5MGLMgwHHcbD88gO+p2TnTpuBgSw8
b1PheAgx/J8R93J7Zr/QuD9XI5sAhwa/kjOpzr0SKAfKpoC680MI4kelHo6GteSS
w1FQNSOgDjhCXM1pW+guiDlAcAvqrRKg/oDj+aKMsm9gCR7lVDMGdzlGQ7aHiFZm
tgBDkl+Y51Ka0nx0FwgxWvawx5HwQIA44tEhzTpni54GRzWHY+XV3UEsBX+9FtRQ
rZUnyVNeQKqSMe09Mh5jsenwyGsFQB52F+jU+idY41pmhk7mOjK/sEaj836aKOuC
fJ5eACJzVRPH5LZAKvsK8WAszrgXX7vUCoQxg8eKr+R/jTnoYFO/9Iho9U3JqWYi
1YnIFxIe1ROpnq0tFKN8xphfpAzbYnegBnePOEvAdNb5rXyWnB4u3AjOf6rS53d7
xd8ZKmZR88OzdBue9/T0o4qqDy1oaWxO1639zu0TNiBkDUz4t+UECkd+SsUMkGkD
INoGEmDdFigLb9X3SwT9IizsfluOY/56yAlOKu/JgoEoeAOCWnYiL0Ewhekq48JB
c2gg4aEuMAQm9o9A/gO4Hwb32Wv2ivZTA3cHdBsp9OXNuwuxmBmsHqvvszYl7G41
5y46kU9hVutmMo4MzAHpHGCzyxHaVJ7yqfbIpRjfVZ8LQhFUDncmHk+Tw8U7jVq0
Sh09DdmNcfsIcuadPlVY2Xco14QrAvcpglVKv14al9Mpptrw3B/JxNMXEOszwNeJ
8in1yDnIxp+bJbiX7uCrfziMiBq/53HFw1+oZ+vm45jH5d/Wul1VakEZJP9p05d+
JzcyOQCkTevccZOWG16gnGdanQlMQ3HDe/VASyc3L0kpMfrUpWDIBlEoOb1h6GPP
ucdmyX1uocCBCezA4rCN40HSwi7xPFkiQklBMkiudR4niIs7PfN6RYlNiGk6m2WH
cEoOyhcU1+YPZQ0Ceszf7CHphlTgzXJ1CXl1flxqRnAWrp1EyL0kbgiEmO9eTiTt
aCGQ6beZmD4ZfVmNb3FBbJj+v3IYEMiU9PZHWsRF8V+ul2IIOxJ1IEk1Zdk6dEYx
NVYwmEw2D/Qv2Uu3wSNDbjLHrDD5pCbJ2VSiQNIuQdf7xKOH/FOYtEYuQBuGVeAK
17sxylX3pQX/Q6SY2gRqsowfcc7sYP11zVMoGoWykVD0d8Po2EZgMoNPe0EapvTd
XFrfOO5OOdU+2w00CbBu5G3qF6eAABR6ybFt/ShRJ/+DDeklE9IKAsHE7sVZxYu6
ZQLPEAfpkCayjj2qGxDjwzSmE2zlEEEoPTCiW6ntWiEvd+VKtyCiTvkeyruRJwhQ
67rEloUqf7tt4TUUpSXn6ju5TW7RMYpzTwSoH3GdvUDBqR8b2mw0BI0/uBOw69zr
qiM0a1OSJsNG4Nq1NfkJG/qSH23JJsSD2P8N32Y6cjOX58/1/qFXt5JwqvkHFhMf
o08FZNm14l7jaCB8wLKoYuW4irM6q8BkBF+OASmgR9xT+wBgX/ZCSnjuXcpZXy5k
QFWwQLqZcY6diiPGd8aX9Fsq8g3cFuMdhJ3oD6ujvQbXXN5I8NYi7cLeinyxOfeJ
sxFIjgESNhkO0GiB0NbEdeVcHM/04nFoMPMzi5Rb7c//o36WeRpue+HIv2ydXJ16
0GgP+b1MaLCHOQJYLi+bYvWC1sUAFz4r19p/evMVyKbqI1sbH4SzNbOLXzkn5UM/
RJwyn74z+oF2iWs1O+qhulRpiAYPR+FzLLI8Nj4c0BG0aJkGBkQxYEvQ4CXjuBDn
OeoUS/dP2JoX3+YNMnzq79et4i93J1Ki9pX6d7LiZ/1Y4YDQ1hsEnSVfoNxjQgE0
O2K1nayTn/+uQ1cOuHYQaKcLD/aQlNYl7sQEZPi5qrTlFADB+BHrD3qkRCGg9HYx
Ep5IVimWGR69BuHLm3UIcFnx5nKDVVr7y/U3PsfsyAo8/RRZO1yzQsFRaS4Q0XQx
svkqRfrI36eowN3fohKaRTbElkpP+g/3ryetDpJ4crAw1M96CKdkOaHWt4JpTvPH
QlKYqaY6/fiMW4QAJbN584QQCFfz/yCtlx/ZuoHbC5o5q75f/xrvcZc0q3uhHiUS
YOYPgLpw8pLxSvxqnh4VTxSBql2r0ucOxf5zzx9ujMJLEaLsGSCA6waKqTIRtLSb
AQF6uTkYIqAdqItdeYPhEg==
`protect end_protected