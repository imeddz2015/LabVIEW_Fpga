`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 12080 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/59UwEX+aE7FohaWu0/8IpTj7mav863zUNIsgIH2BWb
Uw34kZl5aMhQsSK68elNYCLoridczp13fXKCx3fEfyKUJue12Ij9mbYnYBuu8i+L
rAOzoClkKE0qBZ9pt2A2frgMu6SYsqcp9lxiUBu4u3B+FjBIIzMjYc8LrL+Z3xBI
57EGserhTTdOL4erDITwXpXp95hcqaHNW5S9aC1MZCsbGnDzuohTwRw7LoCUipcD
idZnyqHmjIEqGF3vEnZuBIQjAmCSGhHJn1qf3ymGr348DPGtkGuMIrP/Adf/9sPZ
ny1Pvdqs1FmTJPHURD525yejHV5U/akBihVAUaMIhaEZhXV4QANmspIiwQAkqh5Z
hL/Bxjx1fiGaB1tPMGYNvsv6dZaQy7wHkmS++XpGIT+bLWaho6QyuF6IcdSj0//h
QoH8kXPgxwzbpjaPsHctb8iBqfr0uq/QbVAkCenHSRIxOKF6foNMbVerM82Ew5W0
cf7EA7AMomnLHateqJJhHxrp1rvu9eNCOzfqMZqAr48/Rxt2alkq7ka4SUIAXOg8
hZjN/p5rTEFoD/Nw/SafxoWHyl9ljRqHKgyXXriJzXT2nTWFpzfsWWjHQgK7k718
BHUCRbF8sV8lsKs28WR58OCxbOPsRQz6CAZebjrdCohDH3MIoJJr9pbDAq0YvFYi
zEp1gd0VAzZPumx5cVjUlI+t6Jy5K9uSf37rWTaP6EfpvEPJg8ncyYBtfJwcGj5B
GEZVej3BDlQW5LvKlU37MFKA96qVT5xTtd51A2kVD21LmRbVTTca/Mi5BjGLM49/
ApK0ddNoIRXty9KaZjFk34Ne1aj11M1a2XH+HaBYrQhMXgIkymvJsBlHy4gxipjC
lpx2OhC/tDZix4M88vt7dd1vSPLuofmY4A0uELISBJ7OqsuQRGeirZKTL+gBWyha
c+EjpwOCVHepaOcJsI/IzMAlhBqxrQ6MEb+eCy2IUvowjnWVoaf67WjJF4NMzKV7
a0wS7pcgp2pqe9EnXwJ2s6NezQElAmAM4GeOxBhEcOaM+XAMTOeNVRJGzpMSRr1e
c8yn2XascLMw4c5RB9wAKG7hWOiMoJDW67zVGtnkkWcZCQe0rsfNwaSlgBqPDBeS
VPVIxJIsxm3gaJvTSyKZUmVaK5WrbU8Qu9Vrhv0xhxWwVs1iLpXYGeR6sIbBy7XU
kdrQDpA/gm6GTw9FdOFuAyHjciP/IX7LUmyWM7QVI2LQW9QP1JGv41tZvEMmAVy2
8+/lVjFTvpnbkf1hkcVaYzS6zLnx/c2QFTIsey7n00IGwfIgIdG6WTJ5NSEga3iY
Ek65CujudS4RV35IObgKVrhC0nYCxSQ7ZuyPyBf6HnLAYavbu7A3mb7Q7Px+1Hvg
y4Sepxq2dhdbcMJD6goQzOCDKxV1Gl5d+pVVl5XaFAS8DDuOG1Iz1vE3UkceiH7Y
o2cwwsrjq0z1KIBmlgu7EIqDv5GaasxBBORmpdlXu5fwdT3hCG2WMnbm0gHYYS36
8a1ITXiem8hR0u/lMR0iQECeu6hd0JPYYrR5GUdLREakYeVywygvpoaOJrb0cAiM
aBJP9e4XOA2Rg7R64j5+U7ONPYX2ydwfYXJ6mE9AhoU173yJXnSfODaW/GaqJjLJ
ax/bkH+zsbbV733VnSVyvml74h3fFBlKzHEt2ILJsLbitugFFFxnxlNBtDE/7mwj
Prv99axYts3xpe4F/cH3SrpfCnacb66P+fYz2t8QljEjngRgY4HtBzXlXt2HExBx
BfJ5oHyGyv4OxuHfYjHKGdYlInqwaxtoFYTxVIedAPzPVLHQuN05JlkAvuW2fVdL
qAwVUvz6I3mAoIIgadxtOTVm4PLT4wrQsVh6Nja6HkOd6ZgzEkIBT9fJUIn8Ckg6
DJP9I4t/EJ5yEgVPPQJAzrSHhAPFJj3N1LwhfXyYLIfCi4GJvFtOAW4YLX8v2cYz
/5/MuevHgJG3nMNsXhx7Em3ANBwe0sQUw5VDYOceccnJVg7vm5h0nzTybijXWvRq
rE2URznxyFabPj053wjXbOK/p77yVAX2pouW4WCtrnLtTrToJpAeQjLPUZM2/Ga9
iLeWR+eKUbzT5G4NihkovKH34hWdKgCfh9/KjBwGxo7HmBz3WK1xVJREBCw73o6X
WyDYK/MjonG4gneB/SEfVSRWFRGOdcXMvFnrkjIHW2Bh3djbJmOXhHC9McQ9OF04
Ab/CI3huYfeTxdxER7WG5OC2IEyh2Xmr+4Gaxt1ztR+XwGETpuFygimT6JFxEPmn
lp+YXzFYQl3gNOoV5kJtAkzYhAXSw82/ZF/2oP8WGKpn5sZy2LWbo3ZFpz17KPbH
cP/MbwTZU/3bZk3oJEG3Wq2TTzLksgCVjT/6bhEfTfm/0Vrh9v11vSjv5mMJxF2B
oPM55bEnrmRLRCL5d+Ss1ARi7uwSyzVdAzcFN6nfeoYPkZ2FIr7XHh11cAdiZbyN
zHWkEnFmhltLDD9Ph2rClNanl9Pha2m/wvBZyfcqqBAICtXiwstUyB9oEoxRS0Y2
wrdVL7i5VLpMqWKTgWvzFeqJC5QDFSXOiLA1DEy8blLxEp05LboUdsNAbCuWotdi
02/F7ivCr3MLi9FwFQUYY7DKPJB4XwuZqGgVX2CZ229XYCVhGNcRYh+euz6/M+Pc
orm0Yk6d9VUJ3QXrIBxWXCCSYmyQRd5Btc5dQ4ZHZK7n265AZpR8sLO+CQse43IJ
o/rxIjzRqOSizkcbwguxGUgODdv9cZU4D2H8Rbsitr8AohyatZlfCwnH1gYgq3pP
8C6Kw5idAQ4RHcXAXaPJOl74jbtwRtTS6Wfgv+BFpQTEooWHopkD8ZaqQzaklun7
sca+ANxIvS0z/i2N3xcUyaEwvVH3MdbqLpmt8JRayVYkQGj0aM72K323cEKFNNj1
AljSbKeOHNK5jimZDjSV2iLXHG+RqjAA3S4CaTOkI+zmHNPm5p6dKd0reyRXcYoI
L6KvAa25VfCFeqPAHmmNS5K62s+n65pi9n1cqTATT8LfSzi4TvJixBjXTh4KsKF6
YKIZ9yfOfeFKH42CtIgKtZKX6muisLKD2yI4HwaTuq+IHrAXb6AdLSKiePtyN2yl
YKeumlcCuuC4oEskCGWtvBZCgH9XVmiCpD7q0Xa3AAZjwznGLrFsdZrkRvDkgT1l
0oeqraWJqaKdkG9N0e1gQmCfljJMPT+v+ZGo7RI5Mqk/fXZ4JxhSZMBEq5RKXtCV
FqMDA77q77iQbL34DvwxPz1hKCwzPLxMX1Q6kELK6bIv0RjsnkGWUasGWSwquKIm
rqs/4owQkZ1U1/d2uqQbTWb4etvfHPgZyfYeGTgtCeocLzCo1PxluyIxtekIycFV
2oV9FUu3OUsG5ClftXST3gnbo7Tv+n1F3tII1WNkXknrHdsnxpZIxrwzGM2IaQIT
iw9DPDu8dN0j4qmC7tmHnb2RGDKIyjpb98WuGoTzkwHA+d8154860eRYqnWoK9uj
eEby+i1PXV9e80nvMMqmL4HU3ETGCoAyB8RrSKV1p6nklh3CGXNbGAEFmFppvEeg
yZUzsf9SPcd3jpT5cSoLaZ2ZqVt2Br4phdE2DgJ5eisdWtZgxRnyiVIJawVO/aQl
h9wGvIijdUt5R0eP79GYVnaIZ2fF7NOmuF4/AgoEm3XIoCw6/EnOehcJj6Hto1dP
MQyjhf5nltwAnBcVdzF2TpGlSPkOAb/rqkz2wY+H5TtnLqt8ftTs6MOqs0Mi0/mE
8miiRh+pKlp2hNQORNop0ZKKbs3pRvXPMsolJRavSaW0pcGVreSL19gswffFJfVX
THzS8XQFzrce9ZHbr8l4N2vTRjf4mKDq8fl239koSCCCsv7XZuIO4Dg7OMKr8Vqd
wAytwCw3mmwCAaHLEF3iuntSJEnrJMMHQZ4HHxT4eHKdhzTnTGE9jBGrmSG9HtAO
DvcmyvlJkQwZmmDKynSkLdEhJhe4Iv6+Y2gBzriZMyokzrcHQoC7uti563dWq3xo
jPYRWL7+1tLkjNIJH3ZKinHhIFzNTjXSbtx+X9k8hTInq6rRuaw59Khh/FH7ILnZ
xuZEXubnAuJ+Se8vlIdI9xHs8OqXcmDvWU1dQIH6I1C1YpMPsLQlT7FJGhWvzdEU
4a1ejdnInVfchqI8HJlLUDsmkgy8+UXexRWUAgWhG2C1pRPsrD8UwBGG/4va56HK
y0nFVMWBMgrClWL/I+TqAjeRLjmgCrH1wdTY+BD7v6tAImhZ+YGpvrA0VA728el2
AkJKX4iqgN6/wKQno0z9/MDKiHWYkf8qgrTztVd06qzluyzP57xpEHKZ6Fo4InqD
vsr+cc8cMrIVxtq4Ile7ypVbKeU56b4CPA3jCPPqKPBmV5M30xEM9T/U8JK1e3K5
WVC8PKmTnZrBQzHp4Ol5Tvw1GULNNhDHOC/l6xiuLdDuI/B5Smsj2pQtgLWaxAvc
guKyhZR8E/8FSJvYJ0HeMyVm3bV75JQ0DhcpVyMlcqWgYrr2MNMvwsZl0TSK3G+A
o43177ARNE7H6WlmxFudTSYBG1BeQ56lZrlhzf39Eb7E/kwrRE1rae62dpxXHSQI
i0sHZeuLh0Q8wBTWxGTdL4hn5St6HvWEyqHHsZo7sjIu3Fj0IPkfk0OAX7LTTWXY
v6md5qb7imJxdtKBzPKSA/Kl4etNpAJRsiGHZYC9LGNgCcMI0QrEokbLhn/OkPAJ
FbY//m5e9QTQ7UiCTBnJXJEwSjY6jC9JYOqHkHwCU25oJlxVQXwy80rmQc0PGCB9
BVhr9X3EAf89ujRLLRAWtk2WcbiSkdJVO4eEcmlKyZtmo5oDKcM92s0ALI8rKBA/
41O6HcYDVLNR7/7OT/U/VpN0VqZW5SfyqVT83OHnJnLvfkUBqk/FvfVNwcpy0pOc
bAOsHVkhJEzLaF11dyndOCYnxTB0F3EXzZFWsQAFAX0b2yhY563hhX3UfdTwXwQZ
NP2W9Fi3k123SPBy6CEo15G9V23HN+GhFoQroBjWtjTjdmjmohYYB4DY12OqGliO
6isoZb4D7hSpMzzr7rouPpXEhlIZm4D7wk7Z34fLsxx1l/BtPxtqUIURakMMniQr
p67PKPzfRcLJFf76jtR4ML2IP5tJv3A/oHmSljsSOQ72xoldbsu+Kgv5UR+JlWBX
vjoz5ehCJloD9R3/5trrDX7iz3EkxDikUWIBovXVAamrPzS0ITVZW8q4aKLeCK+u
i/4p/AOXnxUhlJVSnwd8XTedlcAoYCgA/GTseAjwAAfOfeyA7ZUR9uqsBRqfHlP0
1SHAiO2gUuLj52Dzb1wvZ2E08pqEIcMf5rOZyInHjuMOTeK8OwucSp1/GJAhBWLl
4dSVnTwW5dXg4+gS8AgRFCJZ3Gs7JyK0Aw/7bMNmRH3dF9H/KUh8pxXbib+jfPKZ
COk9ay6/mIYUAaxGjZKEn4V/HGy5HMDvwK05SCSTMPtlF/urgwDYwzdW7ECa8lEu
qPVZIUYbUcV3UJQxm5KmrwiF6cuTmzFPuZ3JZfqiG41do6V/CNupxKlVQa7d2OkY
U3xhYpL/8SToLJXA8LUpY688H3OvBoMdG9VdWxA4yo/82rrxKQFE+0UH9ePKqmRi
mbO8s/HJIGvVJ+hZz/Af/alJhHwqrNScOAYB9cM0E/Zk+XuWqsVXrTP+0cBvYXTD
3Wt+mAXglWM04BFBShY8IBqLJ0GFQC0Thgp/1HWJLVnFgDYDHi8MXFCRQvb173yA
82DkvVFwY1UHnDQIikRNhtT0jSg47mODPebNEFXzJriSfpfGpg0I9ac/xyV8cIrC
9YSp/S4XeJJE2LAgrXkrTxzjipb4mGHT268zz9dYQCpN65Us86HISuJcmU5feIXK
JJb9Txsn2NnnevDV8v1NDGzaB+7q1GGQ9kE+6QNPSeW6fN7glN9Ute1nvpb1udEn
Fv2yGjhpJnUU5HEV1eNWSwvzGvhQW9xTCWDfoibWd2tt7IXrqrZBxnoXdThk0d14
u1Xmap7SDKvqlTpLbsmaBG/DhdmkONmiB9uIRDSIWAIkCLj0/iVUX211Cf8seen/
gA3rntoZzhVhYuLUhtRxd6wkoiTokirFrwlHpvMAwhIvFnQgBgNO8C/ZYgE1+jdI
aKgjsI8hx+74wJaOOFnhMLxg3FLfk+9l7rYOYpt/d0HR/vwynly7rUiSWBKo4Bev
dHDLCYeq1bUcSZInkIwx3pwKYrsYvEqXb5nqi8Z8CQeoOiIYoCV7u3njxakht4sg
a5zV7C8Z9WvheX9DRCeedzZAHLYdDrak4sVahfRFylw3oTOt0vZ9BBMMXvLcZqN+
h6dLP/6PPNgHKFa2Qz7HaGZlYftzl42aFa/TM5g4wfX6ETcgXy1c3YsbE5CWPkqV
k/xPXLYRwf/vMt75NefxEgP5XJgm9yfWze95G9DWX0eUXD5Dp4kzovTontt00ekt
CX8dctcsO0q4oEuvEqJt7YUJAXSsfJhTQZV0OIW+S1i8eCECvN8zC1tSyr+QuUUf
hEmVNOfTuvQqOjTBpl/Y9A7boroDvHCURjRkVEvE5C0P76RZoHS/S/fwXNst46Mh
q3zOiDSzNN4PV2Y4va1R3ADKGwF7+nhGXENdbl0UDz3yq2cK4KsfmTx3lvv3EVGF
bibjDRM3zI/kxti9j7Ser9e2VmHtlkdaIoNLy6FSXQMDVhNjoReHx800AH6lwjgr
LF1zg2zlPbbGutnhFZTSZ/XuguGoXqpMDmGmKHswHxIdy4P5o2qNZi7DQH7nv5DI
fQRwn3nnLlWzCITXZ/ECMdfJi1Ea7YyV3Yi8ZMuTiMdwjGhffPu4/ZxflK6WPqhJ
XAnCrjBK765aKS6AkngAATxy93NSMgFQakYwtsmGTZF2/6nHl/17rMAQDKUnMPkU
ZlDt3Lk0E9fT/n5qStJwjNiXxFS6jxgpGSAs+MIRYFuhuNb+XRpBsGkAAjWl3REx
1+I3FGrmKbhybLuziaxIg6Nw8Kariq6I8GLIfagvgDqvRxDFgmSEHJXWV14mNhu3
Lgs7gdI7zr0PslPNTn+0596PDPV8KV1SSwXai8zwYh015O7PwTP0NsL0RwykVXYr
Gc2UQqJrJhzRmarc7WcuLofaCs+jFOl84VTunT948lKFXkenpGLMo5DbeM4D2QDc
wpR9kt0aAl25xSoS4acJOWOcHEbd/06FktlCCzaNvvbrKH6nECibK2lFWpeRIJ+Q
kyEJy6IJv8uYR8PNIaCfWsPXiZZGt28t3lIbc4tkWeWA2/LkDxux++XGmfn2XZRQ
Mqc2RU8KD155WwZG9/Z/A7Yp0gfMqu29V2LN9VHDSUSKGfOmuQy1QSKS/eehjtJf
YTQ9Mq1e1tiiiB6TBBb8wl0R/uO5J/9QcjTaLV6g3LKQg5tgLZ+i55sb/LAzT6hB
d8Lm1rJay0tJVypVc0ppFdYiz+nx2D8zg0Xps9geGA38KJcaY3cv/M7Kja2+v/zA
CjGCFY7iLlBDahVRpKoPUbW6s8izVjss9iJuNKR+kknX/XEbrTGaGjTXeMZnl3gR
/36r3d2Ov2j+iE7sq3BeADB03mp8ZR2RER2GyzQHYfJ4/LLJWE+0+cwybQE1CSrv
55ZATSOqnJly8qScjABHnOrANZ5TqKGKYz0Ny8KHtLqVUapGWqZ0olMoRt84Rg6i
r0aVSTcHzHRszZC4WFXmFfCOIIacQnDhhuT2FrnkhqiDrZM74ssL4FUfPoWh5B7y
XOStuZ3yuzG+EJHH2RoOiESmEbnpxw5O3RSjBT2DUgc96Bwslw4laIejM+JrG8HX
TD8vYBg4RfAMi3PhpIY8uCavlAOVDcPd1DmtyLvQKatWO0fFxkKyoFxeDhHafx/C
HnRaNq0dIQgBsru6qB4A8Wb9L1VMyxNkQAYzru0jDTGdhSGFuAFiN0+nHpVJMBOj
gxBkDXanzOMSvmIF6iwO2fmTOqHqawJ1Ty8AA5U+khi8W3JLJlsOs5bHo0lLn/1t
cRvJHv8dV3IVP9E1YH4mq5A4NFqUAh6NbX7d390GoIh6bSqRzlvElOp2JOZ9184n
GuTqaXFEl+KEX4ZyiOkd1mwea2esRuWXJfPoenIikHve6MOle+q8VGHdp/x+ouAW
u//QA/MVK8zLPwozch3zbo6u0+MF1teDTfAUaNguKS47/vebBWnbIIT4lgyFdkj0
m1dFIb46geZGmKdLhB0EggsiQIdRYKVZic60vuWt3w+pYPETmAZdmQDDQ5KgsfDi
ON/V1yt8yRa8Q66NTuDhlPPdKctdB+5uCecJTf4RvOPGv+eej03P/T1Wy4NcQddN
hHLre82BLRtHq1Inrb9J/A4OdCyGYV5RLgz+5XBzOtkx9HSI6mYmA0az1Ak2uHC1
o2lKB0I7Hux7wtQtlJOpryxfH9a2gdS6XaKlRM98SPUnDP1DPSHBhv7LazpVcLwd
l9MQ7EYBQRj1LWsFkamI3ZVQGUcyDb7ieR+1tafTZEzCiQIskk/9I1JO3MTd3zAl
2p2GFESE+b9v2scgNidsf9NWPJyTXs+EZKPCacebA5YN/v4wnwc+pSSfacUMfO9D
vEXQZM1cy2J2nom4f/ppKcNQ43+oCwR+2/JtkAxdXqt15ZSIguAnEP1WhLkLlIsk
Df9Gy6KVYeNapZUL5ttBMjOQCbAIgrKOIgZuCDRK0jTHAXzf22Ybz2g52L/vP20v
79R6nWJbXEQC9hJKeJcxoAWb/KvJFd/WanUxxdxmzWW8mkeN7FPiI+SMGMrGwCFE
M9ZLDKYZSHaSIf+T7kSq3Ra8II7J/CkJwzxmaplwgUeqsRGMldExFl6tJB/JqzCD
X8oclTgcWRN5e5qjWwcnCDzutmECPexPi2ShpDUyr4nbnHSKzhUR20wa59yarIAS
oFL8n7nkzu2K4PULomnuN1CQpGMHcO+Pmwdp//TAvLPveYOoU0u/h+lVzY3mgpOp
KmiaVTsPJYI4NbpO14MtPQ6HHSC05c0aSaYLjmT2m1iM9IJSMk38+6hqSXuY3s/V
OCdAgFbUGKIk3rpuc0izf22foCghMFMCVMm6Ms2gfqnE/JANQcsRkNXVMbYWSq/a
gcML9+XseJqgSiriIdv3t7msUEBIQqFFxEHjuuswpxmkVJ+1lIx5hHXCiCGbsfQk
kELcL2EtZfI+IsRg7zenWwhdff99Fr5uG9sBnyNPCuXqUuy9/E+Z2+d9ss7HzNVb
9J/AA4ytY7+UVTYfwYEsAUxXyulu+X1L0NekW6NuqkDxIre1Ae0EMbjRlbRB/nW4
8uEm0xRLyrPCqRyC6GBPJZqrc54dyWSs69NjDb6XBFuIbqaTQpp9P57sV3VhlYo4
owALR5nXPQF7FnV7Vm+Uybw7YmkcUoHTtEEhxcYo/HYu211HSaUqBFsRoEvhV6/5
K6aONuNfkWMifnkDxHxsfAM9peOsy3lLeOPo1UjZOEdNwmj5EcyUlsR/H5j9stbU
SqLtxdzRGPuKwJb4IS9G8gUnQGcvPp5wT0cP2lfQd59H1cXglHD/iMVRhEf5VNJ4
KMOjW4yFKUPnHxw3iOLsXKXWnaPrbvOlXlT/nfVp0jBL4oh3IN3itC94zao4RBGN
yQKD1P2bdYfnWbNRD0KmEi1UQTaf3E6a+feYibSFYDr6p0pXkIzZSRM9hp1E/REz
2RQpfBe/iuq2ZbIwGp2zUoz+0FLX0Dv6ZplhZ0YivSUmRIveooq3x6sSFham5eIq
FjlbS9mouInaC6wcBNoNYFX+945V2wLtK7mFUHxEJT8HHQpk15gL/loMeV524H2s
ooz5MsRRj5ugJ4TLIaDKEt59gby+13zuouKNK0qzkXyRccNBXo0r0s7AgQtHos+U
a/e61okryfyHZyjfemytHC19/7nzMCxQyE3D7b57XPQXaLmAGYLudXxArABwEvOH
BwAcPn0zTSep67TbWP9VNoHQLCVSphRg491GTUdo2X81GBa1IH12wVr0oaCh6ShU
euQik3sqBzmpVucrwugxHuJXVVvsYzQq1QIZ1xEI13iIm73paNkH3crcfN9VfQ7v
7ceM7T/w22bdG5/fqVP9XG23rpnbIVuqeDkAHegUu7AQUulJm5j/rqcSF65gG3K3
TJhjjlaRfHylXlXpe8drEBGG8q/Z3FyDsG/4hN8t5ZtjCRE/VuFEnImWC9Yx9RcG
HKZL9xXB3Lkm4xNQpURr/csNTfs9w5eYxjoSAWZyA8rj5mEmZQlYswxGZHe0AaX6
gCpbGjkFDWf8sJ0rpJjw5KwmcCrJidTEvgEziexGyri/IMNhDDNe33X35YZ7O18u
W/HmE7+Pc5Optp0DJvtPTQjqdHE6gbt/4XiixrAK4VBuVF12hkB2AzYsn1HYero2
9FiMzQ3HSU4I8RqoEsqDlUaSRh4sc2aATO4Yq7jpVZJWoOFUZJog12bHdp8XExSQ
+3PfEZPAJaIw8lfUASoUfeyI5ju0I18mu8XDtCkKh1JAft78XMlpxN2GdULsTrFY
md6L2zQV43sefiaQz2P10Zd5T6k9f8uSse37mOkXh/bKWg8ZUALUP+KuzYtRoahH
pby1CyZiRezfb/FGVnNEpc8fKt5kEvSB/OEZpKE1MilBoJJCtIASUXp2foeJAQV0
RYJt4zSBe2pBbiDaqyzpDho6NNvUZ1FYy1AiEXSn6TEEzYNAEhUDwAjqQYhcDs2p
e3jzfzuw+MltsxBkD6fX4ihlQbPO/M95RQAl0j/JwkOCNNt4MKQsC4Q6V9yaPYVI
YJtA5lyR57Nxh5/Bs/dgkDpgYC2NY+5PONyZ22NCSkezzX0hGW9YxwcF0/nz+54L
L3uMEAfBesVEW/33jR4HEeWao7v72DALaFO+WP7aCWozvapsk2DREuVCzizNobBA
1JSBcu0XQWwfc7L8lEOaFbarOOqAFdz7v0opGRwWQx/Jv5eUJPGEQRz5iUNuMB0h
R/9r8in3eI4l8RbeOigOPwBhxZ0wS8UKRJEwE9+i1V70OE3c5A04LjhWSQsrdDsI
zNDqZ9nTbhAp5p7auOSV6RKYR0z+XDL7pRTttUDmyVdKdeL6SXm9qVKyKW2UgUTm
7+OvwY1JqWrnLcXcA85hGWiKWIlTB65fs+83JnEmR1gGhInqvlH2Xrg03I1K2XZ6
5b6PC1gJIy8FAgHTmkdogaWm2Zqu4com1Cdom3F/4amkq84LFIAZYLHN2409SDwt
LfCh9wqPUedu4nSyqF3yzG2/SPIMF12hYez8ic7ZPV6ySIG3R8TfRNwPsPbhRFoO
dJTnaeD7O4TPs1KyNgfjLe1BNFtOszqGJq/bWivCextROpqNXii3RaqTBfClmQuf
kxOf2ZHYyZx8VnfQftDwDojU5BjRcMerwmXM1v9985babXxsMnPjykA3dTo/zqaE
v4rIeAtAdBt6pf/ZpjG5hqFG5c0PU0+MGOm1bVsIby2aypW9v2Xdcwq1yNqjuTH+
ilx3zMr7pa7VX4qyF/76M4ejNbuLWFAvs+h4M0XnHmC1wSPXcYFkMFjN+FLkcd4x
G5RxcP/UEsx9S5/LtXOexyscme7Ln2pog6NJ0cWrVk+Mp+NERbTL4JhBXvGBOJqQ
r1ODIzLrSIFH3BxGflj+soee2tonuRWRjMotnrLvmZE3v4O2Ydm7KLCTky0L3ZK7
cx7pgmfODUhCOJQ/a0DJzhdHwmHgFcL15olFFmQHTnHHHqt1qCpd6QxiOELRbpvP
7O+9FDJuCPDK7+FihoE2l3xeTSc5RR6Z66su6/6XFebX/iVaNgmw48zuMYVAdu17
m/e6xtcASnrhIUNZI6JVyPzGU01lgL0pasY6V7PZU2O4jW0QW1w31+09ei/8/j2k
ookIJArHZk7jlLN3NE2yiax8u+KsfpBDIb8et5Km44u9uk2az9S9ZNQDX+NcE7ge
IfLMqY9iSfNzW3d20ed4fdd2mvUacOhXzatGPlffert+VksjiuG8IAa4i9vtwE7u
A96MuZxMtyt7vwvyU04PLzHtxNq64P0OvbR0IJ4is+ztpB7S8GNQblJPRt5saICU
x8wTk4uD2AEdPmKSmRZiAWqZ1U03G7qJ0vvZ2feu9XaGS9lEIOgZZdeKPkhmVcYZ
cwz/D7s5Cnk0fctytvZPy8FTGpSRRZN8xi8SYbaFkoIiqRg8BHJa2yi3Kop4DIp4
qYYt5eosB5zdMhVgJglJw8D+ocS6LCUm2dmW0/aahmz9Ef4StOGOD6TKjNc7Ojk5
LZgKHT1xluGMLLl5BGoUrPpKH6GQasv4+37Msrcn5rlArnvjrPPYMxZPoAXPe+pN
1b94fOFod0NeDPhveHCb/5KsKPlEShxqVZbOFFN5lfR3i4VG3NgGX9aA7X1TLPaa
5tcARZ5/kntSAcyGFsT1YPDsAnCHu2MzLoxhFPZR/THrKCwwVe7aVKGbZSKOesud
NgIwXzoDfoB7+7R9souvBLe5kAPw+lUK0g4917Bu+b3JQmV+PUwITCIn9604iIuw
GO5IdRHqwFuTv/gHUAlFCyxIauI24QM+MrZLLBWQK6Z8sg0YEB6PTPzyY4V3TmWG
eVPlHRwYSMxHZC672KEUx4YObUS7dNWyMgN0U3+tbSa4AF7FA/JQYXdV0wq+wx0K
sgi7tR3IZrAlmTXS6M8COc+E4lpIFZn06sh70DzosJsUkpPqakI/ZVxjhp3VP4k0
7CMz1YjjQHFyzWiOA7eGLbby/DCayujHnsrbx1AwS/Ab6NFdIMARjOv5VMt9akhV
8o0lsx4O1vv4Cmqs+JO0nHywqE+2vYuIHYwvfEgVab2dhRGXErlP9pNqJcIAik0L
SyZpTaOnpUTmOmrNewO7uayoAI6gBWnfbFRHX9qTftvU4W8BPqqrhHREiMjZ28vs
o7CLhvBqvHRF6jjIpVvtkDPkxu4wd2gvZ6jTV9s71ls5z43cxUvlFGkyVH0TELsI
S6Xj1bF30h1qyaZBTAZ1QgS7lY3vbX9ria3Cr7u29IdCg5DjiCUFa9pXewrrdmw6
EOALrF70FETSYbMoJQ3aT8iQ+CgEngoJ6Ad1EB2ZmU4Q9ryMi075vf9fEtmhzLXW
YM7i+OMhtBCaw95DMAw4Pmg038ym2BR2Mb3pQjYuHmGNOo2fP+mhwHH4fsxxzen+
gKX1toS5T6Jt92hNKWgQZYZb5jqGMLkkDTzZciYScn2dAoLnZ766EheH8LejJWk/
189awq64q+ZGUqK+7kiMYdIpHBc8pFcQSh8mkGd02IC6TcOyXfX2GISUFIRT2Kas
9cEQRPw3+0XOWQw/xppcmWvvfrtufrcwOUlVjt+WdFjT5/2fOGrrrVnigzQkkNSr
xOBlJLAb/Wi5IELWdSzCJ+pDZlpkcVc4rsWyNZOf2vTl6Cu742tjRFTE377dYUAK
OgK6xbClrpK5Zd8xvVz5AAlIS+tI0wh4FSqZsFmjEkStoYAWEo9PRJU/HJPGmrJN
9vdyBgFX0q9h2l2dI+FpdujbhuOdu6QN+I2dmb6Cn5naZ6ArJiaSLHAQg+P33b9z
6h4IKDtHdbXw4yyxOf81P2qVRdRyq/htvYdn2Gp6TQHKyiXk7CNDfnzSq6ag19L9
PsOLj5ejXioHR1kgBTLnjxhNpqmu9MVpzrBkZ0TKvZKoWOTw+fAY4HC+Qiz+jEJq
jTN+V196GuC0yrSPiFev36kK/QWwXamDX7LP1B76sMcc/dmOGRGyCspPNQOrctIp
yZMD9nr0+bRLb3a2op6Lx5W+cteok4tXbey+92Im09pdnDubCU8HoRn9YJpI1gVd
nHgSUIFy50EydY/mpNFy7XuFUa2WjfM3HofTgbewxEPp9zdWB3+53YMhC/BXGU7/
dNocGqUCBvqoBe3E5zOqgRGonXSvruzTn9iWpGpDAhYWHMrNPvpIxmMrjR7jigf6
nTQdHMfHmYoGnl7XSuc40Bdw+KQtAbXwuO0CLzk4efAWxoXyzKcdV8DCyCZmSxei
pPdBv6gDajgNe2X2DSHCUTEdxvdOEygkOCl9Tjh5PBiqE1IiU7gAM8Ypm3cWKUrU
8R8CenoBFPOTEZwXNhnDPB59lBE5Z6UmvMhw8gbj1fpw1hsqZSV9+bwfFUtI340c
Mi3HQhwpNOO77R2RC8o7zChBC9UEjm3ODZ5M2aTG128Cjjdu8S1I/K7r+soYZKyQ
ETODd+1R6jbg1HGXC1bN9vLG+3PAMZkTaHGk5wIqY6dinytY+gwbcYYOfuXQPXLF
yPbBC0tlCSH95soz4+rdcKtHGcPkkDVqnbK6A47atg2YuVqSvSiNZJdQhznLFnNk
rJUYlY1eAe8ITxkXa020y1N0gstwfByjneNDpPOrYgPSoJrpYd5Tyd6n6Cdp1Uxv
Pz39mVFKowmFbV8y9TEGkksehUYlGHBR5G+PMgA1J73ksW1qdaesk6ToP+S7YN6u
twUeoYYoV2MiTJP+4YOUJGp7kGDaWferqZ8ofVgPPuKLJSVXwth9oujHYvC2dEnr
rU7nTCKDj7iOfxKrHvQDg7g0XRbcPOwxbekxQkB3g/PyeuTMLCA2XywPG7jsKb8v
USIIgdMuaotlgapECIxB2SzBdllI4t3+1Fcih3vmOXk65Rn82NO+DLAvDPjXWeh1
l5V5QcaszHg+WWdWY8NpVHAy6XqBONRCyFHCOAKPcHcDBSXVUKPKhsmmYQzyWvnK
lXv6ZNjJ8X7yEORUEiAWh+3eKB4cCUBr56TVOYJ348ktppNODHefwjdgqvUdAAcZ
w95ANii7vykKCOzw4DHowRWMWQzfGdqVHuCOai95Hn+lYte4omYnZWu/KU84oT+1
2kP8N8z4wE1+l0hZWjQGK7ahSbwwX2jggsUt7UGaqnoGwTYO4/IC5v9U/KXiuWHE
SHmBYRGPRM12TIYXRAcQIKXeN0/BuO2kMa3ktagV8TmiyOe9f4k4Je2cz3mdsOkh
/YNLNZlKXZ4uqGpE3s9HKO6QbF5gc0NxsX+b+8MjQ8ugPaslJYCE2ZD2cvqvZKfc
VGeN3IVTQzhJuKdMnLXFemO5+uNZ0BNgYFVBFBN6bPLVlniPzzQWfTKScpHqOGfO
49u7WWi+PCxUD000aF36HFWt4DvcZyYVEXoxqutlMdGnMsq2n+hZHs4rV3vn8eg2
Lgfdv+pIdufooMGsjs+kwfX2pMH0Ix3ef837sm7KJbvwTaG3aEj5ZdBNG5FUloiF
4os/7gPTc0ltVTe1TRpFC7vSq+KN53nBCu2N11Oot29looJ9UyWVFyz5B5pTuVEm
9myXvi68z4nCagC13gqH10WLeM/uLQ/9M9jYfveusba+mbTOhzVAhSLCdoW/oDsu
YM3C8Felth79IpUDF40ykZ7SxVC2/0qCtiYXO4prlmVRSDhZM3WyKbAlTa1yYczI
RZ3Ze2Ei61f5fQ1ePViPtvVMio9cWsK9PZa+X5TR+Y4Vt+0O8147iNnpuEIHzYJ8
NtmQCqAC4liBC8fi91VT6NipagxPl/RnyaaTXui6EHBdsJMxcCZv6ZzExF5oHXKQ
D1eWe/5Jc6h+BuOqUiEY7xrzJg483Xmd/J+x5hAdNKzgiyNKBM9kQUEb0zC1Bjuo
sn2Rq4U0atO/3shX3hjsXsIBhF4KGSpmYx6DnSpRnqQQkbvKRXwArkGRmJIzTZhq
rGF/ijfc+eaUME9+v1uM7ZS7eb5dd1gvwfwG/MraFKatwv4rlwytq9IyOliN91GR
E/sxfO3U19czDLSberdABPdAM/GhcDqxlFTvCawj6orxgS6RP8EXyAm1vgG/42Dp
QOGHtdOejTehYqeIKNYDsfH2CWXn/ZdGkpkXPGH4Mog4jtwP5ajhEOG0/5D7azsK
H8POawGkGaZI11iIndv9Rblv101y6QYXs5H2TnOESOlnfrbdRmz6vpxKFlLJwXtH
8fhyvTDNOJp50EPdNW0GZsnAFp4sJADW2cnLB6DtsQPyJiPg81sp3zUJR18uhxyR
1IX2isXpJYVHWvr11eOSpSuKqyY+eGha01Nc91+kIZjykKlKAeEWP9RS1fBBUpgr
K7ZoigPo4cXs9AUIrTlvEMvzDQQ9V9+4Hb1ed/fe5h3UyapNQIKYrtTrd3R4cIuF
jScDNqqztcJkKME9yE0463z8McykD0LvxV9zZ6t1zsU=
`protect end_protected