`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 9744 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/9huKRhRMtvnNqb3Z+UU7TahEoHV+T8U3P3ufru7l1O
3DlgtZzb9QxCbOjthp9+wDkjygH0eUfDrEl1ovhZG62Dy2soqUkD/L9mmtBzQlK4
YN27aXOSRU5yMjqRccoh5IfqA6IoIwSqMQ4kDH/4uzF7f6eygq3Z0g92+/YuoSak
YwYEIEWGUjX0/WgKfH03ZW0/W9jMxSyic4I5Wm+kNhFOI0DSMti8WpEQSdgJVuaM
k1CbMXK4sv1UV9FvyC48Q3xw1WhJWPgFvHrRpp9I0z05BGbtkzD0cT84h6nlyxDF
bIrqwtCr1qU9pQdOM+tzFRO2DtXO3rEMksJjIE9NMK/AB4e8nD+ZoXIEJmdynChA
0jRbSEVTu5fVK9R6RPUK5eLCUp184p0ol+ccTYOMXfbUVtV7kFY/QGCL1aK1+GRy
QJR97huww26WGpQxbKzX82afp42thrPi+/4zQNoVlauW4TIXCOaPZpTCsy5T1R3M
W9Zca1R1QGVBJwADsSpeFs9qNuY8bC/AjFHqNRsv4cJq37KX/L+sE/jfm/gXGisk
xspcfmhjbXRJ5H4O1JOUGhA5fWuMpN4d3VXVbkZrhTjJN2ePdxLCQf9U7cbl7VWu
/K1DeY6iR8EgH/tqMbKkSKm0gOtfaBdIL0MxXHi1njfCR61iRTJVspbJGgpOUY2/
nAmL4jGlIRaMJz47AR3iyOZanGJ9G/dfVjA5mgvNHswK7Vimsc6TZ0nRM6blWmG1
1KUTBEGDx6WVg8dXahFnPizrANVubOHwZmOMJN66EZZ41LeC1uZsIEqHOd1myY/v
H/HvgaTUF+6XS2xpYWPwuEQMc52/TW2twgH+yPVgoEQevljPDSaScprKHI+mRWDe
dJQVd/gSwzz6vEjvq3dFg4EGqQGacQzUbre4Sf6g4e9to9ndLjVv5+mvP49p1DUl
UXhkzptXk87oXvGMeaQF1azbvkfzWwYK/y+/pQj9RfvyMaX7VLwD95JrWfQgSC/z
y4sQ4yVTFjjaknCoEXbAsC5NSiWSSZfzADV0fyaysDuxr3AXNAbGayiQOHrXRinQ
EBpOoGhDYLeJHe6TvvvBRd+8EiX2gmtwjTxV9YhrWFI2T24jE1JsvrKzB8GjZ8CQ
Fa+1FSpt3nrMFEArqJsa33DJf9y5Yf7KFwPrfTkdEaEXy8Sz/Os2tTKar5MYMQEl
seLkOqXbCUAsUe1x3CeOn0J2078PtM+7R/MUctoNSCPJwTsCLakwbjRTo1YCgHmP
pH2U0AFtrC34y/aXnIDZzkNxFiAv+HW4eGMJ5N1gm2R6W7kSkMTcg5zRnPbQMOSQ
F73wGMpldhYHqKQQzZZ38pGKSg1gTwdyZOzLSOmuxUvrwbxs9gG95itYoJjVUYG7
Lb1XZgA9gpCFhYAKvV7L8yo8JQqybXMzk7iVVoQ5mj9j/v9jvbFqGqaTzXENP67D
3AiCgUkrN8wuZYgzpX3BIPHVBFtbAw0qUuDUcJ1TEx3RX5NvSZ2L/xZd3KIb2fu0
WdHZd0prfZuG/TrZYHZQuf3owZ5SsiehsSsSDX2T+7EyO2n+Lyt2RwAk8VT/Mov6
syxpLQs/NIDBs+f1QHP8x6duOlah/CV6g3gZqPMwNMrhKfS7FXxDsimhsy73mMqK
utgjo8675g7un15SdABo8W/yfrN1aDBW13FRpg+9FeqC41dyxnoY4xU2zhVGbRME
vnHEFsXQkWB8uyv1pcNN0J3G5cqjRBC41JR58VrW9wAtavUC0hZT0KFl7LqKq0S8
1ofthLHFYzaFr26V3ZcDLsyYBkRrw2pFjTZ7+3/7pGciVvtZp/EoqmX434KRkMZn
XvbgXMWpHWtWBTlRoxaDZpWYWAtV1GBwJYjPyGrihEVOz4Jinp2cc03iZgvRD4KE
0P2srb9hebV4/0jXKo/PmXgu0iE5qhVP0QUzQjYF8/0ZVpy78rqXhj2Q6eAgr9oX
/vBjafnfH18xKkBskkDoxsYKEtW5Es9HUNiOGpG3wkwLCXv+9GH0yrqHDK58iJww
mkte76O2fWKzTWJvFWot80WAKYx7sPOwu1EV5RVaY3ovEIROmQszmZzps5JXQU4w
G85H8D9TEtC6rMk8w6ajVF8XI+xD935qpel7G2UuK8vqV7VlUhtwdTTr7UdZWeyQ
vOVuel6DRXnHBQ124hJYc1qggTEtyYYJGKNtHPNqGP5htqWspQgSrN4FXMXCjIJK
p6CeovRX/d1nyambcLRIZBno2DNKk2yWRV0BtEv19m1gXDoWoCq0R2bGTW3823IB
NpHcpETPq15DSG5DFxSl4zesy5NpwtWtHZybW7oc5DKIQ3pYVkP0euVeCB10Qn1S
ggmbCgxwDi1QdSg1HsBeYTUJDDychaTVTQNFLfyXp2HnAGLlm7Tb7kGaZn16YlLM
xCH+NuABTZVrceJX/hXXcbhg6bY9S0qHIUnHpAF4lOtNhzLOTRyofgpo8Pdl/OYp
uTfAJ7gnPuJX90ZxdJif4kyiIlaqmLlkZZ7Bz5GHFYK1rpRr3MbYWoPVHdiBHsH6
ryx+pD6vLhbEl6pPmmmOaxWxIPD3AuMq91rdZh5L4diM9/P/LxDzuN4aOlo9ad3C
Yy+IPcQ0v9hsyvWeXIIushIeIfsn6y1SsrqS1/W9KqlsN77DnLCIyp2TDQ66eujS
hpjb1+OQmZ5sr/ZYslY+2ypdAii6K11o9VscirzffSHkqf8ksnugYKXz8v1Lr7ZE
91NlGTe++EAySuoAhlWnIEfeHgTAIAxirPHzN5Ngwg2tb5GSS0cuT+OcHLo3aF/T
DOEdQqsePrSgxC9QmyuhTFQHDu5W/538nVo2DXBDkbMVxHccefO9oi9ojPA78hzO
whOofBp1MDa/dfFiUxJYCc+SzdKH5pXb3R8VDP5LCOgUjCnd0s0lcJfyaH98If0P
dvXy+6yZXUEaijmj++i6OewjL8RIUHwc+9qG/Yeec4vc5UZuEPZ6VexuSe5DutbN
+payQLw2rcaNcTeHqSM6D7ovw0H3PDHjukeFdGvI5HOYGqeebniENoS0JN3+tZrs
NPKRra+2eC4PdHRcHU3tsYtEeOzssqK5XGWqJQKvxqQeoUp+XScxCFC7bN2cyv/t
zOkhP8NYvhccFbEqjIFrqPInrbV8r+E2yIPBrbAyYQg6oAqSE8aBJBe93QlrXFtT
0Iz+WyGw5ujDAw+qJzNDsVrnrRaWrYRS+TELUyEAx/YGqjP5UwH9QkXNVdqQv32Y
7hhPEkqgiKwSmwZy7ODgZqhQ3gK31TQjER8w7zrwEn4oN0032yaSPFkgGoY0mvNP
dQcxO9bnLoQ3/VUEnoJaR8oS2hdiLKx3BIcHVR9fii0+EXr/3yRp/lwWj6A4IbJM
CPyoQQPxT/SOJ6AoC21Kkfr53qlwFuiKcrCGHQF26AgLTK1Nj7ohJUGO/9quAan8
3EUd23q8NxWMCnPCwXA7W9tAaovmnpI4ckEAL2CDIEj9m4k7GJjBOrhykep+fYWR
gntMNIimV96qZUI6xvo63cI9ui1JLOIsNOlWp8zXLSnKRMTDsqKtbYaCJVhi3N6k
dcVLhr0UJhk07kEx0zpPqQcVE/gvgSPns84s/Vq7QsQW9uVsBTlhG/LCgZMtevnj
Aomh0yts4RDSaMjSBH6qjT7JBnkc8g22gBfleo3hKnRZ5HgtKJiDqqc4JVYGAiBD
YHqgNSIYJkVqKUhUlnuU7cgpYv9zuz339lbHSM9riaED8He7M9tG1B3XRzfUnKDX
NQcic1U3NQTMOT/1Qx1m0QOOnOJ4KeCNF9gR/9d23K+8zgBfIwGSCZWpEmg3WcaX
NI7NJfyx8yRapBF5IwAVUxRx3ABRQTLABvDgQOIbzMIccX7+dJYOhlw5ohsOc97t
r78ZG0Hxpp3LDadfW2rle11rX6IguU4i0GG8sYMbkru5n6AiiHuKefQtN8IaqFN1
uSnBclnsd0F2IoF3MORMb50bwUf952x7arVIFRRUa3Q1yBn2q/cjtOfBs3Zw+ZNI
yMxbgl4CwmVOS51M0IojVbjRtPm7oNxAv6+VBapoRI9/S/JDAOzv/jpWIvuKTm8o
m/iVpCPMf1vw+Lq/KtN4FrKw09n0qStcY3JZPIof5fy/AzU7f7DWFcUbDWqYOS/3
s9y8cwB0TDpH8pWK29fgZLk0FSSnj3wQ9Z/zzCUrm1VBnrJEWGMqtQQFYSEwdpo7
FB7JLwZP2GVLi+4FI3qFkFwz8NNnAci9pIYOPEa9jHWi1MMorUwbzjw8U27YikCq
ZlSuW+6QiYIoiPco9J4NupV1xRm3qu06CoV5I4F1oQl3ILmnsRM/aYbQ3ShktOmZ
ksOLgbVlFvw0aW7lLa9ApHtwx4rGv+w62PCJK9zWaQsw44948v6f+0PqmS82lfV2
0kEqDFQpVqGVxJeWjp1w8AmZcvcAfd/Iy+gVVmgc458SiK9KooVAUHZIsMC43POL
2ayMSRMcx8Wm+z/gxztrRng2yW1txM0/CD+RGWw3sRmpmheeaN6PHIoMdXRMJZE5
VirZN+HUSMflvAehmr1+iN3txj/g6r8Nzx0u/SDBYTnOBewKumXNDbjgHIeY1YNS
KMaVEe6cKKeel9N/cYDiAFrAKtYS+w/hCp81GP2BWdy9TTUmUJhE4tHKWdeL/cKJ
LTKZiahxWuwo4TwvVf8LwI7B9mQ6Tc1/EfZnxzkqj8aNdnUVJYpng0I1HSzx/4s2
0WXNI3WlRbqRtBM7mf5pMvFcLEyU0HZE8RwXEiUlTn1RSOr+1zHXw0w6e2aiU2UB
wEx04Wmi+SW21ayqRV2z3psHEUKQo/red6oEU5cdNloRbmPoaIgJC5+uBh7jbdlu
Pb+5zGWTkSiYOEh4UwwFoODOibaLoa2CKhjlFeZZU+l7eHi63pqyG3PeAwM5EZVW
iMVxuSrnGawCv32g32wasMg3jLWyWh6sUzV9+ngghw1TLiZLbi+gly4y68cVoe0v
6/0Dnak0Fxpklre1kQQbuZjMoX5KXjlwTqZOe3AAvkNN6KClsUYIizsWGMHqA63j
tfAiExr5rmOOEwjv7PV7S8oXGDp71w4O04ri3APcnI1HWZWs083ylhzNJE0SXZnT
4xn3f/E8vADXYEMfolGJJGr4BKCjKthPAZk2NNzc2JkuwqZAEJNnVgEDwzGBTuKs
CsSehhBumfAckV5Tzfl0ZTbzhaVhxcnjbBFCeeuLlJJd86E1xprAHZcnhvwCTG//
oRX6O0YWLyXnL1ylGkHv5cRYkdv0sj7XCXzYjfE5J1rtJQNlBy0Cvok1PwdpxsGg
d3sdi9Jn0233WXV7ECpWcLsSnFbIoD7LvzAn79KZWfImhxhlE7f63MxxWfd4MArW
I6Wq1V4jOr7qSdoiXMpsFuuLcbGBGP5RZ0CM2QSFu5Ifwy/sl7uU2319+LyKlsLk
+S2NtydGv7ohuujujnN8xz8hkCQnl5EoKInDup/NeXvdvud91OPGuBuayGLN7KBO
iKPtG1vF8HPhIvlJ53FoBeO+O/Jm8fnU0uxhnMoqD+hTGBk1gtZG8wLd9MCfoFmi
vqQKGOjXwV7iolfcJqz9Akadt2wqjEjOmHX1rxIgIOwHj4JIKl2hn+8Q5LpJ63X7
eUsOnZC+ckXFmJJ20LH4reXcSkPPSYp1fAwo9QL6WqjempEBt2/KDx1bwY5363IY
2d+wpJc6kGMVzff6OxyIIT3vN0uabNtaUtJKXoR7CvL5YsmTTz/F6o5zW15grvwR
PF/x6ZuqoLuwZj5jfaXjQo5RMabMQivtuUlJpIvRT01RaSJHczgF5A0Biz+3qXaT
ANt5eBLb6Con4VaOa5Jp1tlMQsPFwee1KCEdigxf3Sin6HGoy137jktzmy5krXOa
zsXsyFGJi/BidjXS2r/I6GpdY5YiF2LrQbnUlzaJqgG1zSuasBuzoBrKjGaq+Ae2
U/hUuF4AE2TUCgboS21ab+dqLsdYyG2oqF+zxhkDl8gplsgu4FqIri5CTpPtrFj3
ADgLLwJDubbE/N6r/0QSM8FgzjoKKmZoHjPP2JatuK9+60QpbAyUFSdWmtvtjpa2
9Ja0ZVVxfXwPINFzIZJeU26lkkKiRjQNFDt28wTG8pMfkKukom8WS/BtqM/yHVwk
UG+eA+hQiA9REteyrqFB0Ua3oNr2cRbZOwh/iiltthce6TT8mOOrUrwctMphtFtl
PcRXaGfOabUQOrvbL2vijvjzIoR2lQ6fCk3X+Owd+4at4l74VCxiWT1OMu76X1Re
AOvKN3P0eKJ0cSumg9TYkPakblJamsO7TsbkbuwfRz4LOnczds5eM06cK7JioHR4
bR+wIHY0mE3BzfE3fcI6rFrtQ+wf6xw+Q+FvAKPakjX7jSOcw24zarSYC0PU0/YJ
H7LGwPaWuY+XNN7uLJb4DdZ+JuVVuOW0kwmNESdhmBNm4sXctUFmBXCuXcjrfamk
DO67qnPNlJibmUiB3lYF7APNY3jlPU8mB9UlffxxUmpy+d7oF1vmeL/M1vMDhQiq
30B7Rw4yMJ2+WfKr13tlFByrfjkCDqABuHMtxSSg+zmuCC0liXJmODr432arVSe4
cWizH8TWuHmme5FH80LIQbly2tpJGvJK6V76rigOxiR2v90HPb7TMXyLvYzoMDxR
cJRdnDQH0J/Ql/V11fQ491qtgpKjur1NVfA0D4bm9+mvTTbF3dyYp9zzB7joSCzq
kLllScngP+AXSRl9TRLdos6yCATHybEFcSWRBxuWJX4nBHCOgBM6eZIPJ3CUXNA8
1kZ/epLowREDK5HxbmRpcqQzSaYPfUyF2SbdLQWC5fLzLzhiWbqw4uj+NaGfXeev
n6wWx41NGM0/tvl1YDLa28nvZVaihs/Wtkd+eAUAeo6Xl0QlFTdGn4Hgpwna4rjE
fRsicfBHIK6/EN/9v+rkiECn7iyARxetS2qPHsqc93DA6mkTh61ZIcLqG1Ux7Osp
ZY8JPAa0ukFxXg2O1gF9bnkrgwoH8U/urlqUImNWcK5WR14zaJ9Xzqdrcb5+URwB
r2xdVe4eCt3ZUOOtYBcQsBLFuS/5iiWqgSfOp7FS5pUO0XUpz/5lNM2Eo+GhCSlf
ZcaBtwZHH3PZWFZJITSeBJUnlHONQ3l/Nt+Ime1bO/mYMelFY6TUi3RqdSgxRWVy
ExQefGq/HVyyhw0sSIxREu6GKjMlNTvsTn4wGHVgzMXNMlSMb8KZQkGxNFgw4c3B
oji+FwDQp8CvkMQ+++uMrUjBjW9Vjn2j9VoDHfsHXRKR/0BJeD/pIFHf5CHb24Py
/PKTO12CWkZhkNhzp4YgtqgD/+XCkJH4nQizwS5V6CVZVHg1PSIN9XaOSNKkwd+Y
4J6NZDf9LZQd0MRYh2MCB7EEfTj2x6SGjF8VmWOaMblaG1VeYkFrpz4A9cp8VP4j
kksNcMIXO2ALADZoijWRbtLIuyBHBJ8qdLg4gkCQ2mBpDj5+XdpHVRw0/r1C1jjV
9729nUHBGsptZz3NpgYnKmB+wKTr2mxELhLeWHSrN8VLA8l6HY16TezHc3KrVVvR
itUcpKm3hfNzxTtjSfBDC/QYPqNnjKFOq/jasBuJFSJCldOSBfR/bq3CymVyqU7i
4e+PbmEwsyslFbnzYsOmrobCRTH3KTHEO2fO68svpBNtqfK21YBW86d/MvmDzKc1
U5M3z/n0mVAQqjmtcMyfdo235rsIudQPyQ1FNLSca1I9OQ6O8OFDADhXh9cDC4XR
yCn5dbFBdTYFcYP49g2wS+00hM1smwxxZM3HrVA4k3MGvforxwOEL2n5DGX6IcPn
VuJOW0jSZ9P/RTdVqdsZPKAz77NcutvaWAziIkZqygQfJe+9im4QXOZ7wF37eop7
Dy416DGfYZcfVD6pUuj07Edx51XCUHLa1DviFFpWWGr+c3kUZILIlzMN2S9zYSrj
7m23bU56wJpmuLVVzlfa1zBecEmMO5tT/pOZs3FiP+7FOBa4ui4vPhePIi8Gbp8p
Ote9sy6ItspUB4dyFa7AzAjhCzmGx3ZBtrbQ8CHHfpwkWLp1BfYvw3VS7uzVbpT3
/wARPzwp6OZgw3ULFslsXVZmaSKlqOGqzKCG4+jGtkHWJDHtg3G4iS+tfC9FN4WX
KikOKQ0sDEKoy4lfgq6ZKsWcSmmEKNVBJzgF2vubp/kp2IX2zezGfPpWKfN87eKd
jNnHngSZyP0jM1vMmRop1qjQS3gYPmemBmC7vBuAvZIe405uqvknnNQSOAjzbnrQ
OK5RRk9oa5EScq/ic/J8cpfFlFQT/LEbFX0FG5nixH1LneWO8DVOFpxc9NWm2Wdk
/LY7+kpMfGHG8xjWVXob5HXWZqIJmKPKA4ERTCzMpf9je9OlrgN0zxPOIWdweqWe
7t48VNL41tRsQfDUAmjvQT1De4ro8znDnxCGtCJP9HceicSWWEFbXY15NcdnvfHZ
HjhnYasrFG9kVjeN+vcGvE5ZUlhq3oSmGcTh3B1TbQk7NvRn8g3852DWU0FgFKlP
5VLxQkZ1rVqsEX5BsmiUFrAKGtZ6lrXL+Tm7+w5SD77PnlOtbQDjW3dqntF+9sfI
OORLBZC++jwKIvKb2EoH21ppS8cgols77D8O7Gd+mSguwRW/9VgmDgDSPRVEVXP3
iOrJyCknW9fqbP41kDE+4GEgCFFQMPSiiOCrF/nAGFvtWMWvwsUPHlHptMCKq89i
HBi/mt5EhMAnJnbJgWxsKCiKN3OOhZa0r+X7c06Fy7PnL6M3luHvqB6d+7I7bRyP
h1DZvS4oG58w6+ZAq13BqTB6mDq7vjw5FUwl4KUABiqI8lEDZge+pWZfCPH6deQ1
NGhyef4i09IKLQM00fHRj3SffTIp6mbiYZ+c3p6mwbeJP5guy0gjoSDP8EB/Z1Yv
fvhAXdDCQnwNDpvUcGsU9tvzWgQn/5VLH0KxW9g338c8m/bt28O2pFfRVZC2sDvv
3diZUz+HCPkXqrT6qY/Azo0HrQeThFp1qhEkqbQaJ29cOmkPttCf04FIwL0dyg/C
68mJF426LVUcui290juIR9GYsqa/FFCLGn7AiOGVAnggVTuL9NtmsP9JWUWyVcSn
ZGSysKndqB/pMCLCgvdJb0GtJPox5d022wkCo/WEDDOZLATX2olroF2CGo3qGwjm
JVRT6lnMQ6kFNYyoIpFegdRXuxSr3PmZhpzG3YLj+VnvrIZH9KfE1fd6vEX5OTNK
z+d3lUuGb1HIrOGQLei9KXgytZDiNiiJtA/ptyAxfDARM6EnOLYVIoyw9DeShe0a
3h5wg+svJsOeQoo5vw2Frl3r59gBjtYLEbtG4kU+d/S4wf39HnQtLGbuZZ3NYM0D
aWhnp/gZAbvQQKwc1davDFyMTl1yo7/lVG4RUPgITiLMElH6YimkW9E4KMW004kx
QQh2RfbPJwoJf2hZJw13r/TJ1hYkBZeBE8d2S/9f4rHE6BJ5cnj57ZvwZ5kJMKjw
N4ictt7dTMdC5nqjrf9lEh/BH4IoxJFv/1NGRi6P5hrnKz555K75CTS7qDU856QG
LydBqQDIhSOaMPZPNdIUgmUub2+GZRIbf6j1ctGXibfdJZFXiyVPqpGS8zWcO+Ue
5w+r8S2Z4A+GhtYj7mATwdnK5bIYYeOvnZntrZzu+Dn1FYyO+uBadZ/ge2x8LbGm
rC6aPvCFCEzC47aLzOc3qn/k11QWrOTIxuUO2O1Ibb+S3Mj8G9Ur0gZJ6EKhBOUH
pdfD+iq0/P2mvtYFbGiZKnEI68Xq2ZW6EKIDQMkKFEpf9x2wMnPD94G7qkSjRpOB
4ATl9gbElKYtcX3+Ol/G7D3te0rElb0eQL/i9XQyxqWicbnLwtDkGBDllc60Vo05
n7mCBwt6jwzP30NpL2f8D39EbwvcWDYPmYOPHkm04Vv0CieLaqfYns2GgIAxlrxC
2+8t3QF9ULmg1AS94VB60xA5VbElaPvopDMFJPuVSTSk415hSLDZK0dfceFh9L/r
gSxhAOjyWlQsZ809XV2nsFN52i7QLAlnJ6hQG/sQjblGC9Rl9UFCR3O5NJMWd7Vl
+S7vfMWQI/VNm1nS2afBrIIXLiWnsYUoSLdwUoscLL4yxIp817bh3bMsn9wvpNAS
KbB9nT1iTXQaxFktuRJwJaKM4BfibBzo0Vy6h9i8ko/EMfedntHS5LOy/kUwaHiS
KyNdHwTPg+Tl6M4JAct3gL0y8+ZmlQqRQJyaTSQyubyBnsXHIC9heZawye0rNBff
EzJAGvpo96qILPY+bQGD4LmRN7UM5p9HguADtBPcDwMrVe2C2hEXhwcG0WDWwxg1
4oZ8jotpr3HdyxrF4RhPA8C2gaSy9HlIUNkKhBdkIogK7C5QpP3Fccu7VAjPNz4H
714gJQ2FLhcCcrHMZnYzyrppqhbJzap1MljUl+kQjnFouz4wqY6nF8OUvdfwDr0i
isq0JCSX6msXEFaJO6tSodM7YLKTsglFL1WGFBTaFrzBo6bcnmQZF5ioGPsU4uZw
bt3y1PrYBLodVXApLGHWUitfck7xGFwgGqyRM9hPhzBVGztppH4gESFcXL1eQz3Y
VWHkXDKmsE+SS/2LGxixA6GgXaNHQVpBNzUknBLhp9tsFEOWS8KPHY672FpxBidJ
zTUuiBV8K2PtBfO0DdNsCihHi+V6FdEhPG9dAuSEVVuiC7hacn3/VTtW4lPgYRTk
Tyt2XN9+O3hX9NneCDiEa/AWz9HP2d6rl1hSFdKGsDgnKeVR42EHxWEt7P/FgSwc
A/RZaS1VRM+6T1hcL1xgSWC0JY0iw12LivXIujIkaqW7Qvwx2QM7+sR/fSYlKHOM
qXzrXcEY17PmM+94yKtRVwlJNpf3X1kgqC6626SYAId1LCeQ059AKtduF54bp4q5
+lvBpsF/yc0VjgkVwGgldrKi06PoMVhUZQt9BWg3uobkaWtMb49pgPSwS7gl/5x7
IUFv9SgGimDIt+nvyZDuFUD9LbrMCo8m4wtZS+ObreONl6eAMO6zVxxFIpVSDpHV
UseLvPLMOkO2vQyTlyYBrl01ALfBlZHjglozHlVOIr9XG7KYBqQMyvjvnx/K8V6u
NcARlElR14VatvyeX4fkN+MJPukP+GI5GMkeNLcjJBAHEC8kMthsSOR1lwNiz5Fg
ONUQrpGnMpZNAyBe8QEzEt6MX1ekmYAaAwTaWl89nVyA4QJx9lhk+g1OnghBMxPZ
4YJTsvrPN0nsJGX5pmGBvIXe806c9MPV9InSuODtIQqX3tGiT13ZRarvYDyYoMtY
7tWp5++dt2CqePint3St46VqM/XUd14rF/F5MktNy+emUZzyUx68QpQ3I2YjU0Vw
yjnDIEgylKxmskg587kwmi1KOp6gs2xXSFlEmY4NQOOJUzTEKiFv6Rfp4jLjZpZg
QCnicIdGlOitERz22wKxdgoFg4GgW/9WCj31ZXMUcJTyo8Ny+2C8zPR6UMwzVg6F
Xo7U7AqB51qpNH5Tp1Mss1h0zqe0ZMkkfsgBY3etekOW84TQsqxWbq1VwAMmElhT
BYLlNutn7gsSjkPwwpmk2v/6il+cfr0N0m/iODGNVF2SvlVYlLBXj2N/PQX2puUB
lcEu8JXIk9KShy0AkiS570uS3KcH2J4K0T7AnKblM5wnKt8wgwMLSa91CIC/EAw8
41OnRbuYxuEijPSWu+KHR0UTXUrIcmvqz/wpqtsm1beH2+of3K/0EZAKCDPuHiB/
sZQCwhlB5E7mjypsdqxhT9XDL98SQyCgcKL0uswZ/aeCI2xfhaLZLWo/6ujBT4RC
KD/7+rYJ+cI8zIKVoO75flf7jBE7UNlzPu3JisaGtRtRc3KsU9C90sG8RaIC3vem
OWq2gYnSE/tXNCn+LXvh5LFZREs9c6/YeD04DQVHTgnqvkx6B7yYK7pCkVisHj3A
CLZ65FxTr86Pqh/QWzuJNffgMoKabd908/FQXmWO1ADmoN/3EWE+CDknj7/1f4vk
53LwIuWImwnXdi/OJvkGi91KIR97INHwHxR13G0uINM8inz2eEarHMU4R6rADdtj
GCGekiXfuhopBkimdDLt5BoWE0S6cBCcpO7wDNvSRr5yaIIhXvvCe4DbprYONcJQ
A9EEcVOX1qYWo6JT/gGCxNT6+md/wP/XZankEps/7V8p0iGR+FVzusYHkWSQcZfV
JaIBVYOlBqqt3hxTSoIm/o/VXSqfvMiaaLHr09mFcVcBEADvdnDWCJT16ozQa4JA
EJ9Sh3NWDmVwLZYMMItJ6runkZoKlmgLJXpRyh7HiM8adZ8+Saux/3MmQhtaxFpw
zx202jOjlKgGxwtz2cuWEJDb7/6Y6FKip/UHqC5/p3NA6qU/xaF5Q6urIRbBFV/z
5VBWJ556i/ziMaSH/tIWIflUcyz0BZBSXreZobqgaK1geTVKvGQAhIoL+rKhgvlu
kZM/V61te+DxA2KEO8t00ktiaA8UnGoTOG1vi7y1etaYCL9zSQefsVhWIdNOwZjz
crlPPKqsRdUqaCGR0q7keFXmJfnMPXIdSKr58UlqxR1k6VEQgOMIcGHHIJ/+teBF
ypx7KrIwEWr+B1rxMsjZxt3VP8NAcxSU8HPZPup5DgRBK3o9gIS2A/3HH5nkW8YW
veco1dGoHTYMJmh8JePgwom396RmBXphst4Kq5pt0EFDUbFYNnQo1XcP1SW3dwOC
m2Ure57nN6a2p18RGiQxDGYv4cGHgEiW3uwAHZolCSYP7xcBIfof6y+ZpOih4egX
+mA8vGxZAANP/Cs/HnacwQm3J1Z9Cvj7ndGi62/bJDlhjEF34MiVxpgpWOwmHet7
gTBzKHrLeTHH2a/AdbruoCLUglRKXmUUHZVcuJXk8hxGANw6PdNLh6qFL0O/TXEx
sb6iAa+st8VNdAwILIYmlPWcum5MUDou36FM/mj0DxfYbdOVihN3u5W2q+jtkOv2
wLoHvFsLEXeH/TKlG6FUGs0J9SrJlCb6wH79qsifxXGDPDU3ATcL+xujeD8y1ZsX
`protect end_protected