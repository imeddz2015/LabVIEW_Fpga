`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 3280 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/9huKRhRMtvnNqb3Z+UU7TahEoHV+T8U3P3ufru7l1O
3DlgtZzb9QxCbOjthp9+wDkjygH0eUfDrEl1ovhZG61irtzHhDPS+qHO7xcio/qA
+E1WCVAu1M7dlBh0YKMlrzZcgbuo6l8ywvDiTYPlrVn9g090ZJ2o/tc+4raM/4Ma
awWeMnL5iHmDpL++WLEZ0q4gKRRYItlMgLBvxZ5LzeA5ZyDFcHWCgPKPe/kFF1vy
ZT3gWBShk0FT4H/VXxMQ/gxoMhfX+jK8iGpW8mjm2+bSsIPO+riknRqWmOpjjlLa
l8gbEk3tnIKvnuYDKhyTiMCyQ9FJfZPvaE/DGxs+42ATcorxT9S8lUwNHFoqGYh/
KbuwRDZ9wyJEBl/3G8I3wyG8eHNRfzWuFVJPPgRF/ZV9M/RUONOo5dyp9HBdkJV2
kxQR4LEOZQAGXJfdM8zA3xayTUFLN70eIPQJUAcD1qRU7WhiM08UAAgn6yZW46M/
7T58PHM74jslCeWNRfm7BA4BtGzZ2l3WVNXKh/OTYcZJGha7eLf2vzE6pfRO+isD
7cvFvaibJI1VBCBPQodzwAOU2Du4bVzAU20ls1oFg9EG0rzx038ihOaFtKHU2QS8
fGC5PhrETSvOvDVW9vc4WwxfcGXEbXDa6D4uohyZtPmXu2d1h8iPJJN5L3F3h/W3
p1506qL7Uy43o0LnBIiGRBPk0GzzNicAv7swhGVHqPechjEesjLqi7HEoBrL4v21
37UlW6V84JD7XSTKH9HmKGb2dRtwuYP9WTHiSUxpuzJucPHJ72lPqLP4uIBq9j6B
hwRSTTnXxl5JwdyY8XALhjl050xkfZbEbmgb+3R5ERBk1BrwnYp798dThdk8q0cU
xlm8HNqlABxwCS00CXap7GjO5oUhRf7rLUAX6EVG0jaCmw/IjgMkyfxRaHpJbvId
+opgAcgGfDFKrNBqOMHk8ISvpAkeikv9OJmJ2yeWzrDIcPbi8DytJiDip0w2Xz1G
jiHbBXkDAqsvVCneevYf9+DzZn1V85Jk9jEilaTld/03MWkx4xggBfU1RNi3mKXV
0HpZ7s/dsI07I8vG9YczsmuaLf/5Fo2IL0e6BHF3cnYA127QiGgDfCXFTRg7rzQk
8B9ad6NcjLhDqClqtHMd01+TUQLPbPtLhV1glPSFhMe1b4SeRgCBBxuuEEnO1/At
Vn/1fDUmi6CM2XyAfqyJvooc61iatTWQSR55RXHBo/7adMpwyNbRDrjivY+6SQQj
qN2uLGqVx7k5HYBadZT/O+Y7SBiz5MihEjXlrLlTUMS2KrJDltDvQyggiIKH/Gum
lz+lW74NmqRBP/ROZ+TMfFhX2dbFzNWMAxT4CvbTE4bikcu0cG3NQf3IT8o45BlM
0ixHhWdWYBKl+QMgZl6H5KSJZREzHM6G1boojaobIjW5FQhRJEfA+6TdaXw8Vist
mb0pNmNEgcdPkm7zn2Q1z6CUYGTNNgdxeK9NCIzYjSrl6iLwazo7goNocTVSg9Y2
tP1CrUwdyQmKGI9li21W58ylRIwzjYCHnLsCW/iRtHcPd+ikCeJq9NKaopssscAU
SZ4LgfwAxcf2OorrB07QO7+m22q46+uSKM3wejnxyK3IpcB/opQd55m2qox0YX4o
G18Cwqc2PYecIdfxu30qV48ivf4tDMD0fuAKVcA1RAJwi983R6WCcXYYXNX/UXxZ
kOvxLkmNQTGlMsG2aGdy2t1ZoeEl+sDZnoh7NSA5Nlq1kAd69Fvxx37z4fqc3rOg
yZG4sVSaUV5hT1oMkZRhmmnsh+ncsyBkz1LWv8Uh3fm7AIFaVJ78EJ3v0Dlm5F/+
f/Ayl9pwD+XKazgqCYGZfou7Fw/oVHw4l/g3uEEOf8rkjP0SBQ2qH9EBKtGV+J8o
3oA1Krlh1GNkba1nNYgu8o/ELkBk0hs/fPeXjoPmG2u5ZYvSr2kYfyf47uN0gST3
R5HjHGN+UU1PS9q8Gg7f5pbjOjhJN3eNRiJNF5ervo1Rk4jSS+dGiRNZiKwxZF1t
SEFzYEhTnFrD5/23uRXk8TVBc841nD+5GzU3mCZihJI/ot68R8VHCBUP/JvxZ/BC
QobbWEXKXGTxj9FHrHBSKwCD5F4mIF1L6/H4M6baor9/78/JHE7BOfww0Fwi6hyi
6WMZFN755kDb/xfds9YWJ3e0f8texInN8Y9FI7l4z4FNklOfJs8pzM8OGtQdjLqy
nB+UoNG5Yt2vJ9dm6/OU7miBnRvzz+RtCp0REOHQbyUfTjvL+gJr19VcqlfR3hFP
X7X9EzOKOSdkh6FTND3EY7mpWO4BlT/gumBHH8GlbKq8pOnNnJJygQRKC+0ETuwZ
dkhqbYbkPwqc/NHdzr1xdckJ6rPzXTYHML8vjOK0Im1TTsgB/da7bG97BPlsZwIm
6uG0j86tt/3J0b5r/RrgeBIrFrt2TLdZIon9skDT11EincPON77zNJVgyMAQ1qP6
VuJQTuE3FoWp0CzaPhb0cW3aa8rZ3BL3HqtMyV/6eeLEtSrzgJ8fANHsnIejyxwF
1GFtI4VDSigbljCu3eVfDVkuTJ4NBNunQCfBB4WHFPVyR4Gw5JiVdGGWz8XXp4le
7HiSeMIUP6zUDVBfYemS4dLepaoNz4rhrLMIt5ZL5WtBAQs3zwd5QDp4nstx3/SR
Y+36HTaAo3tj0wK2zQfhutgBRhEUwa+KzvKdRB98Jie9wxb9Vmuf5c1jQHDS3cYO
Xe65SI59W/1pQIMcGuq43V3k/n9yP3i8UFWrBcryTwzX9C/+BeBIuKdDq5xZ7Lsz
PdiGZimZ2tYBph+VFbblqRHUNv7354ua9YX28CP2sqcZmzR9RbZ30jFDujOJgwrF
NFYr9vHfd7WfODx2adWmIIxR46spGlaFdJ7WsjsgJC0v8Q+lVYye5KKYUFGHkJ4B
Ty9xEe92FaLYj0ylBA/KI4aBtw8LS4mHosWF3qp/rj008O+lOXR2HBvzSnIbo0ei
XCDrKDVQ+VhaV/iMirZPSFclS5Kb4wJiolfv8Ut415qUSR4JfXmXojITi6vcruWB
lGKXYMgZPneLgypu0abdm5Sji6HWXqbDearFqxliFV/TMqRXW5EVPd47LCDHqpu6
TlasAwOT3ms9pgtrkhsMGS3Rlugy5xGSasZNsHdjjYoaQol9guv1TiEki4G3ud2i
DQdqZmwcLfq00p3R0a+Cb1OOr7Dhj6VPEGIp7Mc2sYZBF9N1xg8KmvRGMJwN9VLM
8ZNocWyo6lRYMFheoGw/ol4cw7ZNK1iGbgWr3AFtNbKL0suliA9Q3LSjimMdfUGc
JLQXDVRMH9m0vpOQ9Qo9hwNkhRObTPg9Kt4KFLIPlZMo4Rtbjpemb4YnMPRNArf7
orNxDqaLJfplxOMwFOiKiSsoRBphi/XVU/+jfR9h00t58yojOEE0SK8A3Bjc0SQg
ojh3vtslIuC04cZvXm4yulmqCW15gPRpT9KXXHiE5rxtqbC59GcB2zlOwWci4np8
rpbbBKbhFtgJHuuo0vBWJpe+Q0xODH/6JZSoXVT1idgi34ZxghVpxJMZ1kJg8rEn
c3OmSVR+vwN0SFiDZV1hH/kr67Tk7fQ/daUObRCYz7aj7XRogQnz5RajDUehQCdo
0uARI5esiAxdVCgCDem0rArlpQm2u0XQ5ioSXC+HD434pCbwLjlIQx+QPwOBKXJM
PhJrXY8t1etJ7T+3idkf23pyV8FQMp8URdP8eOab8dkETrZJEGjKObeN+kd5h5D/
NZgPghH9Vib8iNjAivDefrisbaeBcHxiqleqSbUgd8H3iimsRYYMtaglt1y6YT7f
mzjhVRHKGxV05XDansrMV3aTK9Fgfv0VMXj+jL+NhWHfyosD9lgC1UyuXzjKFNTB
y/VQEs4rpLMNZFTOYC9oHhgX94BulSABfZFatEE95VNsYoM7Bi0+qF+TQpx2MxSA
FwnQF/tZwngxfyXNT+WWCwrltzYYPxJXucmQdCTOI+pGwcjwj8KpgLv9qu+s1cEZ
DnmYvfvNwdZEnTYuf1QoutOlByKfLNtgxgGsAn3dak/FKsRdWl15eErVNexDx+gQ
fWYDLGCrI0LEGg1AEUoUlGcxteiuycCltA1uL+K/2MmhtrwMrMUrViCWtGVWAfUQ
2PIEcxV7aI9PeVvvQK3V7j5Nf5i8nt4I86//ZsMfO3LsRAf6iRsn97h6Qso6NaXV
dTOOoNvLn8wS4fMFTn6cd7QeuijoUDN7iInWf4Y50J8Zwswh1x9h7NCNnds0VThF
E0jJDF5iP2/ej72lXof/AJo3NkSNySKI4+GJTkmWIQxEYXpIqyD7MmcqZlhaw2AY
L29lFm1VQZfQEglQ281K3Q==
`protect end_protected