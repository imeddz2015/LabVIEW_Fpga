`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 9776 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/9huKRhRMtvnNqb3Z+UU7TahEoHV+T8U3P3ufru7l1O
3DlgtZzb9QxCbOjthp9+wDkjygH0eUfDrEl1ovhZG62wcdxw5bCL9pgdQHinz36a
kQL53w502ndqhsWLs/AECIXN8qIxTg/WW75gypP9EmzURm3JBgOU64sRd6Vzz3QQ
ELpwwxSwNX/vfCeq2R0IS9CbzctaJ/hAPmO1x4QCDtAm4sB0IM/neWMLj/ssv2mt
CU1CC197eLW++UjB4ZIIlmNSydxRYZPZl+nr+Nn+oD9AuevoFQIkHHyZ6yokXbb0
L/uT19hRfuHSV/LJFiyC/Zxmy/b7s9LNsTz/BKspBOUqHmPAwa4eARr2MAM2POK2
kLaJPXQ3UDmL10QQtz1WjJc9vfeNYiBp+LrJXaqJ4vrONDrsNzdYM5ORZyPTAclf
/yo7sjB4g11DiPO1fPvPZP/sXiEh6094nJKlEmqZaTh+MRq2J968P0beMOI06JLu
aoIWOJHSKjzzMILwz0H3hgawcmc0EdMYgBXS4qCMxscL8O0rICBO4J7xpp3lGyXz
MMDUhZ8c0CMea4cjWqyqd31QHoPspIxCJxLKZor+dPlI0qx0C7UG6tOPwsv/apo0
01MkCEMJIDm5Y+U+T6qvFgCQROZ5tOdjpaeb4I0Bg4UuQg5TgdwcMd6Osmh9kM66
ioH60vtD9sdgcPohqTUIzOEhxXgKvqhVa0WjF0oBjjVctZnpH+0nPP6prDYmrL8D
L6Ou+YDwqFJXSm+0+tFLnqYeZipHOHgK3nXxu23nXKmUsqC3mJ05hkVJF8ZKWcyF
tuf3NoiFm/nUAWQNAkr1kliPBF2xYuI79hj6I7wmJI8Rtd2khuAnirU+tlvNMHXM
bE1h1PorH3dujHfh0nckcBr4Y820oFjNb1HbDrr18fBznxlBOlCmG10szgaNbgzy
YxLkFwoiML3Az49aCA3eZSuHbk8RgYH+JfVrtdUfV7r4pm4e86hbSHP+YUPN9SWf
byiUBykjDuEQFHoO7mA64ZDrAbalfF/j/uG1BohmkQ9dIErLb+mwR9NU8Y0kTxfb
UjqdFavAlUEWAincNpVCQleZsjA5PUfqL6t0bvtivs7LDEAaSVKeFM1ZaB6X7gwj
nx2+SzlR5dXxvzg67PPFWatiBZRSV2fJYqk2mpo01jeQUrCKIQMeWBBb3+Sb9oWL
0T380Gja/5FvS0tHBF7AnDrAC4yi52biV5Qn+rwOuoUKKmM+gqfvbftS9Dgv3xCB
4OACEc4prDlpvQ/rNyitkNIW4bn9vYv/J9w/ehVUJHfrEZtF3piWj3FmLUWOUCJa
xpRzj0CvEbsh6rHmlmnp/ZSmHa3q51dFWSt0TjGefbIG5GqEK9AaDyJYKDcE26HT
O/SNFwId7HZ9mIf8c4w05WfSVcaUYXLpDKRS/B3TPjUQc9ACiiok+eGKaUPyqDny
gH3QtY9iQ1/UyZY9HC+VdXhN9kxYpuVXi8g6bkMH9LKvatf4D6ONx7Xk2pb+2AnR
0WDxCHOYLnbOe5ROG0/AiFstgSHmBaOfd0E+G1sNcwW+CcbPuSRd05m3s7eibIRd
LuQum+eZ2Uq6n7XH7z0Zh74VoYO+hTyEJCnp3LXlptThlGRblKTXoigURCfywo9n
CCbSRtbra1BChhpxM/me9DjskbwIXVz5aIx0t58/QlELcwZSvFxN9cIF8F2q2Psk
9Bh+xEX3BLKJ12PLmZvSnmPdA3dnbejwYgxWg5nGAqNlBdTY7MoxnjNjX9kbUt5Q
Qx8ATZSI4sKEn1Q0/VOJyKSEp2pgl9oqw80kQ4bwygipVkyYxKKdumlp1Qw79VTy
pdgmG9za8JrhViUKqzTaBX6CuAcSadeYcZa45B4kd7r2Sf/oF/7zS4KfJdTdYaAb
TUJKZPm2JRE0UA7A8FU/xylLQatkPg2ZhNGtjgE0e4XkyqyMxKfLjRsVA+Ejxu9L
je+pNitEuGrffFGdwsjSymc0kobGaHUEBwqhD2o89atgd5K0xhJheaEv/NOglGFg
sNIS5ps8FN7WovrqittA8lR1nqsk+LRrxA5qcfRv1694zzWwEx4uVaF3k9DRz68c
oyfxmgpvmtrNTFvb860MWB/G/D/OMQJ7VZWRlMoizEHE+qCaH2Tnl/P9oIAYNgUk
g8urqWBYE/pglrPA7hQ8KkyCoTcVLzfEr33vGXe73N3hVraSCAFsG4TOKhLJXXq/
psnPudT7kgvSekTdXaGjXJawN+vizR0pbA+puqwHL7YU8VtZ/oHcbARQJtsxwHma
pLFSS7ImGS+rdiEkcPHSRIMwu7oD/j4LY2pp8Scypg8MC6B2vQ0diMzczddGMqt9
YM3uM7m+tPSytN75PgOzzsMRwRUnuoPZdo9Wk75cxBwASB3+wW1u7YyoGAeJk1I2
RywTHkHxa5o/SWZ8CJpsWR0OsKHsktKh2MT3gMIqLD+TW86+4kEKKrAnBlXOs9P1
hR+F0SHStP7o/ZY1iL3DgfgRNxdNC9gJIhr7V/6McPwPI/CJIyeEUaTt8w5JvtNi
anK5bAAO0ynVMKwVX/LyRXqGxdItuwJsm3NO0J/DdzrvkB+SKXiKetgr7yWeUMoZ
94ejrjr/aqhjBdHfVi4YMwiiOkgwUd7R4EpmKR3866PacB/78Ncb2j/nDcffwpaV
2BP5ba3KctbML/jI9dxBID7Px5N12fPtPkEn4h7daLwfWwoj0nf7Q4X1N+pYPpme
fmkwTPW33Hi5yG/WdzZYrVcwF63x+A6UDllfuKMvQstKqVpyoFV+J0zx7D2OE7nl
eh0slz77CQZdbcUYYbAdtfd88HGfyzkPh6Ef4CNtntQQ3NBOgUiAsnHt8dO/vP+7
4RYKFNALzkBK3eps/gqWOOIu5upLfOQ39A9oNg3bQUK4EFF0B/xVzrKegtxhCUWY
Xg0Td7hDzSkMmpNHoHw2vk0X6QFMe3a/LA8JTKTuRs8C84CPIWt95ZIEiu+HagU0
kmHUQc2ZbAgJzLZfXZDFKgLpqj8LJnnui6hfUvZpNV6SM9NYa128ObIh2DM83QOh
zedd6jU5p11KIPyfbezmuA7m6omclvabK9ATLp/yWN8QvNRmWBndNa9FpetkZowI
1sftd0IZ4GlkGd0+kemRLUbu7bx5U9NEvZx3Y3NErnco6Vb0U65ih2lyNohZ7cWJ
n/++4um516v3J0s+8IFMLbKXu2vBSZaBNF1aWRakb9CPSLLLPz7VO0QJLXUF9cPk
kspY5RjO6lc4ljD/u334GwTm1OSjppwjlRy76a9D1zC2akzM9/YkdACInZV8ReHG
GhiCjjNDVLpb4MBh4sF3CGUranDhjgHN0W36v/QCufCVUfP8RRTDtQfur11uTu2d
yPMpainbjs1y9mhB21eX1EUtGZ9mCvTj6Nfjud57gyX8x1/IYCvS5chcyue+dOHK
HY4H1b6hWI7ApMaeFrUJHy0DzKYZoS6uqqivMAmn5lUm1us2oHbxRHpU64q2e909
9y4WDGoAViuiLqeFCISBvfk4jdLHgG6B+37/3C3kedmxbw7aymy9uNnoxonsZIeX
l9fYt3//LoiZbVqjXM3Cj1TjFjBXThECxdtfNkdg171m+344UD0A/TikKpvwAqn7
fHLu1efgK5L7y+lcJNoqzYhCppWQXCBquDbrnI1lBJChXxa493h4qTdv99IP4IQh
75vB18XIfe/CzDU/J48l3d3H8gKx6Qn3CX6OHB2QC63EdDMroOuYPaaRQvjGzP0n
DI5OT+FIQSaJKJX3yctaw+C3kOCOrCXmL/OfKGtjMQT7qt/OswhirU9FnaZR96C5
xGS/cdy0AUHxcqPvJUPT4mSJijdJXd6SLPLJvynSbPTYWX5XJ1/8+pOeg9SoVt6k
6b948sLhQ0u95bLhFJl6Icau94SvvJCRwMHv/R3a93R06s/1ekYmpYtnQh0RObbR
gUEaGasQVVHqLTpb2q84qOlyUi4jynurCITxL8+N1mIAzlH6MCaK/cnTL9yZsQNW
UaxWDwk+6sYEMlv4h/DekiiB0cQ9gU/R0eEZQ1cb38vWYUtYM30Re+8U+XSzE/BQ
aFvCoHcvt/+9mTowWCf9u7B1RFoCHt3VZDMlY8Oxnf+HcMjNakLm9Ic2Q6Cm3oK2
lw1V3gmHCQ7+f+1bQQmTf/wQqv91snHk7B4IkfOM7GjQru6WViyCqHG21Pjw82Ru
099YCBPSTUo315EnMB+0sZB7hM60/9brX3GBDfh/4TqI2BG6WiqYezhHW0KK9zmj
iAUcQKApg6E7KuNCVCSQX3RqMfMwLEen/bTcesqJUs64DUPKalu3u7ApvGJc6EDV
08wG8BkpJFhxBcI2wAvv8DSEtGmw23zQfKHYmIZia+0AqAddsemCVdXZPpPg5ruF
fJrBdvPhYdGp5OUZJAQxeFKYAerQ0C6rRYA6Lv94hpo2TpGEYwi4GNI9SFVTnhq0
DdttaoUA/q1Txdo/LLcetO+yE8DbTwl15PUDGStVDd+f1B0hpg9fVPlVwIktuhjh
pfcpXAg9D1rrAKbQUpDWlq4Ks6ej4lonO2uKK+3lcDTiw8HJ0CEMmlIcCmAnBwXs
If04EjtF0Pe+yfvywRJ1OUC8Y6Ftg9QD1C1VTgm5t6KBufOzwk18zXvgzrBJqsQI
6iHVYS/g9Q2NESeyXazpgOHbaT+5U7xvI/w/Dmmjw4t4mNB6yku/TZICv/XX/T2Y
YZHY3sXLibt8MuHmj3xkiPhaMSiq5FtZY/G2IVRyFN47LHQIX9Eha4ABxqLsbWLp
N/prCAENJoiJPbCXKYbAKsjjCAz1fBdN/TCS1c3I61nuViuYgEWei+1IpztHqfQU
/5JBn6Am8D3FQ8YXzYky6fozAKBsl1WceWx3QBAIZB/f4wDraBWGCDeIXwxyHIj4
wyYAXQeYWD3P2rWVgdwejdN0MyOQ/OGNI6OV+fBio12JtN4g61k1TISKg6F4GdqB
vJ2aE4m+qRVy5LxzyYOW5IaTZ6UNfip2xnVPboDnToyjWQpx7ATryvBIk2fZUtSL
LfYol4Esy6WY39s39UifetP19ah7i84GIwWinm9SFfiSNIybsiZ/9pGs0nFmtZFf
32mZOF0g9B25pJ59/1PSOexSGMcBUxXdP9EoGsnTOAp8UCWjmOs6+UsxYq+W0Fyf
RmyNqPN5Q6qdXNhHAe/whSC8Yi9i8wp6fF1+X/foUdr0wsfjheVb77X16RlZLK6I
jdWQq1hOuBIpPseUWZfbE+oEOBDabE/xNKjfHpor73PC7tbBtbD8Z/n0PNBZfj6B
geeemS26xcR+NmHRTOMJWpvD6KOIgF9HdIAGoOPZ+dSbTSaGlJM3p0Lqk9R1sSte
tAaAr5a1jpGIXkalQThGEhiLUPopmwnQJ8Mu9IWc0Fi0XJenh5Ql6SUsta6UKRie
9lqH48ygie7k7uh4npLwsCR7nXpoD924ce3AU73gZbhLsir+MUFD0JlVuTmyTkmd
PTCcLCnsQk2VCcf/7oAuICbjAlU93mH7i+d6UM2ZVLM65Gl9fIR14ltIy12G3+dB
A9p2G+FarAh+Wj+7qRcOIAO8SssAUdrQ9bdW/H2G5t4K+0ecTL9n3y6DuhgHN5qq
DmaneHokJZU0u3V9hvsFuofJ65rrP7SDObe3NARJ58jfJmfVh1KnlHsQYHyBynxq
iFcjX3igy6IjY+aaGIylHiy6H28ainlLo1DHxO/9iJHWp/OXB+WxKd2HDGB+0POa
KvQy0OnbdHf1d/Cw2jW92CQAQFnIID6sS/YMO+GhV5+HGwDQzkeI/s9Uw0LvkBO3
soeWfyfOq9S6xAdmldlK5zdsYtFLK5lSI7ap9UKnmRbzkJewE2SWOJaT+L1rswAA
8tknSImLzsmGaDRNMCy3WpprSW7jhUlbyrAmbBXUDBw32PnWwxbnOUsfuyEUFYIy
p6yJyXw2n5Fn2DRQr54s2T36HoVXUgkd7XLMKEECXGsQN72dmnP1sWP/4erj/LRe
4lz14L6FfO5aq6ZZts3wnJ3o0PjkPYnEWhWQEi1LwZNimQtZIadz4i9Y/EoqoDUy
oNgrOlGMIFlSVgJNndjg6knmF9TfY1uxMRjkM16fv/yNXscR/+00vpIrOeXAG7Jq
WuWagHPEHWZH+gpvUGy71FAWdu+8NNhQx7Uw/K6D8v1zBFqJYmRpu7xqisnC2qwR
9SWZfsGDGn7Si4gSyKyrtnDp36wFT1BbrE0c3nCz9Wx0RGj8SonQiUAY3Nul7E+5
KVrunFnRUIdvAdCUxCeTaj3/7Epsd/vl2+G68WIOC6j4SYQUtOWz9RRkFp4k5kM9
N0XKWCA5anSpgpropNDHMyFqd30IXKfvm2RM/OkAcemxhmFPkSCY6b5gi8CaVzVN
5P/rZHdgxULhZHjcx1JC9Gqg7FBQ8B6lSdh+SSk9/q9PLXzg7ORVkDmJA8YBuYCq
rmXiaFmsOySOH08+PTBEKt+pRNaEywzwo/rU1WUqDmU6IoFv36nGMDUXzYL1045v
WPw1KIZVP5DWMTLWl6yx7KzFgv6MDfnSW9u1Z8KReoftFKT12ShF1p83ZXR5x1rd
zlHRNGy7ytMiAS+mOltQoYA08VdygW+56fcZPpS0w0mPyY15fPsOZqhlW2i05+XK
HQghtAFIDPUeq6vonzKtrFJ4HsCzipSUVgTQHXTQtW57YOdkoZLIkh5mk2xhQk0P
htAb+LF6tHXPTU48yPaCFODPeRPT/s7/pJfjfuvLmNJqs74U1FCKlgy+UhHK83iC
to6A1QUeXd+sw8cSeyb5MoV3S6UhrLk62oOJwTFDA63lovk0RVW+RoiG4uGxP6Kv
F58RY0ljw4niqx3WC0bIGuOIXw5JBdSSxUDZL4qd/16esbbzDzWkV+YETR/z26tz
egqpsDaNmKjbnnuDZKG6ch1Ul2RqDkeWbTzmJJmnBd1V0bzl7WAGFco2JOV0djzG
QjCVRcrODpfZ2nUSXAsMfB0mGjttJ5AcFp3jlxiTYYqiZaNOdLlaTlia021yzv2A
SjGQEv7HyNyb2/MGgXsp61jhjZ2ZAsTQg9q1fC5nISoZKLOCPxKbGmD+YwZE307z
Xs2k5d+WzpjcK0fiac77mrRyWTiS6qF9kWL3blSN+LkPLzI5lHUoN3GbfliJEzEG
wdYj2XkrMnX5dK/dop/Bbb8bCbmH+0WH6lG+uUV410tqf9ZkvzZLJSgeVldAgHxY
m4fSL9299M8TgG9H43/zo+MnQ0qWu6xGYjnzdf6738XAktpFP+t9h0eECMpz+e4v
LFrqZpP7K09thtJe+B05Z/HsbdilD9dm4+F5ep/Dm6oVEm6aIDd9BEzTBuP7iiAP
rCNJ+LzrFcJViINzU+iToR+2efPDC9YSXiR7SAjqeXXkNj4OpKjPYmIL4kRcmRjS
1TG7VxyKyb4ar8OlzT7/gkW4wvGsXC1Eq4YQXr/D8RU9YBiVlnejNjtLfhNZwCyo
U96toq52jGc7mvpq/pTpUU345nKrfiphhGeCUl3yJdtmN2l2YlDE3Piulak7L7Hw
ShITEylyQeVHn5nT/NzeWxP7r6Dv2nh9xSLXJ2PGaSAXyt81SOyWxSv++fXJpZCa
SRKBX0uO3IQeo7b9CeD0imizOQf21gPBCe5FLdvlsjBmvEi7mae7CW0dHmdQIQfn
T19T8MCHoIzsGTaynfTIrQsnYTS250wGrqn/vfXnaYrt9Kvuy6WVTiP/ciMJpd1K
/jAGCKuLnKy9QS5eSeBd1kBBajMgPj1kSOwqsStHn3MJikqzBEJOA9L0D1LrHJ8n
wUZXe96Jo15TfRzDRUt8JuZ746B8Jc9iJ7EUXtZoCKXDjaErRe5WHmL0L9vYRiJ+
yQvgPv0DgO9AHoaCQGoDjGS6QgtUC8BOF9a//z6I/Xa567QWF8sPrpcqgogikgFC
vRiPZWxrFZsEDVSGai4JIIms9K25Deppr5oaql2E3Sb2fKI4CvA+uiprXehQCJ8j
0S/y/Bd91tLnRQTbD5TiHPuAzn8heTglmqAL2qctWPJ4oEe5v5ZahjlRjBrbV4rt
uVXbFsYE1B40OyboKSO/SlI9Dq2xwkfdwcfa9IbLyXqJgRaR1Sa0GFmwEGMvza00
v50ZBJrgSm2PiTrOg3jGwSXo6joSTZT+BQQQHiDDXjdoPDtt1mMrxc7vossB2DXA
/8fEfHWKPO5jBgLTzWhQvmvvAsGJyOCMzHjICXx27gQ1ridGh/CavpIGAZ0Z/r1I
1VdRfggq41+LZkbxdWcRN3Y5clgQL9PBY41PtoQqF/rykGNPLCuRt2BSKrk0+I++
SLUwDpWr7tKCKl48N8BiN3ZLA5OngUrPiahmAOqcAISueXcdAhQuuNJ5ysIHNwu6
UkCoagt30bBKQ6OZpFRb2+rwXllOklSURs1UbGPuRsaHNmuTupGc5+/ZMSbAEf8k
0YRhmL95E5kX49ns53NzXihXgq/M30ZG9Qemz65SkwjiG1mCCsrNjRAbS4pd3xx9
jrUtZsRtknMU8JMvQmf+hvlANUA67/D8ldAcMHCYYUaP8g2rVLcQdERhhfLQN3A1
ScFZTcHgGVDK1kdZD2xT9PqmLWWJ07kqbxdze4hV73hwJeWG03jNGeYeMfXILNeW
J1ZLD+TmlYT3E+L6ThkZbH/oVHJ0jpPnsXz+jJ6508RIWZ3W8tpqobU8ZHEHoRwX
PyJMILzwuJk15Nk4XI+IPPlw4vrMRsgHuaIBpi3tt6bZMGMWbjrd5qAU8UQ826By
cASMyGKs6Yvhj7zVvV4RKWHjRM23KDogX0f+kVCx/pEKzIQancmgqphjGxGos5H0
oWUbTaKLlzYL9DHCuczmIPTEurRIzjjQnOswEOGwwYocJ9be+YSYQfbV1Am0Fv0c
e99/RkrtELVGt25BfwfV7Nf7DPI06sSw2dhsSOB1u1L8ZUFdOiBqANeOOFFvX6Cm
Ts1ia2ua5uzRptYc3Nv8/cGToqaRHlJTPLydMMl7v7sHdKb13o3hvHAr1qYt5PZE
JwGBL2/zG+ggQi/ExtueleDzm77FqnbbkFiuC7jD85pMUTgfvwwgmNNk12lRp04z
vjanRhYs3L069x+F3ghDB4fJQwlR2pEVZCJ11URmCsotnzoKz2mNIUFfg+KcHCjh
0c3WjcoI/f2YVMGyXLa2lgzaOtHuIWtLeyG0fOdRV3ozCtnQIFUxXkxKkGzXJTNO
XFfBLu87taBoY52p5G73iuldAxpwk+XBou6wOiWyIW86HJPMyj+OH53ZCMDV6ZAE
20YsKBw03TFdi7zssMLSKYg3vxv/97pbvMZA+1OGrAw440LL1VcuT4gLU0RLfRQg
+7WWwl9Ff8SthbQ5vzTN0PgMs1TYl081ZTMcPk7PmYCCIcAnD6qZYEkKDnruNCVc
3EAoOCepfNQd92ubp69Yqjaje7oZ2yndOhYxpRSZW79Z8xCAOWOkda7JN+GHz+Dp
gVf8CUffrk8z9jjH58JFyd4iXQbpvS+hHLWc4YD7XvqvVQHsXi//jCeH8eSh2fjk
rWqP2z8BbHcMLzj3cvTCazNdnQGERC7oK1fx2+/9fQulr4uSihhFut76TXOlmzNH
3EsEpNJNDIowhJ1D3ZX36pDKRQOiMMn2aIXMu9BntqBW3wFTVTWiP0ejX902Cwk4
qHkrZ7i5Tjpd3Q0q0+vVm64hZ2e5btdToKiiyPCi/JlThMF9Ud9cF5C8bS4rFRbU
xbIDoIXyC5amlEiqtbzwSLGd3CupZ9jL+USyLYrFoex0oqE7xviuCDXkP+Jb+t23
BwjvQPoQ4S1/5ZWfsd8KsTLbuZX73k/BVf+9bLUOKfcbZfPbcx50DUO2WxYWXIjz
87oYTNkZ8o/G/DFw7pULkK4aPshy16JJuPfBTX6ouYAm/HGrpgKDAES225Rpwgh9
B1K/K+1qfLKHpCpXnugjEn4Q9vjzB5PcHV/vBVjnioCRrEADLRBkDHKI4Z9ivsYN
DiLLN+TkKpaSwwS2yyYTpyQS8E/iHQStyLBvMUV0f1nBPxoJIV5IGo/cdPp6wj8d
IzjVdxEh7uD8m5dLVXV/BrVgp2XsoF6NkhFebWybno/F13v7y5pf7U3jJSZrMADx
lQ8PHD7jGyyOjT5Y2D5rKQSB0BMreKbSXqV8MDvacYrKV0KJKEo/Xvz4lg3YVwGc
TVsG7Kq2MzApcs0iQl9KEe1+cXVzoJXk7VAGZmkFF8pIB3Ek/nbk7EiOQB0okwnH
ykc0CtF2JxpW7n91NxGJQH+TEvqk3Eq6qToIU66tmauDy8wntcZkVHlY06RnSG98
Qta8CwcGCAF5sETrDp/92+OiNgwaIWktLJqxte0SlpTXWdR+DSHKHqePSc4KmBQi
w/M8aBgxJ0xQ9XgrOn6ivztHFmmvu+E7Rs6VEqJcDyI8hDsGBHhVvmjOC1ikgzMT
euuRDbNdoFBqo92PfD68M94XjQA0D/vXKdDn0897K+LHFAao6Aw4hl3QS87kG6kT
WKC3BBX20GUGwt+PLl+ljmMoYO11FhJBL0mssT5opvCvnBqOTI3hQl9VbeJvTkew
nGf1MNUwk4a7FsAPLYRfIfkkLnwqVJLmRJSEOWXyNirnI+HHn2uuGvbQBKTDizRO
clcMsJMDofWgYzk3tke7PcJ71eVMp7b+1TU1BwddZap8eBIvJBQz++vTtnz+2KwM
xNuQSuYGCy4Vrn6Rw7XB7WLgl2QYmmQYay8wRZ/Qla3pkASgxYwmMVK/nEG5HHsn
Ks0QDoXoaLphcp94/iEAueNd7KlZ03RWxdp0M/RlL1e4KGuIffCi/Bd+5KFk5aRq
7ROI4xG0h0mmX0BWxgqfQyS+zfH7mlfTjZWX7fnpIF4q3oittyu6DVfsqH2lANL4
gXa1juGeGayyF4oQPfve3mPq3+qOCiiVO4z2Ci4SRst0DrSEa/rNydIJ4fgUQ8/a
X6Q6xwasAYbHtyZTejsMzsk6Vs7CRUX6BmMz+nJmCm2FZvcKn01BoCXboanvq3kO
VmHMp9P9RcS1m//EUCyzYbDJaUroecWrkekuJy6gy7rJIXKnIYdpajLac9aIcwz+
+xHLmeCEriXr7g+1czp1am8940i70EY6KPQgnOiSa/dA3nb9yVIujjIXA91+kvMs
1qKzho0z3p86jOhAFkgS92TkHNE2H9uGpuZT52yaJAmArgwtnb8d320gWIIGy7Wg
co6Z7dmcj1fybBk6+OHz7VZkAaoFeFytIqL6Z8XdO37YdD0Kr53Z5j6MFx3p/AGG
iNWNM3AoEjYQb6JlhG8joS6eIuq2yYNd6Bg+Sq2+T7ToqQRuHo+CbS/oIyL4OTng
rVhAw9Y4VMMpPVO+e+lCK2U9xaatl3D60f+ww5JyA4jfp9mreYs/k8kJOksinVh6
jBtTLNba/tBfSomvqFv8y5p6+nNabJb5RlT5ypJtSDWAu/gwdkKBMeeVslBu7Y+j
bsNTrulJ6mldRRKWPZvl5UvOYoR6DHGK/xvffGZKoq2rSj7wJEfEfIFkj0BSIrWW
K3dpqa9GYR8cxp51KkpOan13nit5yvUJ4s4T78goPCTKVs3sla1ihGjtExdGqT1C
T4ms8mYCUxDJ6XUDxVGuPyTbFyga0h0FnYbk9rOPepe2dFn6jwauwwzjm8KLd/P4
Vk3n6Jx7smv/5nn7hrUWWOpQ1yTM3+r0NvIX8HEx3UlYrArfCgjxUTfXy1B5ivgv
4vJf+0MNYxXu3BEDIjC/iYyk1HQTS7n3rnffzj3VJ7rZc+HBAZS709hfR8FxuO2m
1eh6nD5UpD52kE6K+qfv0tzURZCfUe0bPCKgPnufmyF5Fdh8g2vzgHpe1pMAt6rq
SKzTq/UNucaW0xZ/aLFP9fmY6sjqHiTDxkD36DZFfbESWq/7KAm9LY0EbUGgkE72
VPpzH9a7qui5G/uMx9ECtNJiGq1yWiQA04uwH7gX2GQTwT10ITc/4c1di5QqY2hR
W4ZQXoM4rfADW16jXT5w859d/NvXs7znljbgfVwnjm4WDmSW/xsfc7bWzQNclXXE
Iae6oGM4zDq4Bt4OlS7hw1+A1Fg+uG+M51YRw1xAdc23elwK8Cg/1ozqgpcZEEEh
Q91rWUxryYyMqcwbaFNUDp/RsdU829GIrkGYJjiq7b8DB70YHBDohQ1/dCB5WFvA
yLh26l+52VysuY1kg4+y0CJJaXto7QuAhgCV2HyvwK6vDBR0uSSu194DYIw26emo
pCCm4HRDLD2x9E1l5CgO+xI2ytvU0Md2U2TYUgKmH+4doYbAVn0cprTlIYmpU9cV
Oq3HLRP+y4wNJw5zsxk6YjXyexMZBkTxHUtbdJCvXbiVfr9R6Xv4vt+NyjpmBqFB
J6OSe7mUI9LHor7K4jxsvtHXFpNg0sN5L+9CB28wnS82XCqF3qU7TOvkXuyR7lYr
cDU6BK+1AjtB0QPL57wGnC9GyrqA+6dI0Fu3p8jhvuN2WosyyEW2VvW6cUCTgfi7
DBZJvZo7XAIjIVnbBdaJtmtQm28CazpvX3zSt43geNvxW+D5MMv24MIBOYA5t4Xk
FsiHW1hmmvJxR3+vmHKqdvcDJz7CHxTfx2C86dREKxUqJM51FckpIIyqMgmHZmD8
qJ2jfxzlPkDL2VAnSLTxacvyUgpOkjRWN1e0jGDE9KnYVxRSfj8gaIa9cLWfuPV5
QZmhguc+xOz2z+UKiQyBdv10nun3Td1qFFdz1G09CfDMsqS6naWWMU6VGaiG5aCV
OcK0xlUAuL/SjlHM855WNP6lQCRRujQObZdWlDtCjfXbTtqWeKPPUprKplKV+RFU
WrhmboTzuE2DBIhjvQVcIZr1ho0H29m6SIJGNxjADHy8NXfk+VjbC7iDvV4Tk9Nc
a3UJlUHT803hv1m3egp1avLhPwPsN9S8j2EbrPLkrTbyOsMc5z6ogJnIIVpGzblr
BiR25Pl7hahwRhKRJ+MIwYtxI3ZiSg3cX48TWcX+XpiLz0aqQfO9rS6iWqs38slz
H2GED1YR/2uVPruxlkF0NNJg9HSdb6+zfEBSkigAyxA=
`protect end_protected