`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 10880 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/9huKRhRMtvnNqb3Z+UU7TahEoHV+T8U3P3ufru7l1O
3DlgtZzb9QxCbOjthp9+wDkjygH0eUfDrEl1ovhZG61L5Dska56mP5nmYufCCL8C
Lq5E6twsicYP2J23yu0Euh3KYymUqN4u1GK2sv4Ut1vTYE223VzjFqmoCwy8izfO
ZCBQyw8j6rmsvfM4wABuW7nQ5lgJmwr+R2z2gipg4XXenrt37kGhUmJAnNNTAMmQ
9x8UlI00G8g+xpb9m9Zg1om994eU/D7feDiGIBn2UTy7l54OEAKAoqLtijB72Bfp
8HIdvNV4Cg7SArvSZuksbpbvd8AHCqoV4OsH5raJa4zJHe9EEERdYcwptXES+RgR
oh6DsTsfpkxs/y2ztpHHwM8Yx6AUa/8wyPqckV+vL2TDNwyMCJPUGtZSYEjsMhhL
KJfzQWb9fCFWhYHyvYI7Qrt8108ZO0YADh/grfOs6hOzqpuXpQ5G0mX8Bi2OSFJn
1bykpYieUoLKPcbel5O2S9+a+/s12au0Gs2BxTluXKsWtHjw+C+KGyzYwwwRK1Pc
/mVXgTIolwz6bYpBnyLnRy/f44yIBLyMnCxm2lDkSZnlxuGUO+BBDeem2RLrkBW9
rGK2YzIkMG0yiVjKDh2j+AH+r5P8OZ7FtkiUnNdajzKl4Qry8XpC33CzMjjHlqsa
i+RkMxzIxFlWAegc4sNe5iCRAjaGG1uSCBerKB7uGeoLzNup1owqMvH4yX2/FRIc
j3aQjYFUEhUOcTibcjsruWIqnMG9XxzSjIrbSCQ5i/nC78R4kikh+fYNigTYyfy8
3CHviyydfZLM1V1eCg7JfJBS1HJEunwQ6ZRffh56+XtW+Z5VjwG8xiAE/V75mCoF
/0Mna+k5l5uFahNqF9I4VR2bFdPiEoEj2KqNJOq1LxD2mlSUg+OK7kcF9EAxLfYA
rmr0TUaI0aXH7Hf6kuPgasEzMg70r0lTQiu1+mq8R+girMtR7csFXoiKmgEmn/ss
H/k2kJYYiEvL0xgJiCO+7Druw+qa5LpJvj58DInZNEtMAe2mYJzRkJnr3ImLha18
S73JJ58HRij7ULRvp7GuXQG8J4BuNVWFRyAOx++xp02y3rWt0/V+l/s4f33VoZzT
RgsA40PmxukLFqK8L7rabUB38ppjnmXBPD7hMDvaCTFE1Dq9Iy1MEBO8jMp6Bbp+
hkHXvbfIxxYs9a3ucxlkX5CcKhNKEKkXfcHmV+68d0XLiGQkLx5ABX+85QP0cyPb
6X4BQ2hwmtliNsgVreGn3fcYwZzsv2pWlpF8rjJk+SAkB5P1Pk4hRHeNIDksKYKF
i5D8/gZUFfaXJD2Y65ZbGHcKxCmk50WuthTWuWGnN//ZJTvucPPqt1N5fSoqpKu6
EI+2dNK4UMvaKkEDL/RN5VCLGMaY5sgn/eH2em3HWpprXfXjWezM6ok7Le3rsRK8
eZSMdv9MjnVmt3tNdTc55mLg2Odn12Owd4a/hGP2/IcDKZ58KfYeQPUrx7cQZSAm
kxTSGGFo5LNeyrJM4oD9p1ciz1vxkykJJbU+yBsPDx7mhSLAyhB8kkh8vhlKmMW9
NHm3mrNwP0R33QWEGUYoQ9rY8hMnLDlPi4bxY4eGgkwhodiXxRJ17T+PYeP88g/+
EonK+ZyqHodThyUuoq90Vn7msPwx1tohSjNL7dPdtLZyzYjMZqsnQtogGZms+fyv
X3B+RuHVHgkLcT56robc2r4REBwX6w1sb0UIFeofKvuL7mILWea2io+vBX2KNSpG
J8r/5hUn1Zsl59mvaYLTicAtoW7IySAaKXOs138hwFjy4fiBsD4kR6iLBAQkGBWA
KRuvnKwOBuzt3CAOPGxJVVugBg3QU4xazseTfDj9n7w5+Lu4zkpsihXOp1aTAQAS
RbVHlXHdUQ+iU16Yp+FXzJgOLM0Klal+QwagQpL88yo5yxdpHOazltlez0Z24KOW
VNRT+R63pecbm3aiX/sxv5EgY0cchj/IT15t1ZRQKZGpd3y9bmhw6niydYEZi5AD
UBIi7VQ1ktgKI8jvdJgYtq+TFf5ZrSBOZF3jFJPfqllNysz5DAUmtclrAxqzeJvy
dLomzuKbbG+Er0bn2ZD8g0HtQvZBbOsHPuAtFmACFSMBZXH0Bw3jOer0+YJDdo6q
QfBn7p/nu5TeVXK29obtAIv5Xm14vHc6dSyGVnHcRYocRQddmHc3QzjyTXzEBvPK
pegiho79q8cc+0/3BXwM5Je6hcMEWEvdI0gj10fHxQE/Dk1M1dlc8QerRhUVI878
fHxMafAZf9RPzT79w2C3hVK/9IbX/o74gyfLojzezEThcvC0nwl7SPXF9vpznICc
svHJq/Xr7YniOzAClqBGABdKQnn3hFeqPOxPxhf923b8FBt8qfqjqgSpMMflwwV4
mNzTDmLf1TXCjLAmQWEUrn5bYgCjRZF5aPULGWboSltPAmRcCH9fqRK+U0HMQG27
SEKz0Dz2J1JZKI0VEeVhG0BmNqrOUPP5sqIkjOSfS4WZAY4oBAOpoe1HWjt/aAAf
ZGdSH8AgvBY3BaPs3TFI64fTkQJPTNq9pQQjXnpqyPOVtfVQggzlkUsrfWiSpvh0
J2M88fv4X5jUlZVyYO/lmN3o8gGwseZpiyAfK/SAVO5p5NFOoZmxWq34BCjYipxm
tRGO2iBk0H3FBGuTaGJgixwIB4kyswuOdRoVc61Ir5mmnL9P4vykY4+LJC9Bho4z
Le+zK3I8wBPcHTqOdkr4EDZ7EoP1pniUaJ0r+0qeA8RvuH5Wn9NGFPJnZcZrHETa
4zxhmQgxFW5x36LUvpf4sq21bVG4rhiIoMFDGCYA+s0Z265jA4R4dLB7IjkyDF7k
ajBGWkrYlBA7Mqxops5WgfL/1I4FTQoevMClmmatHVk87YVu2h0bcxgxZTJWVc8V
j/bgFHamc6qJjJjf3QYyaprNZjR49m8RZagjm7fb8/csYhiAXe0c8cAy99+zJtDf
/QAAY8luYADsEPNTHaBYTpUNmrcxjoYBCJw+6kqJjqiQIGhtHYDscRdG1toxKimq
ettaOb7zNyX0aJKTwhtkOXpXx6FLV203LndqGn34QClRK5AYwrvw875Uyoh+Vh1j
OqZu5LX4nAwPJ0Zi8MtGCJiR/Jxve4PevxXuD0+yP78Sfatb73dTSOSN71Kz/cKM
7Dybya26hwGyTioy2bOD4Ctx91GSkqNGkWNjiNnOxUaEIhk5iV2W+4WR8FZh0Qn8
+54E4AjZjGBhRqfjEP6NbHikxWr82C/h9nEM07OCrh7s8zJaAkbVAnbp8C/sWkQs
HegvgF7de/fLEZkTIfSBgyBtxITvCJPVRF0KblgQ+b47ogRSOR/Eha5en648Zi3C
6JiOSJarsEXnS3+ujlF8DBVCsq3h65wlEc9qPvccksAUXl+6BlO8XUUwuU7Z2QuN
0mTLGNP77eKJl9cAy+atTIE6aw3vPVTzFxaeBfq67kd8YMSBHHlVyGyZWFJVlrh4
L/7i5kOd6VvPWyUORNzVw1x1rjkM7GPhN9xGGUZRoIcLN6Zo9oaDZB+jJf7XjWsR
sq21hmC7y0nxsaMyhLrhB7W9SlwmIUBRX5oFfKzWvmMZc1BBmLxcJ3U8yvH5xoRr
BYO+abTIoKk39kRrjo8JQn264470GF3m1HA8jutwJWn9AcV/0HoSJAYHxi9Oxcb/
snwbT5xV+obNqE22kjGtkRqXfuHUOZfvP5SfYAyhydsB7yFlLRD9zS3XOGVnuDoo
YUjVXVW0/eJgMQsggiH7ZLEUrAoRLc4CGe71pgx0Gf0z3EfqhydTSzyzrJ1ZhljA
vfVYan3ZBbYwTVN1dS1fktHPUrN4tLte4PBzelbnosYwRpb1Ha1Cbwc4wiSxOdY7
24NjVyhQUlSpsiF0bbB5P/cKSeYhq6LzZVKjZA2OnrfughZOAlyC8/sfVKS1YLnW
E4kw/LeDm8O1n59PYtP5u5RI0XGCPB0qnlrNTpmbkzOOV/BXxPAy/FXsaWWn5Zof
3HLiM1X7FJdBXrMsro+2WgnlGa22okpNsSeVUpI8vSIbo05jbvfTpM1Pooc2T0nB
WR96IxxTBzhlbTVwduM+ryp8+jLCXeGWsY/NycxHT8OkFkVufjysv2TwLedqBiK2
ShGljjv6sxQvf7JcbTS1CFAXr6fa7ZS5YvdEZfjlOK4SdlQUg14P7QwbPP+EOTh4
EMo/fev7Mqh4K1/u9SK8/uqGyzAHkUrmHBuuG7wMKzg/Yrj7O/Tsqi21r2ZbiPKY
6KyIeh4B9QrRD0eLz9CrNzhN1F7Lk3LFJlKNJTn/aPl2lMo2Fe9yuQO++w800UWm
O8CkP3bR91Z1qZv5mgBB7pDFugBFqvr944AcWikZ/JGZ9sSKC5cPKWbYNwiFotYU
CHJUeyQFpVROU/ApukWGc5CfULIYwov44xg7oXas/OZLq3116DZPEjWJXofIHLKU
I+6nRt8kBeyChScqCyPyxltHWH3245G0X9iQ916P91yZF4eNFs0dEn/opkIENgAh
814bk5hb37KW2P5e0GV9J1CUdg8TdH3nq6XsYW9CQWWn/d6EUH5q7bs+ENFl2Ex0
D/XfhBuAlmkNjLa8QHYcVvwekFyGF7e0NJGi4+Up/+PPsTrSgoLy8Uv0UH5sStbb
36t6b1sxC9DE6lwcnMw4Z5Wwhion0XADwiqvvI2e6JY+xgCRixEtM9+JZvfgluuc
ZJPLeIkpwM3nTH6vQ5rdussU0vam+UpVljsNa+4q7A93fa3Tz9lMPe8pe/v46bOt
tHrF3jLaLWFqwKbEnsNXHqa25pu8XhE8CmXNQAByRPZQeVvxUebfYpcopW/jtooA
lYv/4WXzC6MVW0/kpIWKTjW50DZoQcSJCusnNwS6g8920SE4Em/ZMu3n9mZpJuCt
dnLGdGKzFj0NxGdbNy+6oMO2X6x+3mPsNkW6YpGSs+0DEm0QtTzTqJLX48Uz6rmP
DR6uuVsoB00Vah8k9KrG35AZTCugMsFeXADQo69oRY4ez46gbUIGVqHpfMaOntLJ
tYUx52tgVMeaFu5Q251a2fc/goMweoR/UhHUj4P31b2ZszgIimMeSNk9fInEVy16
emadBSKQdaCxq4d/pQhH5EogEE/A9A7JzCgeOUXZGRwonP1PoFIZ4prMxey0XtX3
qKqiKiYe8eEgVi3Gx0PrJcMdqXtgINdhLoOIMk+9ZC+64hTQOkPuzoxbWZeRuebe
zZXS2LVl0/YAJd34ZnPL5EcxiXr9qR1182EULT+9j2HOzi4cHYJTKxtZCd95L6yO
XJJBHJF/tir0OzlFb2LG7u3EvK2kB6J9QtbEmwvnLlL9uAXUJhm5M+AhQv+fye2+
pWuqpUb2sQ2L5BZeea/MylV9FCVzJaetBQPq3WfQnWIxmLq4SDIM2XrF5wEqHJKR
hJVRIyiraOcu61PWnJ0Bq2N4jntQb6jEy+cTi1C3Tv/zRLn6KDfeE9UROsBhkX4D
Pq3c2B1vzAG5ejHwp1oQPd+Y5wa2aq680yHdHOVIRXUDh5fT+rjQXZgVYgIrKirp
6bpXp3Ndd9IWZCYSntbiivsMzdsAgHY05c6S9U7pe/n9Q2y5nIiGtqMsgvomRfKh
7cr1QicEY/4HB3VP3KBVj1enmWrOkfm5WO0I8tA40BkhaGOogt+iiIhod2lW1hSn
7XLl1OsUAE2oaZPNFrNq7Fe24F8C7WCi6ViPVMWySsx1Idx3+ddc2vTtpQBnYt4N
HkIUmtVwIQ2DUA6wIYOqjAkxYwJXuBGNuW/dKP5Luj0f3IXv/NfiOV9mH1M1g+0L
6yHx1sRs1+JAlbWyALuHs/Sqmsa/w3cNVTzgVt+EpGIGmUSpqqljoneqd/5TCSvY
9ZmLt6rSBo6GscUxrk/5worEN7fUlA0LucShdZF7CGSS6zSwSlRZHI84NM4488vy
U7A1lfaJ726wBMxl6pyoQtEY4H+FjXzYL0jrz6aCzhbKUZuDQNuqsGnfJDwLbJRk
a8hAiitmTTnR910V+rValxC7Sa+vyjVw5xVgvTp6unqeHrvaKDS7m87y3MCLaFCL
ZFK/+bqcszLCCoz8dvxro6pa6m+jp5b3qJ8xXDmHiMJtMUPE+QlhvqULtP8+C25k
fzzjY9ZLo+y1Zd8x46J2zReNzjU299RlQ6CyQ52w9ezoOkV7jOIJkCDJrUZqH694
e5/cuMBjoBgHcEnLRXpR3l13yNOiIaCYWVBYeHgWN7izrHrDfAhUh5jwDTF7MJNh
cZ3pNQ7xuj4FSN/Z3VA9XvXVQ6keRxGegfmaf9meuWWPryP4kNrFmBSt54M+sgyl
TJUKKEBKzNnYbcuoE/+erkh4kXZg/hsRK0t6r3bzyc3a07kZooKvfv9ezhU7caRw
eSsbPAmEFbkbkO9Mcvn6JAXwE/YFn4rdRp8TBq38D8t2ap8Te93mgZrWe/P/04qG
CFwVOM7hpGhFFvPQ/Ss1CWOPSWxchs9ZSvqZPsaawsL1qDRnBsmkYikaCpmMAFAz
4ilEWB/Qz6sfD7vUlAjM8xLz8HbUHzju9s33o3sNJrtpxIGkXMhkceTEcud9tcl2
6eDjOCLGgEKiQChUVHtxTlJNykGvoqIQcjzgLsgyK26TQSh+d+TXKN4YNheZie4f
k4GB5sKGxHJ8nqDp6ERSGLQRl8rXkww6ti0As13kUyFosItNkw/EEOwlgHIdjTPl
GsDqaYd9HdBlW+86PttideFkdJRv9hSZDu17rFfNfU6e1p9e9NcyOk0CyIqU6Bt4
p51ymkpEiFfeCOJlULnFBg/VRijcONjdZFwyET/7YpV3GKdvk3HztN1lNoRl+DPO
X+7HZX2+N6IBAhswabObOz11s7QHXYio9WFcZSiVwh54pT5q2RdjCRMIgwAC4Jwg
uOZE2MqZJFTOA/S18PpzbPALwuqB/U19ona+WFxzFBhLvOGV0wOaUeAfbcSvTnsE
wDm4wlno+PJyW+edqGoP4UdDb4/KbsO7uhSa5Dl30lIiuliRcTV5Do21gAx6mx0D
Pa8bdvPAaCkDmHvZbeM2ozK1oR6E8IO4p+eGG5d41kggYzOKL/FyVle5O3OlWrIc
UMHGBDbcJPq4g4N91hFRnLOE8Vvb7IfAcac1xK31hO8tntFHgEd4AsF6/Xl/s1bb
oVfp2on12hmpA+9HdNjcX2kqhEqwAwMNt7oyx90rWt7DOP8oUCzk51MaASx/jdCF
GqTTX+UJ/ft2BMc2DVs7S+GcCxfSCAmErji9R/RPzKYfvD4TmUgBwcZigsQ26XvS
9ixOxs4kng4N0DS6SLdocPz8X+EO+6q/F9jogHYCNbU0X04fjghsgKRoWJFMw0o6
ExlsibEuJC67umrGrKATOux4JFtfzt0B1TQDBmYAwejPBuRPO9FOWPtLeeUIiRBy
KjAC3BXmEVF+4cmiQigNsd1YPDwlBpv/2tUeT97+KIAJwPQY7heAB3KGCRncfqi7
VYwbyDanrhOg4Wk/z+PtJbJyAOi12iTbqJAXfVP3CpX8x1GJlul92214Bw8sWrEd
1KR/fUZqButL1QM1lvT53gWYx50EuJLkZM8e9vXeZYxbvBzWSjVby5c9yPQI6ldl
gKWR8xWXTFfhqNEh7EDUrZ/WTi4T6PcbzzSGkzVYQc4iGQC9zMsnn+FVeEmzkw9A
8F0mEWaZquxiuvN3o9/7CZ5jVNQsDJFjZyAnr2vk76QKSUkeIBVSphjjrW+/Ky0o
Vo8Hln73DYBtZPnRDbv+hs4wDtRL+pK0HU/mZI74Jk5Zf//Nhdbe5VkNWhoP7w4I
cFYPJitFsgdlmcx5kJHKjsAuIRro2iXzioEJ9C10b88NUfPuPHY3j73v3/sE+/7x
VbEI79VNJjlf8o9sfbKtRi5O63ENAu9SmQIy36+bPxCPU91GZ98NhUpDiijjRl30
Ma8oJPP+ksgm/UXU2ByEID2yq0w+8jzcy+kCpLz6qey0SBAiXMMykWr2Kp6OiqCE
ilGmV+ZnTKUq+4bncyd8VdJjvI6qVVVp0kGhAkacNQZIcP4h9hCPhVqTy0lkp0o4
9SGJGKzPd9tNYwp9syVslJNgsQ7RnSRPkxzHEmRYSmqAkYhLDBduBOcdKpzTRqrs
gmSGDgv04ck5Q5D/GiwvxTqK+XArs3kVLwQ8znjtszn1BFFEeuBTst6cdfB3eAEC
iq5f1nzbVhOe9IAheunQtjVq4btdFcB4GC/MmmUiXg9/kP15HBLWeIfcebXYjGu/
7GF7DEnMXAgRqtfrjJrsMGJIIzpjMaRsV97z1c3yipVHsHd7S58XOZf/00NSXZCj
omo3y85vgwKB3TGSla3+VmFbXGCeC5hC15EkQC+c5GNaAijaALMy7rNqCZWUXGT5
Rgh+CRrwt/92vPqdt1E6XFBKUiHG79xhagw59Mg3fRbPPJjcSiU6/F2J8u7F1BhI
S25y4c4kKFKvcJ9CCZiHHASvlKx/Ml8yyn08Hrp4idfImRXL4f6kXHkg2lgSSs7I
JIZxEngNKU3172OTbSZG3mxfFJMeDgAefbvBSjCmLQhTMvKvte1Q6qhdMLEksUC/
ZpssQ9noF+VrqGHFQQyGKtIDLEbtRBa5Yr3gGDSGlrHEvI5ShNES6QQ6q+8RB36y
L78TEVTAQovx9+j34KHBco4tEef8X7B0h0lTpTJWyTJdkl9h09NQQAMC1g38D+3T
Vl35xVIp+84aQdqH3bagXS1pHZ8o1kE9LuUXrRct8RsfHXBFIl90EVw2786FfJwe
CSJ1vMNdOZ9lBKhPcLI/I/25OZ3Nl7tycyKcVBi08PlPiPHmNJ6FQ18YURQ022TL
Dt6sxFEYl/Ng9yXWHEIX1Kuhwi37iI9QoNpkvvJlqMM4JmjN2rccftA7osoJRWft
zM8+euDMDiDr0IVlhOkUW/BE4Z5D4gx0GdDK0+Ad64BOM0akVZ5+i0OymNanzdEc
ecjaqNi8HJwAur0MsG1u2T4RFLf4UMJctcbNokCSURvLW+vMHO1EAHYRV7Jrx5kh
uQACqujSSZ8zlAS6nBKMvW53CFx0pmOOUIM3OTILwin3wxXmwizvO50mSX2ggb//
CeussBf8Gknj6NONwMryvBs6jfNlLGcrgD77vQktM05CDn4teOoZSTPSAKtpH0KR
gX9/KePs5kMtCzRd7DmKxHUVeKUEUYA/rSqQIfMtmY94Ux7M63MVUKzA6GTfLtZX
cPdjj+BgAwoZ20uW3NJSegblTzqL1hjZbnCvIHL3KGiPc2jzkjzsjKibM4pgxfjz
sxTgLc5dxGtXTmIUz8JW+K0CFg8+BIcANEt/z4jiLr8n6nX4FDE1DyRLjM2j3LzA
UW8flSEiC/dQRfSI33r+HUdpi/fUPsqAT5ia3HGsxEHrlfq9pTifmB5+7m5xUijE
C1SKddtzjb2wmnKknxwPsQppeBwSRxbzmMlPTz7HfVs0hgPSt3T0Gydtb912m2Ss
2Ct1MdUGiHUb38LQxMkwjfNHI+gwvCci0r6q+6o5GzZEsSgYX5LZJDP/+bDjcko4
ScN/R0xk4hpm6Ah4k1wqPqE6cgYiH1jgjjMwVl6Fq+yklTYt9JgwpjG5W+7h7CxA
sz1iECXvkzudRH4h1PiLXwtUYlv0ZZ4Wx6OnyNYoL9hFubPz0LkXaK/wIPehE6Tm
BjRDPql9FqXi7H931Id5rJAlhqgpY6LKUp9BvQS5KmDGWp2RjHnhkLba3bybVQpd
dR73cZjzdlkQcc/usI75MR9xJzsDFix6Ij47T5STBoEc6WxijctPXFjqLsCv+HAG
YymL06JSPqs2kC48WdaVuCP0wNbvucBPHV1kKo0gGGRk2+MayuSkw3IshMv4qg6T
hF3g28tT9HrbVoDiEmFohrEKPYCJf9mTjJzcRKxsUTweVuqs43cTm9Es4wAITkhL
PGu4Ilx7RVc5SKR5sPn/YK3NIYxG1G9d7QY9YcdWNCHbz3X/MCu49O1R33AZf9cI
kpgVz94+oOZZohzaE68g7SRKV7RZB1k2binh5udWVmkL4MdYFBdCMbOv7tJgNkuc
uRf7UDchLkC9q9qpzLUfdJ8yHd87MUy8lrULrzo/phEY4xnp3sdrmtJeElXSZoO0
4PxoozuP12YBu4Kw6ko+86zvkj2gpFvyvzagli1ORAm6yZhfN1o3cKTR4wMtxxbD
T2QdYx0rejVMLs9uynvdu3IaGtyKNUejg81TSdaeXduqIVTdj1zFSgsVVuqQUuiD
1dFw6HQgALYMzNPq0gUxyPAcW1l8iHAuC9TUPtJH+DVKaO5FPPN0OsC8j8yLNTYe
t+UIvd72hJ0uofF8WrpYLmuxuwoY1Kf2UaQrRGOJ3axaC+77yXi39vW93EEC3Fh2
JRtdB0fu4rBpKYWkJumbLW3KYiGgUkIdbBZve2auigGpbyiXLqluIeM/ctyQi9Zx
Vgxn2JaTKBsW+35P/rzoRl9BkedZ6szHD2MXS5o/Y2KDVDbMyjdVrSnIBdOAJbHK
JiXBAekhnb+T9Bi06gKgt/tKkaTk4wB6Z9sq1YIiVeob0n55VtdJMiW+InGl3ZLy
+6cwmTIzKXSvk6GCCpnvgfrqhjAsMIdM0ZQ5PsqN1C7as8UUUwy53uOV4/eQKxsW
1XZ7xnTBRaDPMGT1Z4z8d2Ft2TdpgNsusr+ZpECY+B3W9wO2HKSoPYx/CtzcDI70
+Xvb2f7dz3CI7BBHY/skEuJ9O9DfX6UotNlFcD89aah/aXjGln7vQtcFHaT0dGLF
mSGCjx1jSB5fUtVUUJyyobu7Idgyk0TmN1z+3UxrOMNd+t2q6gidERsW8Zs8bXNn
Dmfv9ixdKtynO6UwhekMjU4XI1UseNNyVfTxsGkOYzqzxyPfwwNwocb+4bL9YYc6
ujt/QEDbRGADniuiVNbLkdlfxtqKz9BO7/ooDnvKATk/DWQricUSSZSz3zupDhGs
G46Uf3/BaL8yLqzMn3w1PQxksNkJKTUKYFJgcEuWgDhWDTCHRJ9tbiIRQ4CscQMs
C4uz+Du38SrI7Z3sfgzXOl80Kp8E9vyQerQ28Aumx9lrw1yaxm/FM+Oib1Yx3w15
5KFtBlm4kcAKKZrOoYoCE9K2hY+rZRphkuCiYy8KkKmKokd63lGguOh0DmmsGqnq
22A6+FuufooZCN1VGPn4onggFHTuLDuT/Tb50jdTGx+g8JQgqWX3uuEL2354N++V
eurCB7DKUiw6iKSF8ocOeTSp+nbg/Vw8hRhiU0OB9UQv+8jfOHX0baJJLUBimc4a
i0Bl2MFCrx5W3NFgrwfw5EtnQbTx6BiI1vxD6BiX6UcIzx48aL7pS26h3/keTF+E
rdyMqunyjzyKL35HOzWGHTG4JS4Mf/2d6Pbyi60CevlcAucrLeh9yMZbl5DQojB4
9lHY/dB81Lzym2jIDrBZfohF/9jbfzXCXEHaZU0WL3wkCIaabaqqcYnCNyEpWSeP
N9HIefuDoX8LJdT4Tp9nDohssItHrmZLpg56cpc1rGbWbHc7QN7amxEiEtrVnEck
YsCrHpxNH/uLayUxbiKdQ1v9qwYsoxKcL0hz+rhm2qFtd5zqFn7PcQb+lqMiXBxk
ex+J8YmwcTtHA4sNapKAvnsPh8YnadFMTtwPgrMqO2lAp2Tm9DhljrM+Vej4j79Y
iILIWXw1UWCldsmbmhQuLQIOF/ycnMBWGBe/4wSt2Ysb7Q+5A5Jr13OQFaoOecbz
3kU7MnKYfJBDE9V6L8uBofoZCI89xHq2lUJbLdIdKJJOHJin8k3ZngU5hZ18qBw0
/WAVoRNFUbx/H2eIrb67Dk1hbHVKZv1XRchE1IAYMzuLU32EckCIfO2SQp6kP5St
pkpBc6tON5rs3p6pRf6b4xXCnPMDHqaokcXszL0NmRA3i6dzkcP62z1vtlZcZypB
DldwZBflwJ4wLjCsvhnB9ggmV6xoQ3afj0E9CuAGHXWURwycYh6fr6zL5iZn8vdt
JRiEKIR7FzqAz8ORnQEkO8JzPqRElwEfyQ3nLBtJMB4C3743tLNwIsMDXW0b9DqZ
eUrpjkd0D3ea5VgzodGjy9x0hOjskV8gf+jZLWIg/EdQs7CAWP7do1UgoQJiWd0K
95KPNHA+U+UnJtcTRG1q6S18Cr1t9ohj8LPGmqf1HAUt0UYv11NRVfGN89fp59PQ
mOfuNSSz8l6G3lClxbyXQ5erIRo3Xp9lI9rW9JWf2vEG57Fm10SNKLsJKz2Xz7iM
oO/4ih8pKZ8lzMOxGpvKgYKwCuH+IXsgmGcxaN39OanGlJqUcFSPSPGRdh6w3phk
qocz9tD/BIiPwCxATRnadEuQHLctdEg2jkUDLgoZPrkKmlfAV0JrC94lTqNX/Hyf
W8eDdVpYgzp/V4kESYNBOcZjO9ICQJ8ns6bPAOPNYw86dtsSiy+z9+I+BWmtsJI2
/OeBkc2A+7GyBVieuaItvkKdH1keukp/fyqMdG6C1dmyk5dQ5oIopq/oAXJEYuMI
ahFRGTatx1sYOWRKl4W3d/k79FOjbjF4rvsxI3EtnhxmZ6qL2vgG1FKCerQ0rn5s
zNd2q9EDSsMtNfyt7tib7BP1MR3334T+DQezjj2EO8CHE99s7v4OTg1TYWKha+Dz
3kKpDjBflVWH4vf5PbEbOLv145aCrlEw15QEMY/p+s3neHLY7X7VKQEPOaIXZGtS
+h7z5vfqWqineMaWCMpvGWzNFvAgJuQ5P0uCMKxyUpq5cOIx5IlPUrmFREasA99W
fmPIVZr4qKDtoTIwllXhMcGL9fWk+2eQ+etl6va1Bb0WSfT0uAwO+/cp3KQhXmIS
qxyCKmpG675+GUqo859Dyz59+EthIKy5reRWizjE7LZcsdRKDe7OZgutLd8TJart
ekMPd7FpL77siESvARvmat2fwBWeqxfgsz8OI1G4mCb3NJeJ+a7qIo0HGjKOEfnq
lD/hMYNPDg0cXbXKIUOBPZXMevu9IQVVGQ0/pKal4ANweev6S+ConloXPLRUaZ+m
nGa1Yzi9rhvqfHe1EQ74Nu679O5j1XEzRxTUf0T/+/WPW53tVaxCzk/US9eH1Q5Z
H1rgDbJdg1o3Iqcu3ilcdFdLnNZiRQhMNuSHszvuiCOrKl36ddMLqTrETSoCuoGR
C1qmeRar24STxE9+zmRaMVLMU9KSz49ngbK50M/Kpp4LBx8YJl3pHn1mxWWa06SL
FkAzX7lNlWbYo6s/8HYsclk9YeHEyn3lwxOnS6flTmRSv7oI6GxvhuFiIX3F4ggw
Vh9dRsP7S8XgqtZUmruOwTzhDhEXVvrvPjI1zP1TjDPzmpIetTqbmjUZLbtzl0TD
4Xmsd2Akq6o2LI54cSJappTiyfn4tpA4T+m2ATRzR+awHYI+9LtrJshtDnLn4l33
NOD84I95QLc118RewiEajH+3uqFm/GFfXEtsnuToP4elgEYUePa++BbOiys2omjt
wcEdfUMP3EtzInDy8TbAGels06xV1L7kTLM+X6etskuCqOz0XXo0MdnpGpKAa7dz
kBT6CcsVGBQwyFka4Uueq3To8NEDwyxwrAPaKR8rchhLzvHgn3H48cBN8a8Q04/n
eB/nESmb8tE1JSfl8WYNWK7nPJydzIkXfIm69xJY0mB6t89ts+VRtbpIlY42u9eQ
SHbnDGrc2nHMTGCTv/nLg1/BBMFiMyZauahufuFxM/CYtP3xsPy9ymbVbyvRFgjV
GcfzhgCVujqJXKWKQ8HBv9hmEGZsdSv8mX1dN1pwQWffhRzB/fd67C1ZhnCR1ljb
ZKAo3Bdq5EpF+uERMs5jktc3WT0R+0M/hpFwXXdNDIc9sz7PMkYgbTmeopKHknsz
UusK7Xs6DXAFaUIoCaEoTjZqySkPq6paB8kTFRj+zHgsfNiSt5qpFBWK6CUK72LS
CKA3Eyj9e7PPTMUZHEehJlSJIHKXjjeayGGr1qMuZncJ1vU90ybQrIPr8NqrT0jB
cwTCAF0pmQ2XTexcLA10qf30oXec4I1zuqfvjTRz+Pl0XzAu8tVspDZSOYRfxDDo
Y5UoXs5O730U/o5HXa+l/sFb8cnwXCQIgkXIC0Q/sAy/FcGHSFxb+WGsPe4AxfVO
PY6FAXbGNDCoUpPc2Nx1hq3cpd8Oe/Ob9MoPjOqiBRlN5jtA8mGogn/5WFHL2A7V
C/+Of/wi/PHzW431mB6fYf3fuppgXNJg584hVhoZ7XjkcmphF1KbLE2qx+BceL3g
QbtU9qeXvZklJcyhV6pl5eA9DfqhqBHE3h99IH7TwGTXkgTpaA/my3rAPOdRKZ+k
oqm1d65iL6Hyskroi1JcjjCJARnw0np4mtZylbG00GON1DfZzYzLWT0/cs5zEwMW
gWKhTm42vmdA3GC2/fjNUvA42rsDXzxiTX3sQwQGrDQIusE9bXUo3cvKfXZwLrvS
KD9dEsWs9TsnwhvQ/EBNk6pdXhU//5ZSnXnbe56/2G8YZmKvZrR1tEsvmAWbljL1
ry6XeF3FEceB4Ox4hYm3rOXMPoo+T1DHyXp4wXVuYzM=
`protect end_protected