`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 2704 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/9huKRhRMtvnNqb3Z+UU7TahEoHV+T8U3P3ufru7l1O
3DlgtZzb9QxCbOjthp9+wDkjygH0eUfDrEl1ovhZG61yv++n6acuonw9uLP45TzY
F5qKq8p75iiL1MD5aLK+TrRPnf6AhUH6ydeJNZgGJI2hlom4Rn9VbktTtE9JNw40
cO+NIUsBOAALW4wd4fIoazM0T5i2+CV51ktR/eBYzOTLhZZVlaQ916UOFfc4h1JA
pU0OHD5QqxF/Axc5GjhXaYF0z3L9Br0PBZkEsSTaadjY70pJSp1nkqME5QlLAy5I
Kwgd2A4ExjNHb/b3cnog2n78qKc3RjGFgtSgsh+wF4Ud5y7y5yyzPgJ655XODgMJ
icIzPKiseH7YE/1oNi8C4PfmW0LNEnRYnG6W1a35CaQkXMilr05mPF0nF7bsGrkY
TZjR8GWDlZ9/AMmiAl7I21a805pbPKU5FwYIAXKzxikNnXZSwYmNIZX3XDg8gQaK
5MRYq2S0/52VOn9BDiH+/eCnLYINinAKP0CL2LbvDs6dCE31j5xyVP8NSmLAY0r4
ZtKLZNtDH/gcGrb6Zh4IRPD9NXHpBMpPV2oI0x8Dp06L//Cdy+OxoyuxFuzv1k1F
IwEdvzkqhRZJqGR3dMVnKwGROUbh/b4C/m6VZbDAgU2NroebS6Dw1p1138pAMPfG
x65I0e/4I81KvLMMVUoFZLrStmDNYVE+s6nRQHHpqhppwovVxCWjyiCuWonJLStv
NiF73V8E++JdF2ARuA9B4ncBAptP1Zo1wDjHvLqyR05ngf772VFJKEqYWls1LH0x
jy26rdfPLA43k4+aY92pbnnIh3GUytt9OgD2AdLszuuhO+bRBQfko2bBBhgv7Mpe
AHudOrGRJus1c+jxP8X9wFVB8tVURYifRjBHIIkeDdQSlBGTNiFQS2AeZDm0uDLz
nLNO/L7ao2JZb+TpzWGA2qxQms7DnZgvpZ4sBpuU82dpOzeabV/P4knJC8Wt2e6n
fnc1tOktdiZxdD3t9ic1jBEbiC7Waw1NAEewGPcgXWOYvY2v+cQyHOTR0JRLpGi9
GtKMKSG0kFraXTqlDHnttyN1R2KFuMhHJQ6FAoXbumnlpN2K01myDmB3TvhI3Umj
GrD5e9zcZNShWt3D+AyXRGTJhx5meexXKacno+dHEhrrQosEyoxWpJTjuQSlLi5/
JYdytFNFG8M6vQKKiifeRNePyv82jF5RAR19Mx77tAh5nrrO3JXh89+f/T4lfI4w
w6K5aQp+8TaiEkGACrQmNd0Tw9jprHu/y6nNSSc4QcVVCAqo0CYcv4v94lABHER2
Hhk3E8vS3TT/rCVS9cyhWsliJpcIiNsoV76nLdv+iuOv2de/3Agv86Krc9gt/z/M
hXrEGVITqKa2iPzVvHmxf8VJqGNEtJvCy3rDSV0WcZe9BlIa9yR50pyGAeKFyLcn
X1/hK5Upo9t1qS+PzqJPjjlcafr6/6j+WksashQK+muwtB2xrgbDPrlyuQ/YpLMs
8SZ5e2nFsXRqjwcKcvmic4i3ePwZ6nlTqDa6/X3BDxdZtyyuMLCgdXOpv11qLIxm
jaxtWxw2IlFyvlJ4G1bavx5WsT3MTVcYgys6X19B2PAGMLKPKZjKX5OM6SygX53V
BsIp0cZ7EEORZbg00MCtJvpLECh/0xRRRJGlUOzWCu6ehgOcUSq7Qjyk+w4+lzMf
Trnsjn11l5J7OxDBEX/EvQ49P+KbQ+sKFK09Hbgoi5oCI23dakl+NfbuyAmNhQIA
lEtpDtwgj6F//Tod/te3RL0Adj6OADE1BiUQ5sfd+sK2lCFZRf3L6ChD0Hbie5U4
toC55tz6PJ1L0b6bdxznPGSH/JVskwHWvMNVc8VSNWe/mpndn2/py9cJH16K0D8N
IBRIb0mNZhRZWaKoQeBfeI1fWpAizmcyTVzv2wbPk+OiH/6m1Fj5uGWRprRyWfo1
OayXKGWWw5UTWuLd2Q8UleCiQ7XAB0ZdaIsMpHeZXUXkRBWWjVdxPg+F9LeuekE8
SahqxEUUQsRfqEMOuSyW6laJmeVSr5Gl6qL/wt57M5G3L3XFx5BPzYvcMGYaNZFm
UdPgBkduCw9gZqCBNvQPceGr4eKptqRikX8BVm9qrg2dExLjlfCjKeYUxaUEmTsH
KsCFcFtUvh1lauh9ahBGicSlxXBudfD1SCKaWYHuySkBD7GNbAyztzgE+eWtDIbK
qST+qS+LPu97n+P67SG5kRUMRvwyQ5891cMUAmn+7aVD89POGdoGF5w4jezGz2GF
EBFGy/IsYHNs8rzOtXZS3h5xxrTRXzZZuD5yPpgK9xY5/Eypb05ZLq50jLIXVpgx
p1hBzB6QNuTRep7aajNqOzmnNqGMZ9lq5R1i/3tDixhh8o5Wgmzia9WIkdc+UJiN
qP4Um5otdBstED1SUVaKiRvIZ9kdX7xBkqjTWIuED+RLIicz/DtlIhp853Dcz51b
n2qcKO2XJpscGRgPIY0/jKPw4FBcyCPm+yg+XyxiErs+t3YN49IDKJK2VqQFzTdI
dF9DcoLeRbr2NZxQXYIvHQt5SKi+cZKs83nhpUlGhqAOeBUoOsv/yRmoNExwju4r
WfuqBH8pEnvg4IEIXWD6Emr5kyDDBEc4OSUpnGOGViBkEWgrBg/Xbd+FfIPnjLPg
Qod3c9c1IbLz+nneCu9EyM4LAVjGvDtpx1QML/VlyR02hpLKZM43/cSHTDrfsrVZ
bZJJCuZfRw5v3wIntrHidL+fPBnmXbj4JFmunEdhv0x005QyWBL4NcB70lWnbxbh
/jUD5XUlnYyN6OQN4gg1xnp4oPLPoBYdkFbsqxz/T4I8XEfI1eCWPNSAAHW8rQz7
99pOsdTS+7GU7Xo7fnKra2WvmOGZ73nHdGB0WR9u0EsVRZBGR/zetcSk1UiHvORv
BjUYV+PBo6vpHU0HLVcY+898nxDJHK4INJNtuPC16m6/Pn2TSbTR9a7XhzWHn69d
yBy5MDu/LcGnIOh80NAxMS627KEAg3z1yH4IqIoxjawHqxLGmhUl/QeSdPIxzUDp
oGHgBZPmN+sxMSNGYypKj6CVAK84pDMAGtFivRhNykZFmVYjyP5NY5bpyj+yd+B2
nbPxJ8hXlswzmgoY9uMd+JafTOONk+EJNERr8xpK0dZPmoN3KFQ+TnjfqhPuJ0q0
hy0Je4Ol5we2QTHeHvWEHBTJDZttj86EmKVRdrIgyxNbrloo/WKgHEYdSa+uS2j9
R8HVn+eWVlRHfwil4FJw6BEwmzASqbne/lcljfTztOGn18usA8cg92f8EqzAwShx
w8671nL0yKFiwJKKc25Lfew0v9/uKDVQdewr6sRekf1X3Ql3NjfoaD9+vzBZGWZN
CvDyNDrZrSgcx4uyAWeZ0866LqNvjP/C4CNU1R+wvjD7Zu63FbNGCZ+lkr9MMLYT
B16aVqNxbfcLF3yVNyhRmo43nLg9OdE75N2oF++8kogpDn+MrWWWUDGTxZOgipz2
Ulk66FWGYyPErj1WSC7+XiRfEWCS/zZar3QcQfVBkGDC1toTCY1b31KwbeuMWv6U
nWGpDGtlNx7XIJ6Bu/Dx2Q==
`protect end_protected