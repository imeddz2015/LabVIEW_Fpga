`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 28608 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/9huKRhRMtvnNqb3Z+UU7TahEoHV+T8U3P3ufru7l1O
3DlgtZzb9QxCbOjthp9+wDkjygH0eUfDrEl1ovhZG60OVutSr2mwucnVXNeoxT1U
dsCSLO46cMjgPdrhlbieOlz0epXfHuxfAt6GwTjU2P9H80Qc8o5aOwlF/+Xftpju
hecD9JqGboWUfw44ynFWdpPmgfmB8EfIQJmb7SaYnxBNozFE5YK7QEPqrTZrAtKH
CFcgn7zmAv5IwpzHHBvr+eSkiw7prHwSavV2rLyH4o0YqNnMA0lxfQcTH+CYqB0B
05OJ4/DIGPidMuE3DbGKmzNU98eTJlM6V0S2pUolR9Bzof/wSltaV5+L3wCfdFk3
tfSYKCWcUTIAl/Hi2dD3XT/1zYNssgIgGmvR3wCduGHv1O5i9Z/4+71R5ks0rybh
Vw5ua4ibEmvD+m50SurA6xrqTk9ciT1yOFS78UF9bLk9TpUuUDHL/aPBw17Tx5KP
w5OGe4Fd/b+fuXVR42umezcqZWYFacihxiB7EgtgFx67AqiYCqiIcp/R3BKFUODo
W+oWenTWUPBY0PsYmaWkIuGS/FCL0jrepGm65Z6a6TFBkDuGQFxlMDrbqIrOxgcH
DavqvDmdnTHfjJNi0oLTToxXUG8nvNIp46zVPfnhcf7YPYAQplVFQjYhV6QC31+h
ZeQl+L66+BzrVQxR5d6+P7dSAJ092jOWNZJKZCz99YOdHEZ0mmFID3eJMIL9J7M+
7DnJNJARyyUm7CmuzAXN2z3X5w3N9WQKLzuxni861OtvsY/zD4fc11D2kC5q7KK/
j+657r8pGj09MVcjN+vwgXRWd+Loz7L8ifi3xQW4Ib/5FtQFtcnaRdOY/yXKyyGO
eJxt/JxjJVX+2kfJPfLaJiCC3UrwKxp+rS0l3EOdbxmTcM9ZBWPkYlE4rUUrpFzP
K3jwlqsiy5gmNYQSReBdzNd9pstJ6FHZybqgNVHrpX+Njhiuc5bZKIElypARkWqj
DfYymCOU0U4ky7cvy9A5yqvH4sMQkWhzfKkta9z8aWlEnDJ9KrNcvW7njZJxnpAh
vdW+4sS+H4HA5tn9dFTnjKaArqt3G1FQUc1wY8b0s7xdPww0Jrg8b9LZeq6Ro3/f
QhPkzpZoDPQZG5Lauzu6GRXQ29pCqbZuhUatWNVybpIe8cr1Gy2eoz+0syThxDIk
YS7m4UGTCgo7OS3ltIpGYgREqh+IIpCrcOPOsHc56u3MTzWQkeTKxKPUrleb7ZWQ
GJGa+IR6HchYHOD/ePl8lj6TEK7ZeJWWyzidebI1rag65VlK/D8tDn8VciA1/EOj
SHNXJocNlVsUnPry/gzIg+Ln8PYMX3tST1SnXhy2jC2Is6dnPPOYb9frpxfaemwo
fW2O91VZt7sjpXIAa58MaJGuHsTDD9kZF7D1C+4O6ssl8nRHIayTpFhE5JSvUJup
Qnzo3QtAV8clpG7Yk6k8Tca0McyWsR4Fg0hDYitc6k3OcpxwabYzPidUDcmoBZ5r
yi5u8r8qVYqk8LEZpYvxBOentkhOcU9cQitrDM2B7kL9YkNPdxVGX4hW1LlLD34Z
rOhtx6ef1i21yaiUJBwuR11prpRqGOWO5fpg9qFwBuzhC2oadd6FK+KiEbugfkKj
oX0ALKiGhs3p1Qhg5BmfxwptIF2JfV82fJu5WXZymXsF/AOkuUHjJNs6FjDrP3Mf
sDSpnAo1AVq480pCITSn4Do/dG51VHe11XDP/vz7jxDuXndKIXU3QFrUc+N3hqkA
MbzAMWdKcjckPSRlTky3qHKoUicFRCRQo9wVNuEKEAlDba7vz4D1gbWjPSREKviv
coLMYGdItdBMTEvn5Yjjm5LpeNBSlj5Gks7YEK5FLDBMRXNL6QqAueoKnxD/3tGh
TU+qe6AFy0it9EEx7sSKzD11stK1spwSKvQivivXavzvuBKJUd0mA5O0waIgPGt0
z53BcPfdprNPKtxfq7v1jHPYey6IyVaQtTu+cYu9e8KJh+oVHpfXdVoVpovOLOW/
5vuAyJRpqFXvSeD3UavOoHTES7RD2AELzP9Ef5KCOmgU+gKIbXEqH7Kq7xjnohiX
j6zvMTu6KKHCyVhDb+JSamHJeiVVi9rjmsJSvxo03IwvdHsW+H8Ul1fSjjeWEagd
GnpVhBpv4DaUWgzyijPzVGA/jXfU6hOVEH4b25cW2GaMTOLBz7MNV0Lj1//0U9s7
qpQ6ahagtPbNHtynlXgKbKcvdBdPk3JEuDdKMQBpz+O8OZ1FRHDzhm13+E4nmn2o
TOd271GoMq7RS4mzcCEV/6c8sgAzayCfhB2iJ8OzHBXmkPWOFv2d2juFCOv9bH7r
rn62ckJe9GliRNqFIcmgquHquYmcYvmvuvwTMespMnD3bCFEpBSBpUpBgI6uJx+1
1od1IxIXu+mxJHL2zqFcB5t14cJyiWBqi4X3zllUsHHXsvzCoo52AjxSTQ+iRe1I
TsKHcWYXHttVwoIkd//ZAtxaB9DkqM5qFB9GCPdiqThu8STCHwrGVQhDni/Nj0nx
5zrbjE08tGaIVS96RtIsjccRs87qoHLGEQg0c/Da7AR6+Zv9SQWUpkAOmRBT1OWg
GE2PiosER+kblfvnVE38pkwqIDjFoLhz65VmpdqGjibdebC+xM9Q1TjkaSbk8kOW
bvKV7CnELE0DBZGqgGCoUa5F5WruMyyr6VrDfplah4pn3+kcrBa4go6eglQ32qic
2uOpNAgM8Hox5l3vt1822eyi9dYJx8VObClbNJbtPbkyZjhRWtFM/eHd9qXew9Fi
6c5dHPSJD64UzT7YV1OfvJA/xZTHU/7hC2WFKLLI/fHfPdfV25DJAo1xx9tlnQRb
tGzfoOMwuEcmLMnb60qei5zRoz+9NeZRdG25OHnSpQEMlqvAaNNwO+4969JwwQPV
6XFQYDZyTDcGoS2qCigIaP74iST6nHl/P4N8ZbTNbXE3B1otLSg4A54grCgqVvep
Fnh7Lg+qbC5snvdOuj4Acb7lxGu3iZLzoWTM/60bA+DTM0uyGI1GXRBjxCgd5hbZ
dngghlneChK0ODgji8rBSDDpicTNhvW2Py/2LE9URAOSOzmMpok/dLtnmRnGPYsO
58F/9wShsH7/BMptHgL3cldJp9Lf3wuqZQIlD42ATriKK9lxBLH4DVeCAIY8bJKA
3kUr0GYGuvORwiYWMQ5Oon05sAQ8f6Vrt8TvvgCOnfVlvUXYhk/HEfijc54QGjZW
2Lper7P2JvHyt9lVLloDD32QdAGEvikY5M6JxqevM+M2YVNp9RX+HT57DijjG/t8
DZW726ubiNR57aUOI6R7ACmgZ+ow8kq1fHBrmeNohg2eFFX48AJQmGX1IE9OqUy2
Vu5XfTEZCVfQ4B7dRF+hJVTOVKQbWNtsaIxgMNAm4m4LzSzU6I8ubPojIz9FKzfz
hRBoWpgYV/PV11i0CS9eoOB3b1zsq3G+Au1ss0pYsF/UHWTBkCiDCFS+PuXYmc6i
VgHioVTJQsl7RfKW+m0aKhcZrdIBnPj4CYI3DmqVgwtTQbeZXx20ibHltjmNZQBd
4LhqkN9kUAQcJ+t+JWLn6V3Acy+68fzlVtptkxA0kFxhpl+mSxhLPc6uO2uj54DA
1rKt2CAL4cenyU2MzvU0jFzVGhY+fSkP5VWQ/NJsYiKdBdQFQQW0kTn0o/7zwoia
lO8VpM+gzS03DchCl+sRJLviYssKFY1iaAGHxiFbQAQVQNSxL0eSHwYdkMIZG64z
7SpuSrvgAXWL6kBSffzofOBWFMXSqSvmFwY+ZzM4Zby4mbHMRYtQGQUz0zmrLbWf
VXSUPZEgELEkTU9jy6B93qLUg7PYZNLQlD8lfCxsGqPSKSVRkfkHssNJZrfkvkMd
y/pU2MbaSxiWcpot0z7Bk3TcryIbcRi59HyianqLvu4GSWIdTuvLvSVMakykCQxB
GbH4OQzvtdhBBDiJQ8hVn5VnbkV1j5DO9q0hbmiMXfSyVgEFuuOqun74XCcglIZG
Cie7HzlicG3JOATj2ye5LuGWe3c712rKGNpH7NNekukLI11Z2oOXgjVwH8KwGmCU
1QkKcMJB9U3gEdPrZs+qsVgqIRebgCyshqBPGadEg8NgUAaf/AIKlwHKgKFZKDg1
frzHaIiSI0UDn9YCuDnqu/YhVoKAIMZEMmxrMKjp7HbVjAsZye4N9QWLfjmaWdg4
pqh1xP+4xo8GVXpYxcK5sN8QmLqe6HJO7LlXeCGtK/m4PVWzDWM8vMJLTfy2Onlk
kE1Ynf8R9F83atA0Dkjddg54SvFpS6NYI3QGrHHDZy0f+JstLUsd3IhPWZ/NfkA/
wuL+fCU6o2WXlq4qS+t2mvSW/k5YznA/GYzS1ErrWUYwM3X5eRHX5UDBAlGvR5vh
mlN4OKFUHkK3Dq7uAJZFGnsl1RJXSq26wnyAf8QdB6ApcFC6fhyhvZZZBa11A4iT
bgPyxoz1WuYvziJK1w4nLJIFsuPKaWXonz/PQDgxs8Bd5bTEVm32jKifVfHWdR4V
CVODX4KSkXsWL+BnLEp1BG6+aM/JG0J8ai7B+nTcocgCrogjp5ElDXnqsW3yNsqu
0CWR5vIfU+0ozouD5kAyIbMEoPKm/nat9L4izgZ2bkozf2AH3tHd2MF6kwpyk+NV
5CVPqN0pvCWQQgw1S6U1XYHhZ4eE/pErqm+tiHPCwYmcGk2WuaayN+9tP8qm/ho+
TgX6HRX4DgoQa/CCq7xKz0LpJv98xb1lg4SAXhHviRy1XwLKwdUXR2hTbR6W3bYz
ZXENWvuVNRz9gOYAWuhZGxZOnUvrYJgb7FTOCoFoMen4TLc++foZTo3Twl1rkRFF
6T5uVCwirLHPudIsTO6e2Esdzy1QDhmmVZ9O/n6X6FCTzJa9W4n5AYB9ZySJ00KI
727Zspv96cNcFeFUqatjWbsLEuMhROjcE613kYBVDsehTM+YGiAa+onUNFiM4jIn
XIxLSwDlgXezAHKlmJZD2QxoS3HJ345ngJjolwVOTrqFHsg0HBcoqBBFAGKsCFyt
XASyxXCc3V9oXAi2GLdEHHYoLL3uDyfsv8oodrhpqACKJQH77tTgcrL9ybIZB0Zk
7DzFGCGnq3Q8dci87zRQdq8yBdQ/4Q3x5Eskl1W9sCMVx9kr6KxR20uFthRy9f57
KiCNgKEUalSU+Jj7eWz49Gv26kMrglcZSVLZl0zvdsqCZyDEm2fZiVuZXKfKiS45
xlWeSeq98Ok0myFpDNdEgjf17lbJtXD0Gt832YtorDNmAUaY27+elbmyoVXI+Hch
s2wX7SCuqzyjQ7QBO3VBb1dP9IOvTlytD2TZxDEkJEltEKWMp9u69eE052XhNERo
BYDAn81VB4N6mWiUkl9HtuujfVJE59OhTvCImFU/wFUdGw4Ok0H8XFYxyDlaYyw4
4TRf8K5rCTMOY8VoC+y8meD+6ViP6tDlS0xxpiSnprilFYsI2vS/9VD5jHdBMaIG
0gl/u3iRwuwIWCkZQTXxXpV3YLg7jj+DX9IaiV8O2k88/paUmMWg5+fXuMsIHNT7
w2+rBsTAEsnK4vHx1t9Qc0DrmxFM3mCAhjX+7U1lJQC1YF+AgqY3fSdoOO2rVoMB
yQ+Aw28kmuczm/lp+n71cIO6rIbNCrReaLEWN0tubxlBbHuidQUOZpE2t4xCdUTU
ckrT1CQKHcgfdVyA8kHwYf0RqGSmUfmKKXyvAE84L31d2JEf13CkmJLzOf0JQmBW
20ZUHGkbOWXSNAst0tfMkFauwihEtAUgBkWF8NB8eOV3IyTqXtHk6jywcVg9Flp2
ZO84kPYmXUU5gJTL+dFH8hiZZqD7hrewHVxuAzvfq7c01kwcKKVqBlNHZf5rCyas
m4FCDwexPgNPJHjNjbt5zKxaC2ewZaGuT68HgQe7ISm78DtYEhCcBa74+3ql5okJ
fH3BZ6P8kBY56yw31XrpnKFNU6krIp1zsUxwPh0gHvh7BFRIoYx4BcP/3fh6R/3s
o7/JrwJ8SdMLTrjJL2s8dyI6mc6XhfmkWusCeS8Dctv7xMX0cD60vODAsyJIWGNq
zketMMeKWA1WWx7fCKHr7uI3ZMtQyh8JqjUPfYdqt4veaTf0tvPGrdLA41unKFlP
yHyyMUxXqoUMFRmWn1CgRFNmRMypph4JU6Ejn9GiZ+VG7qeV8a4b+1zXJ4UNdyij
UghmydbzxPxeMpf5/oRp8meRH7pG0Q6riRhOiF7TxyMDYldDES9Ut2gO0K+Qz6jG
ZtN3CBG+xsg10+JpF57V4ozoI0s7m6rL1XRxiZa/vjqIajodVyl1pXadTjRXollZ
QVwP2iuqGWGVa+Rr3+u62DmV9mgWF735KGN32lXxBGswhjCuYmalCQlLskKlT3Zx
ouKuwQfOW/BkMRB5D6Ua77MAUEX3LM2x1wCTB/xVxd3CPLrlAHknObivu2A1//lM
ziE0NtKKGJ3KJ4MsydCIvQrl6HoZasqxzFIzeLDPke5X2a9pxIYemd6H82iI0dAw
jMh6C8b8W5N/n6ePlXg1fBRfEmXHGvSi0ETFOI8KTi8vAwDoRRIJQlvz0Krzyybj
gw2Aq7Oc8maJSF3+4RLOCk82OwQHBG/bM3gNrJ3hqstBRUnbVnkF4TniYJivsFv8
fn6QWCFKNSuSaFsggnMzOEB17sdt6VXkLYCzJNw8KbZFl4PjSUnPgzLX8NyrBpXj
3EK1HqRKxkS1vveKkuJ++FcZwwPymU2RfnniMV5KHEZY8qw1xMvlTyWjrET7+Sr9
Pm+Pc18OEyuR+Ks1+6jBxVUlryldOE94+R/hNvk4VccBySO/CNIy8QYBfvpNxEOv
nS7OW5FVbAZbCXYKOgwa7GZfBH8R13TtOuf6gpR8RTuYlqnFu4YiV4Cmp8JcsMBr
feAHZExAsoE68JPH44LZnQpcNJbOOH7Po4b5AOqluBC6w1U/KeW+KRG/xup85Eli
+ommNp96dnnANt5pSD7Iq8teic7q28JAcbi6ZRnaSN+qdFubu7L9W7K9Zpb1Ovks
JMblNWe069s/SdpT+VetVHshcxKWDmjQNzsff2VyPevks8EAv2Bdj0uED0Dx0MrO
xIORouN5tu/lP3nVb/Qep7xAQwVFMNTlFfHAbXZCi/RfamT7/4ta06xoFLHQYjlX
hWd1OZfyn69aGSUs6UhBZNn0o+sT8K01Tya1ywuBHL5ChwN6maT5WXmMeyWCtR1B
Sk0o3dSCnXJgD8smnmblNOgB8RV/PE2mWhgnzSvhNhaG302Q6QIwH5HejqZ6Hd0A
hI/aQRBcLV4RTpzJ2Z77+8OjtXN+AKl4zlMXAY6i1Ttr+ESsA6nZKQJ7YBIAZ7K8
koC3AXzQ6rpM4ogHTg/WqCSMh9gO0OKCgTpeSH771LhLOzWp1yvKalP8i3Ib6jcI
q0zi/ccFEoohyLL1jIIDE+/1TjCRerEYR7UF9hqj7xGxWiSZ+XskwCmhDB9EVVe9
CJj/0+W/QDd+ewKyhx06Zi5Q2lVtYg9x7tegwc9LfWKrlbmWHte9knkOSitNiLsF
xjN3gX5/07m/wG4Jvg7nQFgzgmJfIttkfVzXXmtBaotq+e0w0eJpUpdQGqjpKOXF
des0+DtA6/twZvRrEhJ20yYECFOQSLRZsgrsyVFFmOZCsKlo0J2WcdvQpd6VM7CG
fEGYLWSPx3RpjYAH/SMaZ438t/V7zus3L310sreAs/RVmp/9WMPbs8kQPbjXoAfY
tC5fB0TQ7QHHI9sLq6u6F6p17U2F3l0S+NEqykceWcRAHmegfpsnIh3ZIVHse8Ht
YYDJLWhSWMGiwRDfw1q5m4/MwZywrcnyySW6bPSVMfM5f0ntjx88IxgUx6iiEUFj
/11ETq3NuMT/a2PBP2LqjkiO4jBt6r4oPIwLYzV+e9bDB5Ge+KthRjt8Na6x2vBF
O+xkzfcN7LtKgiYzZFzD4Wzikm1MpcTombP8DCjERhXK/OldZHpb5gjBUMC394IU
1LU5RCx7AquxfFfBZ1JKxIWTdI1XvxDeHwPcLAvBU9fqk806vW5ukQYfKsFwffKl
krb2wvAXZXshBSt2guVAfdgDIinjMOi7UL4xPgdffyg3VxpzV8o2JQMzxM2C0Hz4
E5KAJWTxZTAjILuOp07XtF3aT49V9Z4OHgwDY+eOgOoz6cJPaqDfaivBRm1z8VkO
EwA1b8aH2M01ABOg0GEZ19vG9/OM85uVa08ZPOchfEiZRrZzj1/soHJs15kLate0
obvER+njw0e6G5MxZ0tUKedI239xXULDC8s1gZ+6HRXLDt4isgPmwmDY7yiaRE9L
JwjsvYFYhVODC/DkWw3jej1EEyAsjNN2hSFSRS+7gWynFxvI6FefcGZEOWkpUN39
jvQ/1Sb/Kygt2QB78hF/51nT068n62AzA0kv4ccs7DTs2kKTqKMBFed4C+P4HK6f
CafZZlEW2vvx5aHSb8gIUogL5KumNqSSHKL+BwPvwp5e2XIovG9dp3LyjgamnrQ2
T7o/Rb0azvkpGxZsgjfcg+TcPgbQdY6jaA/wHcswA0F31Bk/PQ1FDVoic+uUJbqY
4kvR8AF3FYzMOFakLDLJ60irp9pJ584HfcQ41STRLbKHzLw95H7u6qj/7SZx1WdF
C1EFornVRvQUZ2rzQM8Fb43dCQK0rekh3HFrjz/MEiWbNn3Qh9JN5J69oL80lI5B
5/uS7Yfd8gjN3emrXDALd/51DdT2JmD6d77UsBwHahcusVctQP5HYR1c2OQPpYFz
85tpzP1WTbgGdA8Edi5CfyQISa6SN0mCkgM3dJLtOqIQeHQtQOwo4WHi/5T8KoMI
dBfD2TgatO3P4cdYH/vOVx3dneQhnJqcNGtYaZ4jGg3e07pBi46QI7Eq+b3Uaane
vC2WP5LAD1RWzedQ7xs7o4U+1sU4AP+xDwq9Eu8LhSImUOu4CGXLxdGVP1if+zvr
Pq3+GFII3SMgO4TyK35fNB87lnqwyRhREnAI73DcOjByR4xCjpgz7JNEQhicsuW5
qMo87ZZxilCTSGbObZzj7I4jsXo4y1GeoXJPnSJ4gQgRUO5zghKhvJz9eME2zt4i
jf4dY5Qm+JXGVpAO6dZQ3/a13ui+4w5D1O0t3PMj12lyEL5Oh/YXX3mWjrKrkzgq
SE/tApVWY6buymyOKRuQjWXv9n1YGK0s3mwCZNQ8VEBQwNdx2ELK6UNvZTY1t9VW
F2p99F+Rox/Oo931GX74va0sv/llfmGM9r+qmwKU6dg2W33IohJQ4KXlNv6MJy9I
nVjYtym0Jat45YUg3O+m9mAj4pdqIC8VZX5cEZWDeq5o9sorDfWNt+KcSQYp4RGS
Eb0RqONMbPtJNZIyW8sGFG9SxUZ5YVrCXPY9GmQLpeRriTVnbxZ86xJxsqmOWsnp
6pCE16kF1u405TvemZqc/nabZvI4R0U8IcFXvsSsDsfkWBfwwxM1JgwzxAPcniLi
WHkvZg/m/k+O2WpIKzeWERRLiqxwGINtNMZzhPDme+k75SkygTI9zyMH6kmuorKS
ivkfm6pU70xZCT2qsMzvMwqDzr2p2BZ9BpLZWu7tagkTJEA6XyE9nP9DpEqI/SQU
wRkaWK1nqVSYPkNinToViYFC0Gs4bcwphlBFAwtVL05L0x3isjLy/NFwPmIk++Sz
74HvwB6bE1DEO+Pj3cLBzxFxjBpuSIBtekNQVfbkLdrAP+ITkrGJTA+ILoDJ4l8F
CCei6YuFKlUwOhJc6rifvuxUQCNJl3qVtXrHEEGXlgvk1xAYch8janp/sliqce2B
G6eglJX0suDvm1F7WRUC4daWypFRlTUOlhxNz9AaMfjqNG/Za952oXkPYihmAcrF
QZLHYQ5OAZlVyXGqETC/5vNcRA8UrudhzJ4P89Y1nB3s2ySluSniIRHd8KiuSOMA
Y0npNjvm0hNVc3OEw9ktohG7X+2V1+q3GgaMAmV8xWw0l5WKrYI5as/bWNCelk0n
S/ovaS9ZZgqY+2oi6PUjcNFZQc1168sfsL/NZI5W341lkP5sJzbbwAJHbikfekrT
rxtms6eDxbRKnnsB6qatapyA6qdXOOEIrlL/ngeLx4jwsPH5KvqMi1CsF+q36pd+
IuANco53fGfubb0bLg51qPCrIJmJjzNdHr9gHB+6OqFonmWQfPeSz16lG5R7Uf1F
yBSEhDJczK3q+oLEp5BNoZxdejO6Vif+S13LKvbPnmn+zoQKw/bqJpzW8mrHEx9f
LL2O9XtsEGDlc80lnwrdcZMxHLA0nn+79E9IdD8/BwB9YKIVrC3WRZvwt5M3kFn2
T5/gIslrYL3ShKH55tQcs6JODLpIOHNEPJnw0fKYdd9cufQerA09hVk/eK6dOLgz
j4s/4Xepv5NbzcxUOwMaNUuIPVpaY5y+eZyS7sJMcXTKq8pppwG/laz70hE2bpdN
xljnMcn/N2BJaIHcI+qE6E4+k8bYDXmIgJSzXZhqaG/XSi0JFvOF5IYWLip1erez
3QurHJtTo8L/UR7j7g/QFHXnEZxmhxfXHKkvtbzKao3TPg9et/H5Aa9foWwVIjEI
e2EWBSMZHfzFsAbRjUzIGASOV9FCSE4sDhRtOpGgEmFgajrlRnJcWXfK0wX1s+9E
CqNu1RVA7tpbaYCfqti9hrp/DCWjHo/Eu0QZaSOiK7fZa7NLAw3tA3ArC5uHKibV
qt5kYfLKhBM22LBhIITEF3YLOEWPsEtQEbaC5ffoiVxFcMePZtnZeifZ9hFvq55o
cnb7TxeafgAQW7p/opUMMvbXFcpRPtiSPYedDwMMX58/z8vp+Vkr33ve0Y7aRKIr
HERkob9wiiSeQ+7XEteVa6mV55GikcDELWlUwrvFCJiUXO8n7wf3ZdZR4dkyh3+5
N/DEqdu6IzDEzDg3noLy5Ce9bEvkZe4tX87yt6wk04xuRzbNgqQIfbDlSuCkKwi8
d9xGWxBoXAxe9RFeK9XuDxAA8kvzukETU0kaZ5+wJFQ7MGjeiIJXhzn3GA1gg04i
BHM299lQfgSwS9789Z7C9CYQZr8uApExAxmjPe5ipU1P+lP1v0zt/yWrrX/j0+pp
TtNUQTI3W9wnichW4oBNvEwS6xy4bpizeUi0pWCqOxItEzH6ubtnr4n5Vg8Z1Pkf
E1Qz629POVnIIntIlVW4uL5mVnv0VaOmp7qpsJa8NrAOaVkon56+M274qCZPf7pb
8DwDOJ1DPuA6hA8OjDbQJK3ro4sbQV9ny8JOGB0ntXmI7lKeRJcx4FoXxuDxfmCL
ZlUASyps4hP8in2X2RfjRu5YdD0UTQ3U+Dp94FK8Byo+nkdRMCHdJH2y1TPelaGA
8RYnEPxwggOo7FfHxJcFua54FrnJ7qAyziGB86ZW6+ZVvjayi0FrD01/usovw7K4
40siCFViIFYms6FgCyVsEXiRwCTVkNk3DwsqUf6wyP5c3QygVH6J3oQj1V7ear7O
sE805sYD+EVMcQgiFpNMgbs/1TodiiXJTbWT+ZLhKUpXO61cVqcew0PmA4XcD68b
XIUfPuYt+GHGKoA/uZmgsP/6zYnIMutIJDpm2XBXj7x2/7933+cH/ztd50at1nLE
OfPVWzZF7VNzEnUe30k/rnb+9W0b168jopEKs/gj7IVCny+g8CQDVQawDgfldoqH
gTU5PEwir2fqBGvKzqMuAavfF9itWsr2BJ8iU+tGLIl1C8YgfHcC0siBt8MJmBDH
OqTmWZ/s0TBm+TXOkJQXq5pYt7H9tFXuqinzmN3IJnWyQngJUXeMgHyQthSxjY4k
jH9dMhZASrf5XG1IgKgytw4e7T3aZSGNu8lx4qdzVzzQLX6wLad2JWwj8vxgvIVU
Qu4KGMhLh0qXRDV5vwFGN1HzadYjLsrXIPvmstQCmD+/zbFuDPK/AAsAV+wYZgCw
+lp6vQM7WAkFCbtw6hUAAiB533Bn7kEANA/drgVzY5undRiVoLCOF04gpxQXbkLi
836TR65KoDoqRtxCkV27AuW13xrDQTUWs6TOglQ9tjbDglClqqy+u8JRj8ZYCMKS
yPsAbMgt70ka3n92tGcQJeCZvPUYMHizkP5jZvYa7b1mArYqp00cRH2K4pE3fc0C
ssZOqcg3FJ32bjdlqCT5KDoxtuELhGXZDu/gz4SFAV+YcWKwqS1F8IZaj8sI05j/
ywWi73yHL7ehaXyLmwoCHW0d2Kd/O/QE1OJWk5J+rlM8KIyZvtBMaC2E1IjWLJ01
5jS/tADDKj1GDtt5FWiFplAcR8MJT7yGIpGFuYO+9d0qx4YVZweyBA1mYbYtJ3HH
9dshQyv+BQ6sdNUhT/ywwXEW2wTsk309gjiNgBS6Pek8zMyoHxj7sTRz/bNr4v63
HLMg/rvyvjH+tUl+hsL/Jf00XEpagGlgIJHU6vxQ7l477atGMUkEp9KrBimqtQIM
Ekl2zkInGGa20Xd5GMEuGlSyukJirn6Xn6tvA2YvH4FuXh/HyWxCI2Yn9QinqSGl
jVi/uB6vCRhdCpXkZWDmAYeAreRKiOYgDuzcPRwmlxJmpvqf1ry7MK7/sCHhH63l
DLy1ulYcknBNVq6vnGAlAlMasOQ5QQd1i8v0kAIsLkMF6/jWDd+Hqb7Y0h6NGs2A
Jdd+I93aR8B/l0/iskdkuHVXz00cUEcPofsKvnVY/hZ13zBb3ZAB7u+T2y8dtaDI
4jj1iUyIyryjxSW0cSTwDDPegIdoJ/X/K4dvr2SGDyeyb8IlqvcYb1Fo/oHVuNDS
rzt3yvjeI99RyQZ9rqnx7eiQfdkBRtLjvamAvArNgyD+0sIcE9L7P8oNgoP1F7QJ
W/1EG6FtYS51KutPIP6jGQ8kZcxhrG+RFcyibSUo5touvHgy8QiEPjMOoRP7vi0B
MYmpNzvRsI06WLWwYdCRNyz5PIcve/mPXg2RntaiHPR6bCrKbrd7R4jfIbJuCMFC
Cc67SH2wxKeo8rOn03nmW/3OlLTx6JKuJViHIWHo05LI2YbAvh4OxznjJiJPz3r3
YNg3SxeFdPraUOYLymCFJw15uDU67VcE05FxVzo6OvHMK7YtyuxelkIOCUgcJ+Xq
MZawq58EYblDaH7ZfU2jE7Dol9tnJv4YSs27dXnVEJCcTZ/8hTbYLRgnZih7zru/
RqjxgZhbPcBbYZXRBdqzBjrClKmetgYLLIy/XW5k0EsAajmYqw4bTUwJOflnzPaF
ZyEEJIfD88g90ouSJ23/3YSAnvM9lc1ePoKuzcFCAX9Wmiq1VJl3K7a6fP0bvlKI
SzAwumqEJuCas3QpV4TyfyZ+0J5nsES5L7pT23/sZhHCcrU886zjmqYLvE+Qnido
lSsnojFyOtRHGR0OtXBZuXH/zcrxbMj5fhWlzjyYJ9w9o5Yr7F98YRUlfTmdYzEL
poFv1P1zW6S8Nfcag+3DOZmexmSNBl+f/trjKyp81LkSU6eG/nJmnPMmPVAXnHBs
7je73P+HP4kRLDESeqHRPSIfqyojgQlUKWWajpErYvUS0w+tVo4otl9vsrdhw78l
wqR0q8fLDriZ4woF76bvN1jxb45qP5UzqMqYxEuuPgMBHdgiWNHbAbFYdngcoMcm
RD1uq/3SL7CAApFnpILOCFSiYnsYuQ/ERrD30LE2eehrH7HNXloe0wQRqwTVDX6p
XusB76CB67KQpm1PSL3gu2C+UG8QRPTtswriWm0arvD7kjn9MtL9sjaYsYaJBWno
XdlJyi1RwkI4OoxaXRbzs0DStVI7JuWVLMoI4H4uITWIAK2Sb357RI677Tg/3dT7
Rx2XVtXkdklTpQzG3dvzdwgObfm42T7Gg4pkbQ6g9RimXwtgXKlmtDVomcWcIweF
BbCfL+dCkaEeQcCVfM5RerS4A1hUcftojPWVf6YIigWXZJ3nJs2Rg6TLtXp9B2mc
2myReqOJP/jKHW+/Ss5nT3KyowhD5LO/kam0gm1QqRAlLwaXEsRp1Hmx1LEf9n+4
XByFcWnROxz/F64q02UnYH8uHon7HFL1lHo8INFKivku6G2/uvGc3IZsgh+vHNfa
3tPFXJ0oadf9QhRhxY/ZMwasY1Q59UzNNRVcQ2YcxUVBPA9Akq8drtVW1SBNmCNH
X1Qa3WFSsFgRuawr168rE9NzfB78RbmZDwx8jD6YdaXdniQrwTX12PNfW20C0Fba
DVBQT04Ud5Yq5peK1hoc+SnJjCkqyHljP7zEYqZGakyoRyzLa6SIyfSS7QNSV9cc
7BgJwJdDyXEOypy2PrwFnVYwdvvvOKwNCPF5TCBQJEfJ/5WrgHewO6FNWtuw99Hb
/JamSonsExwMvhm4U7GX05tJHGYKGPNmbsEp1vI1CjSVMGoRLCWeau+zX7P/O/22
DPTNPssLfeRvtPLdAYf4vZn0V4wvycGBX8rONeUaIohXqCMoQTnRdjFrTGRY3HyP
+jd9bi6dTrwuHi83ZIwjgG8wVpS2yaYSZIZzwHWANJeTYHogpVUmX9GQH4dWv9fN
P8+t/g8Gbc9a6wRSQJp0zRgXxJShlmJLMQbApTaal/JQaW8cghLuB/tm6PCs8AIE
mEKYlTz2JEhMv3hcg/Gz9I3qPEMXbf4p1hVbe55Ipl8+L1q7phKHo3uxBixGXRdu
NhcbEkToNq0zzq2Hv+NPdUDzRti0S7Bg9KIGQecnsN4fniN16obR6XIyYdwCvT+m
RcdOUeY9NEvTx/Rh7LLARFWUekIkI4540lU2HOd8+gU0SH6Q5ofpTFd2A0yGMNxr
VpgJTjfLuFvWNk/04LCurem34r3DFvERjJQwoYt6c/G1sDgJOLZOS6DGZJBKlrt1
u82DDbqIJRK3uM6T2kaVhf79OjsHqS+ZbcCqy++XBBTo9bp846nS/SRxRqhTNY+4
4nLFDYs0hpjiWAe3JsjP2eIBlH02234o+PymrEHcUH4mCI69JXaxPYX8/7oW3tF/
9BEmN0HToixiCDRkZO0/pdKXxPSaCXaC3Y5gwnqiYDCvHKywxJYkSOHM5r5U1WGU
BYX17nTxzQAoLCXSNjSwCIxQmopdbEFUzesOV6sIpXn1SeOMSS2F1k9/wn8JH3ED
9L9X+SuxDve6xbCmlMTWB4MCfkxzm58LPNk0WPs80GV6fS79d6Hb3HLjZO/wVWfw
Vm4FuGpwaq+axg8pBZwN6wyuoZRmAGZo0jA/Q3lXWin2Fkia79xka47yY6cdN8x0
98Pzvw1LNg1+1yfEKsoA5LDeiYeTwo6GGDvfYXH7CYFRQbIzY+CSP4CF4g07OGFR
gOTRUbAsa6kA/4O+/emosO0w84agmPf0EnJPj2CrrUW8WQEdp9pBSEj8MGXjdGpr
cELBUDJunNfdZ5jjZqTFlUTj1USk/+/A27qP1+m/tKqDhyWt1Qw/yXCL1VA14p9D
fGGoHYRxFYUSiol/UD0J2lGoUAC+NQcuZKHnTmJnVpiU8/3kbW84lVWYPpEAMYNY
kl7BqyrQv6pzqeMCke5GkmM1y12ucpv7NvrAWFExt0uBzWbl87TTyCcf/hN7WJvX
mj5Du2qn/Fv2yJLZKq3iMEmOkiWzH53al1Gzc2J4T+kuhNGN0RsOBuGEWjwtX+2c
TCV4PZfs3SiloNPubgCLlMwMT3H75plH2UzcZisasyzQxi6wNpklhJpaMeY4j0qf
pusz9Yxz/OXA549Y8056zExtNY92vkXoejBrqlKkpQDmyQzmxvREyo6PoFiwNYPP
ljokNtjeQuAfzcttXV/+qDvj5VALS7PJeqFXDW5ugjslYdN10V546EeFNW/IIs/j
LGAi9Ls9zn/VV72umpivpxBlm5kS9bMI0igaVZ3ZEgtMP/AXTRBE7e7mdjAMJT04
vzUZhwjPt5wYFw2PkFMBz2T9IsfgOjCtybNSVqEiq40Rq3EJf1i8d6jzeRChjlKT
UUtYAhz8cUrsEhtY584aiUkMX2een/piIhn2GPfGS/QRzWO7/i7/SYsc5d4LI3jP
tjAnk8Wlz6h9jfm2esSVAu3IHy+lGpq4Q2lpJbMiO3pyMapkkAcme+GMyoeA7b95
wIPCGjU1NJsMbFLtNsHrbEYAgAQ52ESy+fKgoLAoknYrMWdeQROrQu1vMHlNKFuN
f1cwHpIfysO/86CpYRygCH1ReqL2nxMdcqwdFCq/cMb5z2Eb12BWmf33DmVSy/ER
aLi2PeONYMq4E/jwe5Jdl1cpav7Z2S6fH0pfxEi2yiFQoN2y1kXhuDkxFLMsh6C/
LsJ/ib3ZPqPLQNnOiLGBI2RrPjiJmSB+uF5uAcEIat6Cd0sDIYHf9rUI9/wEcg+Z
uVg982/X0PsjBN2UkgmoG7ME54nz9T/Mra8e3ld204DE4BQ6yqMCItYervT17Oos
xgFJnI9zSfpMW+FqVj7AEfNcAClhgaiXNwDZHzyZB+Vdx3xNOfm7VyLFIJJidSe7
RqbYxdQ7UjgnxGrKpBfweBtYbprMb8JmmUmCINOccb50efN24bANvG+VPgCr/OFs
189JE1k/xRvYoz2T4uAHXQ/xAUDxS0t1xQ6pMmS+OQnoMg/XeU2gxZwOKPe+uTAb
dzLfLw8n22kUtcAP0uw98osXNfYNR3jDtolkew3CDJHu8bru8dVkO92HoLkc0N3f
YTSrmaagtavq1Swz2tsHisnLqFLqn85eTmPdOXcjdOulFsUP4AVXKrkc6JrAg3hJ
Q7MWyClOEWmZ91rRSMYe2QpQClmMveKD7dFvgPNH1xROUHnuJrFtEDY91Hs5VXbF
ciDt1WgNslPZQkowwb2cJmWNBe9/8a2l/1KChxc69EITe5ZFG8JmQb1faBiZdVD4
qkzj5gAQd6Yfl64D17TRPSVIJ8plcFlrs9KEsq7QwuC9FD8ej0JX8i3XqOSACA6F
l1H3RgqG4USFYOLnCX73gQ/kap/LK4QzQD3PHBtnxtMAiiHLUdTqqAtCS66mRHAa
HWl3IJhB1ijNAUznzxbYqUmOEVOX2kxXZnbNj2B2gTTE3POXwWgmtiIotckJe3WD
NP20TxRa6R/GPVm58WQr2wonPU8+hGOo5LHSl5dxnM3v6r3vv8dEyoenSHjd8kRn
vFvU2IfDW4dyOBCP1DxbMZiR/zcbXZWzLbcCEPrFM23uCrAVRpv0eLoSa1SuwA8n
xjGvFNlLGmZ8pOUbA7lY2GyJ/cYXt2TtS9Z9vDU/dBYGFc67IIc0wnvmRfTGejJJ
GPmRlHdptPllgKsCHF30zZ8L2QAjvrbIhmLjM0nXnCs6j7qGrejib67Xjsw9vWqj
tPb97UBvvTE0jzzlFA4bBs3oDhbZT6AdqZie8Bu6pFQreboPKrKLS7n7xBA0CGlg
dJtBV9kJhYUDq07ER6173r5GLMk3H0bLycjKWLQRPya1fOYVqCcSUJ3/GCLLDrbS
D4B48hqoB+6SBq1Bwk7/Z1IkQh0Lt5zQsayRxz6Q0LM1GR9N+DKrpdAr3OFJJNS/
fPkLD+FsOJ673BShfmpLyNfbf6/vxsd/6z0dMxkOr7RCJyAPonM2LbmyOqTeKYTc
aYsgDNdAgLR4r9N0kB8cGzO7QS1Aod6evuG0ro/4Gbcrv905N76qvcyQOT5dJxw3
y+mQimzhyTp6CelEzrs7Wn9vYEzV7ZPCTnOU794DiSARroDLFUBusfRcsNe8FWoS
0PKC0T9WV2ASwRAKmH/SBckeuGf1v9p6dTBhY5qCD1k3nM852FnWm8I5RrIycp1s
3qpDVyNz5tmoHeimDKgm3TG/aAR29loY8cTPGYVGPqpBo3e2Eseb84FkGLSWjK08
xuDMJwel+nmIQrFFzbhtT0xUcjNp/mLBuTlSUiMrWMIl9NhctMFBClgDnM6nN/Dc
9WMG6Ih1O7KBMQXU9/UOUeSdfS72YidtM98V+PZ1JM4FK9/x1PFpF/imIFsxvRie
u0knMBPQUfwXEg2TNWUTP8i3RD/GFpKEY4ruwUOS0dVxbfuGz6eWabDrdhI+GoF9
BSQYMSvTJrORsubSBod7jjiJ3IuhlZyVwYa1F1WTObH+TN3oSv7ln3Mzv/SNK2Xs
EpQ+z5DixvnPpAgUpeWA8yFCOzkigMexBVzeNQGh29ZnpxaeF3uaOFQGtS2StofP
GZ9AoOyBfes68jcD9cbjZgm5eq/VVLZ0y8hRNgE4aZjICLNrk0L5uKeXr9REatQF
z0FqD9EHL4RaR6zZgEecjVc+kMuI7qpF85pkv+JDl2NNMUPmsqL2lNpP4kiSzrY5
vZcYefZhggGkS5KC9g1OSdI2zjqQIp9MST+9YiE1H3TcF1nipi/OrPDnE7lz/cWT
HGPlnqAiG31Cxk+HDZGX3gdbS6VNktcNC3yKtKrTpkVeGYM0gVmCTcdBefhA+ef6
9Xt6TC4YimnQrSezF5NXcGcI3GlS5QOws6y+90/89E+rTNz6KeAX8Wn5A8E5Lxv3
nloJvQGgy2jUzHeWBl3ogtAp4h8DNcrwJAj/R1fomeybL8ksuVoC6qtWIR4bUgZ2
yVWzQ39g5eETFca0IX6Qgb+YXYYREYRxoFAH0du8xU+i36tuHmaZgAjvjAhSYeez
/XnuXmTY0gmUeMgDx43n6mDBJMQmoI/EmvkstIh55CQUegbmZ8KIOGNPeX+Ltwo+
R9knRr/BlAphlxVdVsYA/Lxv5xiFxyvTHjvGqF0s0Jk5QBe3Tg1w01Y6Y355gTwj
ewvd6wkZU0hCpY0uCqcZNaRzUZ6XtGgoRkyZL+dua5jTaA8j68ThfcPGAQCw+cfj
PWYpzExqWrfkVJbwFrsEkSxvB63rLd0pXtUV0iVBOTTbT0icjGu8Byl4BBDW9fUZ
gdi3duNACE8ZijbKMf76P31cs9goTr8MNWfxk6XZzFXqXBrRrP9glIqI4Gu8d5g0
oOwY4oXvMsMAWCY+4ZHw7Kh587vYiZdKtxFFbyxjwLEbqxN5JgmU5vDbyAK7zXhX
8ECqZiWByJTbo4/e+blN3oaP5ptx49vllHR4kftsUN9JeouTFb4DbS+ewd7C/b/J
p2Rb1vqowmt0+h5jZXh6a0TF93cdgCQDKcqDTNRU5UE0XyFaF5Xu/DAMFEloLQFh
wPwswxt4J4UxgBALWeUYMX7MQ4xAFZy9sSrWH9pgETR4Tb81cqMNSMnsObBVMsZw
UtpwOzm66e6apQB6JrVmpA18B3Osr8YWGIrYDG3rOUAhPMa9JuuMJ0t+WupoXPyB
JLwWLvzllEmTC8hyE2P7C2l3jMrL/huhsUoO30f6N1hW0B5shML/GxFIV3M+uUiR
UMYM/DSwcowKDzpsYRYh6xDBo7Awvw3jAtoHHulGOTARs4jg4VQ/LasqGnD2IeM6
cWTIfUPxpdNBTA2itfKXbTZ387BAse2DVwOx9aj6mxjZZqXEMcdcxFqsQact3Mu/
UdzbF/tXtbY3R6MYNGCmh6ohnxoxrYtJKXwBZuXCEcLJc3xRZi0DnK15IRzXvBVr
USJFVuT6pMG5tG640/rfc+TlhqohpOISdcUzGbWKJZpW/bqeg6MRuSCQPDMtwube
ExtncOA2H8Db6vZ4XRrG5f3ZjV5sO59NyVehyKjo1xBZQPQgOmCUQRsB3322K9B+
vEkCpI1lM+Y4DoJ256vLSjNu+snIeVJt1qA6+Jbu9G4JVSPkps3xooEKXqsXe599
qglq+p2nixbKPSYKiTYAxMYgU7NGA/GutA+zzyGG0WyWirQ+i+D/sPqkr/OD9SYc
rU9Ljj2URW0tuAvh3gjVDA2nHwMhf2bYF07zIlGmTcLjoQb7nztDbWh+0bGnx0Na
IdfbOKHyKxBmO3HMVdJcFgvi/3QoPufDngurzLxAD415c/+1Qq/r1k3tz2zTXr7Z
PqxKwELmR97UXz3SyKKdJOzenGgVJgMYfghqd+uzEMI2DU1f4V9coziBUVWAr+UZ
S8KCgVEVvUadJt+jri/2nlgClmeYupPy0a3YLZdmpzycY7jSeMV1dcWZdAXu4X0B
xuSaqZK2WGRfU0+N5lpEG+znxPjHLbryYnjcFwVHnvurwK5LTYMOOGYZUb/mPJWJ
XpTv+He+y/3BLbOLruStPVsq1JLk5NJcKWAOs5khVEpayooxE09BXr7maKmMBptt
hJW1B/46CFBRpr3T3a8ZlyavxhxE2G9HkdvtFIXApfq/lt/huSmSGw19bgPsWzyo
TXlKLvkz6iXY9a0FXKKYqtvJAZvoUpXFeIwSYsPhjew7nb5nBSUCw0aCNoeTXhUJ
CgRtQrvQfWYBHdUKigIbkdl1Oqzv7P2jvFLZIMAqzB38OGCzp6sF2EZ1Tq+exV7u
BRudp7BWZDXsqrzXrUo7y7IzyhgDZtucXHgp0fziOLYlJBfZ/bCEu8ICqtMbqlUN
Bjpo/YVV4o6N8sDDF2k7T30mz1wcuUE6JZANQxNti7ZYXQDKawWXivFxvoDbL9yC
ZUoelbpG9foaABDaPLjLPAjgZZRO1DPst+hqsU44/B3v+k55EEioCsyIUBzGBjaj
D+ghkd6SCTxQD0g5+mlflmkINMCiJBrdlZgvbhSNGvfRJ39JD8sbpcWLiC7rXvbg
t6chansL3N6lOPnPbFjEaiVJxGgp7iT5U0saBebLY3JPQLqQR+9IygcsYh7JYi6R
odJOyc22bf6DkMPUaNk6CC5yz9QkELCvDVLbr6SUbP/ljQmFbc+GzLC0FgqtyP2M
2T06byTJclc5l/t6RXbXpiwRXWw43ylawbEkSvl+ilj/zOVAkXssCjwYkP+0LBPA
0jW3eR9wkThpFUouX00x8dS46GdUeFHXOKp0H8Y+c2emmx1NkBKpyi7hkKgiOEfv
f40XwiYXyeJOzF8+M9NTSdQz23EBvJnlipTvsti1Zb/88GLGc3Uiv9moMB2s1XoP
bIRa4VLToSFkNYBlT9oQKsb1CQcfwFEbNMqI37Qng7mySmBvvmuz40VbSaFKCkMY
uWcnZlbBKawcQubs1gKBvB6D+pkFdUQNj2TT9YCT0Uu/DSTUNRW13buS7KX/0zyh
Of97hkQab6JA3b2MBk6GycCvBYyK2jfv5N+HoDw/NgtvX9NDbqfKEPEEvSMLvQsn
xtdBHqOBg0AWOK7T2SJaRDqYcC3Rsxa4qb8vbWte5GNiVXKeNq9SoNFAb3ypdXgH
1BTLk87z2yLvjsmtMGu88kPMAQx48zBR6sQAZrm6z9lETC3sEcyL/tsG9wgW2Ntr
588COZv9+UbWcj17lzsCKhsHbWXgoVPZXqVL5jiHxlCPirSqpRONjpK3KrK/mKsN
KkObXBrkw3p6EoGsDWs6YNhT1++PVk66WV/2dkLlIxjIRgu3tVOHURQ6HK1p5X48
gpl/6CPKAxq3vIQf2Hunw7d049vL8uqcCkmbcNlI8a+K1JGRGhWMkhdla9qkOf8h
xdrg2OmICdI/xNn/i/54cNWAmLT2hjslqxBK9OUEj3SFfwwqQkyZokFBdMN3QMTj
Tai14BA0FuQnMaVAI07WbIS28sFqzgSLEvmuEuRcYjThoqxnhlJmdOshrz25DnWj
jASQeO5wl2x0KFAUsK+6BzDt1/Z9ct+xX0pSBVPVnjdrFWSGEsEcsk16s28pjN/U
QwPICzXpyaNIhvYh3kTDj59gu7jYB6Dkcq9lYUihadP93EzytWZRTnh3Yfeeqpln
jd1F2I3BgBImSqDvKmwr6Bi4Dwr3IDDlNOoxKWvEJkPQfCyBGdlxIzSUAGxkGeUP
eYBEIpJH6egsPF2dBAkW/sSXOsvG/jFQOD11PwjSM1QUOBp5cnbelkGIreH/SjHb
6I3A/T0RQxa9EjBgMeGgWlKvetN8e1fCvRnMBjA5g1bJSxHEy6tKpDEtzwiCVLBe
egbtF//BkAYuokW8GLXWOntjjVfbwD8SzcS7euDU3lXl4p7KUWtIaeVprLgGovAI
73WPoxoWjNpXvkZlo8HYt4KMlhe7cPJOT+IZYWSVYYxo8hO4z5YBxUGgGbAzu/nL
WMibqdI8T8lyTcH3Ngx0iP7hiZ9Ik3u19irA36fxEq6DJCp7y0hzYm9YQxbDCH9N
GXwtME57IrkJ1rHsLEA+TCSTMaU9yLrlqLFBmV/jBwfuYWTkmpAavZluj8hq97Ao
V1c69//RZp7FWHaQgezVFCZDaPFNaqjPUUbtuoRgyuTbYcP3sn7GYAn4BufMEk/a
2IElr64KUZ0MlW6UXouQCsfQ6RqZyE5Eo+6TZMEy9dCXKo9tJGQSLv5tia6Zgy6o
qjeiOAXTmKOgKBOUyfMUGlhJsTriXJmYdUvUYaT3Wxd2JCeDN0vkPsiso+nSdH8x
mJ7cC6mju067ENT79rG44CtVzEFrtPJ8YdI4x0puLuPJIts6mVAcYQ6Jz0G7YrgS
uX0wa3sFY/gT8TKv4ew1EOoQ2rjOTbiSh4Ucmma2V95BUTrXTEbK1nReLVcGfKib
Pg9/64qxwcOIbrLU5fvNfUgC/jjd1p/QAkY0ETWbPuWrkGmzRDt/6CVkjgT8qNad
Iu9V9WBhOst0iUcd0Jbf/a//4chQzHBQsg18f2IzYQTJZNeHrLqPzdDlzIc+/JVk
ZaYFbw6e9pdn8dY7A/70vOAMiKB946sQZOOepGQXX0MOZfEp4+jUrQBKPSzbkr0W
aDHDsMOfFVT8BfGq1yZziKSr/SDKyE9H8nF9fUz5BVRkH9p0pms0R/q6d6e8UACg
TtsRRMDURi9kv6A9zSVyEuoVSHqX3U+FB98bBm1PUyYePa2mdg+dNoW85LscUQye
YFy8TF3zoEmSPWxR+DFhrK6r1vdj7MZ+2uxpL96LAlnxxaEJsbM7dI6B9ytJXDtl
cz4eJyTufiU53aUACmT/ujwgyzKd2oHL/Kt3iecx7p7xPr5mWb6qwBrBwE/0rJuj
SvBqpdZ9ZWjc5PpXVSL+m18pxwrAHZro4EilRtd9JbnGwBupz83jVNOsLZzd1g+l
jPP0fcYJ63cBHlnYXVMez2EPiHDGUpz66sEi9TbarX46hgA4f4esaS3RxtNxSE8v
n3y8RCAFcTlL0LfVhUztaw8Wlu0C0gMDAMkjb6bZWIvOI+D1pZhXuB7ImIkXnCmi
AQlZjtB+EeLBfQWghJmTQM1ByDDGZSqL8a2HEQNjyIb9IYpHB+D/zRUFTzNtcRvH
HENCUTZE9BG5wiy/e8Yj7aEJ8ysJIKNn3wagXYrrHaVkVhfnwqiw0MclGdkBUqZ6
xEEYvboIPri8maxtAlgbxvNFosgxlRTks6O7mKi353KMHLvd62VJaFQFz9B6oNr6
SDaBBlCqprc306GeyXN3znewbF+2HtK72Q/mQEwnkLUMG9VrdQhcC6uOwxKs+r9y
8mN1QUKRrqwRWRYaDCci3eQA18eF2XuaZgkAk/Oqbg3oae01oTVbAS4xAcQxz1z1
W56z+OZPknp1U9K52iqZH1jQVh8e44AkadYai9qteKL82LcT2b3/HNaAbEbuHlDU
J5j8DNSJEAo+PHtAPxnfkK6CXW1NRvFgsf4XMocEeX33o3HgVlS9WIW+oCn7OpGM
+u5sfi+jduUGyAHpv5fqUwtWEyQ6Qu+Wf1rnZJRns45JOp27TzbI+uikdmrBSoS2
trWgWzntWDvCkJFtsM44gnbCR+O53vgdAsJCOo0PbvMUNrUOVYwz6RXLpknlJ2As
FZ1g6B31KI09zQBDY3TLF94sWXgrXB+kk39D/q+47Y14Shu9rbB7neIzdpN5Xxyd
lTWvIXnmnaP+RmXhAqM5Iwc1zQVjn9wdeKKWVhLqGED19rf4Sa0dMYcpI74Q6xxr
k06TP2WatHsk0lgTl/z4nhpyT71gMAKNh+Tq0KXyg4f5ruZpgKJNJr/qt2goYQPF
SJlO0492RhrxAZ+f2gLni+ZtSYL6hee8Lvm9ewB1my451LPb8H2hlWuSEB4vtj3Q
CnNx03L5kajO5+3CM3UwgR33HhPKbM0aY2knDpDribcP5h3HrwmwpmIFAUd7alKP
boCcGCQ5Ed5SwI3oelNPpkwN8jogpsYBElXf9/pOvSdPJ4xJl95nQ9ofSy25HxRF
50OdWDIvE6MTzvOD2Cjqwlwh9gRQz/w2009luibum2F824/Q9TxEZUQuuHPqt0tg
CBG0ReupIr854RGMTlI9C2OrBR8JqRzbxg7SfgC3TtmmBrUdeD0N9taaHGmzDkYn
wAcpxNdV9omQemVDjcWHulVHhBU1tOrHRqNEGkJY+ovXwn2SQozl0sm2iL35VKOC
Zc8b/05NNj4cfg/0vqh6pttElBZKSrgAf71NXNHydtp5vGrvq5fsAeTVEyKd2VkC
O7WelIDNoxUuTO1JoOQ+yHqWvZgPpAwYy1NhiV9IqY+HPP15DNuhTIfeiMOv7Gxy
HAvWm3+Ge77m3GGTxCdyYoxOa2zh9qoqIKbS9LV+WGROr9+DJIcXhTi8G7khlrmy
iIc8nL2nlcPVq3imGGrrJYXQ5uRVuuSyIoTzINzLhi20E7VsspTWc4usllbCoJhw
ENE3H545amBC2n+Li176tNzukQoif9mRGVAjRNGy/qK3joCIPf2XrR2YSWIczHOU
4UNTbmYwRVjXsKYtvYz5cXz03X9KusjXCl+RrCAgHzKiBHK0+VeSkG23IYJxUE+7
HZdJFcpsmijf/BQEJ6uuWKcaptkSEwGscFXXZVri8GPr+KSy9P8LXEq6NN+UdMTu
LfBqLLO2JjsWy2uzoIFUmIDDiP6mwq8e1o8TWWif0410gDmj4S9TJx+9YtGJemZJ
AOQUt0Kc4wUvbBK5d5OxAD/FFs7ebDSsh7M1ixBL3r5RFw/nzRipGgDmUsuXdMY0
xp+3ARDXmtOMs366ZTDuPqKE5lVF/mcN9v/ckxJ+Roo4rgmmK6bgVG+YVQgh6EAM
KKHKHR/RIUMqshk0ikwdqKlj0NryynpStgfvgJaP1yVNgr8hPAYstiClZq8L9LkQ
GJBUVW79j3ApwnjUXO3+S8Sg0/YLkadwL4sEkNKCqJQgh5FI509tM7YU6rQX/FIA
SCyjKycLcSivdRizsi0sHguIFfojr57Q3rmanEtx8D94FGNw7EwdBhjDqRNOwiAE
dyY8m4j5creu+A+Y1dmfqJ4xwZORWsnm87uE+kSWbfQznqZWKVZuqrY7XZk5D5m5
S62Y2fcmAnSS8an4aWdoKV5uuVf9Gj9BPSp6pkr0C2ZQ/pWnwKxAoUaA0AlWcKsD
7t5fUARJ9/sa6PpAwsHm5SPX8C9+30+uvVS3gi0ZsbMlG6ky+mkqxKDSBQxxZDRy
cAmHKJAzjehDprcN4wbejHRjnQvuaaKSRa1MioZoXsdjydo8+fJGPi6FHtBMhtmd
jPQDrnOIA6GXJiquevaL+GajcQi9gTySG6GpvTEBm5J0dsBqBkN5YuvTCcyWOLs+
XLcEv2GCpydvPlJ6P97+ej+vAr+rA93iGgmk8Uzk5q1J+cR3513ioTTM4ZhcAz2T
iI7Mmzqvu7BrzVdPllgjz6OEXE3V0/BlKcFDSGSLFx2MfflaGd7Ui7RS2FurmzuV
cS2Z6a/KfzW46IucV2UDgQzcYgEwxdrjBZRdUN3bGiHvuDHfqRqE+9vukw+rlDPx
/GcOYcvfrIqpe8ZyqsSUJMIy745wyau+2lyt4ruT9VeGkqzBZrK7fNzXQS/w9lCG
BNXVUFKBXdoIjiRmNbXfaOt9FbB+fxLLJjsJQq8wQtgHTMPw33vNz1HDmlQtXo7d
rbKkVo31U+J8uDFAjhmJ/aghLlVWyn+FwVKxyYBxX+PHCaXMArFBfZJMNCafZz8l
oUiZhWOBpagyMBjg2EJsMS9hHJQ5u+nlpvJFHL4gY8KN1PePM3eLIOn+O+jLDeQn
DMcx1mYadeQEcV6+4+lIgexOh9+u/VbWRA2U263y3jO8C8hd60lj+eF318Hv0yj4
MTFnNIanbDQgP+vVB+O4XD3k7WHOJrSf2ZTH8sjc1F4WFDcbueT8/OQR/m1n1Wid
If/9foKCS3OXB6ZQGQPW9CYjJj3A5/8ljULBQqXtotkT1jn16yES6tSKtdF/zU42
YmZfLi3BaVqV1+NT1lhCY845FtoT26T81o4C6KOOa8aexFnvRZQM/52N4K1f9oD1
2g6Hq3nl0vmAHhOadwWZU9b78R/XiBr8r4yt5TscB4AIppYC2dhBYt4v+yikHd4R
jRE3HDepw0uUkb1BjTOUWhS3ojAD65f0Nzk4+yWwfCh9pVdDx9JCiEGZjzJdED1X
CgdFtZBUklMeWMsgRBbuT4xWRTFaaReiYfCXRbUnJpSVy9RG5JOOxyDNfPbErIFk
h5ugW8uHV2uySh4yRPn+e4lMjKWHGF7cuvIX1e2RPG3nAawERNY9oQteYDPTKsCR
06Ii7zEZdQDJgLDjx4tSFCaq4toCZVPyn/yaEnVVQEdkbeMKKS6jal4LluURSwnH
Amomu2y7oaBvnGA5ZQTHk5/hVK66whPoKAHrxjlt90d7t4CCvyebWYvhByshRYds
zKInagoPl+/hbYQmzFnAe2wnxDZ9gVFD89GHsrmoHlyvKLAWe0a2sjbQ6IQXpyGJ
oSrmx10vZz2xoo8qeTYMMvNzwPTOaWz0ms5tnSXJr5Z++yW7DJVug/KoC4kV5bJQ
75F2opzy61apMA6JQmeuFmYD9OufCkbQAGGAySEQX2tl9vGE9TXaFp2qmBMTEtl8
hWLWZsldZFjZbrO9drqV9eVFDg//EZfgtoo6ygktDTfUKQAPId+XWx/UXh2zlTCn
akfA8C/bRH65+9FqA9KXd2du1lUTU5IbXKBYQCF8ZFs/Kb9OHOwnv9COHWuQ+lYA
dw+asjHR5iF5H6WqP1juKze23CDAOC9pejAWp+ZY8s90fB8OUDRQFv8vbZsiBREY
bghF5YrdGAtW7uVgLGzFAdwdY+PJQ5jDBGvoiY+NsYxRQdkGXUGRFYlCW7rVRkO0
FWxUDVh071Bq0fFO/t6CnyvfvKSqlk04BtUsgDobAGhtVVu6d5jVa0evl2J2H1NH
6xYhChaaRcUlRoLK2wkgJNMfdr3XPMUHTfHWI0a13taiWbeY2BJyddhr4UzPqxBh
i+boZJYUfhg87C1b2tvy4APFlb707UCSHyF3jDxRazspC3M1IwkQQ3+udh/ExcuS
8jQ+X/dZt9EqEdlqlgCW9bnuElpWFGqKEi67HWDsDOnaBA5is7IEJyGwbQYzDzpS
PzERS/B9Kkd0dOh/eqcmpmA3k+1f/+AuC0FjX8T+Aw7GgWxiI+padQlRH+HqrGpb
J7YaylKcV8GXv6xQLhMMY1kETkYG5V/3ahFgBUkBBGWq82rueSnm+Km8kYaTgEu4
K7BE/7bbS+WBHKeJP3YHJLimzuJHYin7belf83noafF3uEEGWZw24f8Bzl39TQXF
ZZZPqk0Aa30n3dgq773pPIpZkaYj8x+nUfXGpb7KEjRaYas6BMlBe56fYqHt8+sD
hgVHF/G33GPBS2NbcKXqaZxiwyp+c6R0u33Ra8KHGPtlghyXMfx9JLsSoQtlPnbL
/3q5Skzp6oBVSM+S/Zd2AnZwEhhOd6qtpPkMkNGLRegt8YJVEYWtsAqRSr7SHj4N
vTaqtjRkKGet/JFwrMfKlQeI516INsGe6N3pGSV8L/7DxUqRjgoS7KTfs69/w119
TQ4L2A1PXWfVDbK4rr7Q2xBB36xgW3Rf/SrTrCYkRhBVdB8flyhcEYf1CL6BfViw
j1ioZCCT5eXcP29XsQJ6C34RKA1bG+fVa8VZs2MbXudZ9LJq+nB3E1ugXJYhrhDz
esakA8IT3HxxeHQP7shjQPBfaH6ueJl8XMEScARJ79d7nE6CLzbZd4YK/z/XEnLk
ZV4Ceb62NLMPcCuqvNqvJqlQ49YTSKtnywEuIrAUXFWncLs4WRY3O9I/3FSmy1ch
lmULHFP2Sk8Kko4k2JIKTAxwHKa3/pWbvr/1gAFXTMkaSn/8ulm1+Xm/U9qknAIO
Tp3Xd7RYuoglAiiAWhaWfZBxWCHHCQpQBmXCKsZwYaIPZtSmo9rgucIsx1aMr/Z2
U6wUhoDfikY3fSnAsYGpqt5fpApnTb4gDOOcFUVr6nUHxUG8wSgCGLXOaiv/BKpU
ogz38mTYDqXQvb/p5YtyiswRf8H6srgcIVZeJAgqFeltoCv6/K/eyCt2N5yCHVo9
INdldK4pRC90AaXSxXm7f/XwsWs7mqL5ncp36jtOe39PnqKHAJJ3sP+6UtNwY3tw
An7LoAmDQKU4+xFU6BefagDNchlLQZfX4p80LGeqvUARPbEWxzr4L6I52r/0UcDB
UUwLIH1zcLZHsdAatoONNDJ4ytl9otEw+6j2QrCy5BDBSrDY5xwaedQ8Y5cMrjiT
5qGxkkn2xh3gvHi0FsExZckK8u2h9kMIRORdWQ/LPQDNQAxnMKPkY7BoZleFZf1+
zTwmF4wUHjdDy5b7OO+X8CX7FYvR4gKMMPM240AvySByKwpDJo27RTxXvERilREl
3uYlGHune5TKCKHHyZZnWGhHMlpYp0QuQga6P3IU7MPDriRcQJP6HR4E6CXneeo2
Gpvelb76U9PHfTIyAagFR+RRSfz1Pp2Ri4vs6BSA8lMnHkSjxYVmh6/oPGcO3ilU
J9Pit7AEwYWa8CoDaDGQJrvfPcRa+9NwUOSRMVOS+eOG42Qt9EwYXC3qcAtoB1ax
QtoEon/SSJf4wnjxKLi9bOfuuLMzCHiTzIquOnBEcgp/dLvcmeh+rTV37na0JqcB
vbvPO11a9e9ihxHEra74U80QzvIVynN5p6zUbLR+6GlC9tA260c+gGR5cofGbRuo
MuRorn1TrzygR0GBIdCfuz7xedICjXN19WblqQYZuGF4zdNgPpSMhoosri2VYP3j
CXAEaEfeIdXqAlh+8M7ODTvx5Dtu4udiq8Y2kfFPca0Iw3OX9Q73OYbcq6Pnuv2/
6IeCwHKSOl2jqUfqO1FiiQ/yx7kIat8Ewd2LIdXDJaqjzYuzbgBh8CLloWqf/OTn
1ttrkWnh3I+f+0aVnojbBgctqzYceRlA69RKDpjH2U0Qsnf9R/dic1gJs1YJQadQ
0DZqIDkPEQo6TOG6Yr29wpad19bLyY5Z2cHQAHhVgafXycajfll0OA1Qqd4QKcrS
CXbUgioJ13BkZUG3UAXZODptBm9FHMM2tkBGDk2Ym1O15Hsn93V1N6WpEEU5ZDWB
6w4ksBke1NfRToEeD4P+r7LapRMrojqg2oIyrg+aUk4FPAXPc83tiU9PmzeJn6Od
qDbSijY5LC8Kx90ylA/oiMDNVzD09YAHICj3/uXORWxWfBAtWLk+6D6e5GCXZ2RT
llpZSaRg8Io0MkTpr8cc/2YFimqpSkpQNckYdd1cwWOaVciisAP/FxHe6yd8olzs
LHrCYtn6o/zfxuGnKba5+QClU2AUvdUJeR0FDouOZX89DGWbRCGtpf7XWtSwFaSt
coQr6UyO9ZqMlEAbCh4SxVcRw12eSOA/syKc4V+nOfr2SSrlmcQifKfYZaxeNOH0
mIydt0KAQ7cEUyXAvutk4U2oV+Ry1i8AhE1Xdrwk29jsf1C1ohXwdbl3iSmSIdC8
ZhD3anhJ5dmP2twT/PfbY2ROBU8htlY9GcamW+d/Oezw+35rd5U0VqyJ8xBKLxfN
IYavWx1knj37EXgPciifMmP3L2lnmUyu9zIaad86ENd3aXduoMwfzZ9ajuIncRIC
mxGGeWWWo3+0BHnI3TQW3LDt/GxNBM3xxqL5OhEKxmCg61BOvk96JzM7SrPWLKEW
H2R/8NMg9egkDsSPxRCRPXhuIeXBCdz/9HR0WxgoC9pBWWctbZtHcdZNc571Aits
r3fJk4d/5FGZGCFQQh9HpYld4m65sZs8qRqvhJi1BpT0sxdUrElIBxUkBWiMf5tx
H/KXA1Wf6pYKOjpuyPFMla35qgx2fbgWfiJrS0OR7nZbQMKlYUJgOPnguihwzdqG
ql+2RZbRvy0hSPicfSbW2ilJl/fIX/WWyV+aetvJrBe/9/tRgaZtbXmiBfPcbYnN
4/tZmOXAk+M029bzt9fBaTJeFEBIJ38ROVHb0pz5f9xLElY5GmZNpZmNdoFe/7Wd
YVJlyrXQ0gEkCKuzDJhnTSXXXA60USa4vySvTiXsbE5xZCP6gXCJaAJgI3buMFYz
vPDnwRNye9jEZJSc8MkAaEAu7hdBvFWz8nXo9VA4lGzmZSTsTLxpLnRC9BDMwab7
tV+wpPg6iCDM+l3AqAq+m3yXq9XfL6BZuGjt+suIuxBzuNtkCmbuaVdkn2XKxxfk
k6h0KklPL4u6M8sCUEGGQedZ0NkrLjaDgKvrargWIf5W/c7oEym3uD5afQGFHgUK
opbubz0LJaW9uAPYcbLatKYJbAUsPvMasmimjQlsUNDnCJrbQfinB1NrTfNk6bNq
CxMxYUfvJpPb1/mr/b4gIYp8izloeY+90q0ybZYy1T3LSNsJeat3F4gqkqXyEBvT
gJnkFKCXA4IkOyqBEpvBCjyXqWo8MNUx6jSLt0FQwH0/7FhUtHQ70i1z8pnG+h9E
093vZygeShdp5/faz2gmyPkRE+9xZ7HYtGPAu4pKN8u1s+5bwQA8RF3eTMmtlT1p
9VPV8KuWNEi5wBAx9OjwyLBGi8c6C4Wt0NzEQKrR7RaDPykZd+pre6XAGY6yiuno
13ciHGlWkSrcalUSWy4rOpN3ZiNbp+yZAY2XjZmoQp4fuM0fd9OJUVMUTHCWWvug
R4G/aeBzoxOlCyJxcnMkxwOes2juGHarHdmWylljcn5ZZHqqa3kgurJx/48ezlmv
pyusWuLFy5vIWU03aPsXD0qvahSsFUJT5VUk85XaNr3HxN/ipoL+vh4XcRvxRaF9
YWj6qzGmPAtifhrmX3GCEhFEolKtTq8AWsEWsI4mPKdlV2uI9eHYipwZ2b8xXPBb
XR59qeL7M3NjPj2gGkdSj2OOod0fNFxGlPPLLpV9rz/9ftTmL49DSqcLpLogq7ub
NENWzcCn9SBWwgrASlaXO3LdsMBA+qvinJ16dEsfiD8EQ7a3nqt/Ah2ZI3fyvOpd
RmZEGOS2TrMYKyCmUkC+kqfG179g90OPp6OZc8/0fRhMPpnIF9OFfQpD9vf8S4VJ
cp7kBbVpEuqDAilqIJolwKI/Epdu2ngkdcSoOB/3n6qHj2fnetsz0SAIOa3SPYKH
ILElO92ZMEtt+e1Kn9YlrGkw8AESVkwKnGUzCUwNx3H1yg15wTHJ7Bt+kk63kjby
NeGmuU4LdyuxyTRlckJlmYkxVrJqExaSMwIYU1/5m+sHDkC3H+mHJPcy0j1PxJs6
r76MnGvH95t3UfbnF5XoMjzu7h89Q+oE46g+cETw+qwCIvTiAY7raWm4RMSkB3aT
yeLWLIgKtU9HoRZwAYTNOF9/tHiA89Ag7xqNAVEeSQqrDJX/Vqz6A1WPrQ70E7Ut
KsCDQlwDi688kP5kAKHXQiNAr/GVB6Bjr04HP6KTWFJzSxcD59qs8mJdnhcOaqV/
0WDk+emP2WzDEoHizVFDSaz7sCe+GbN01dA8yqbyz8hldv9FmxXHt6zEwhhV80tT
5PgxxmHvoYAk2GiwqJ+gy/jbdSRhrx0Wdt2O4m1U60AbYsq1/hQn5jGOYjJkN2wY
SmHZ0c7HohWCGYALkTowexhvClSa9DVNkf8sIZRZfS3y5+KXs+4WDlucmkwNSb1I
eV8ztqg8bE8i7JVeq2x9wwlesyiBCxxPWa/nW20ao2YVk8Ji06LF1ZmLGFn64L3F
8CgrCcnrXqXnP2/VYYaXwEPsDR8JitPEvmSbIeMxEn0bF3WaS5b2YnMNeF4GHcph
DbZ3eQZ5hci8NdlvE6LCKgo7ajtfbDGHriZALne7a1TBZ8/CM2PA5LyEtTFj1KLr
jmDfGKPueMoWsH86xM7tDw8Atv+SEIIifNH/vEGsAH52e48KyvGvtnigsoXEK02x
8+cPOpDxZUF3TA+JDTtb49b6ZKYTs/DMiaWnXVe1VAtIqJ+Cn7KVandor+hhFl6o
+rG481liWuotF3XiHU+O7TxnnRIY4fYg7VgUSroMPNWKHNARf1kCH0kcFAbQ7EnG
kPU0fKKUUk024LI7rOjRydNZxPXqqLx21xPPgp8Z+/e/D8wYS2M3evlsLTsoSwC6
579IdX0izUI5z1fjSGwAj0x9tRomv1c1+O3bgetV0hnwAs3TVw/nB3v8LxWBljOI
p0ydGHzp7PdP1Nj/+eYYHYiD0SScSjIOpM+awHA6zXiMgpQ/SIiIohAYTX5iUJNB
sZvp6MP166weQpliHRGXFYneo8Q0JQAhnDqZv5H8h2NDiDYO9Tys64xMcbSQXQiZ
ndqHSFufvGBPH66+7luAaF2eacAW55MWKEerRQphENiT6x+YJ5hP5yq0cxnik75C
kqLNEjp2YwdjtLFqHMq19RvTHJW0wXs6qTrjGMpf0rG/bNVd47rpy9H6TAJL45+4
cRhhf5gO6CnP6fKf2IgNcsZMZkT8AFHzvbP3eort5XhSUuvxeLjFKDZ7KhtWZLlu
qm6wxZ3XTxLAwfRF9h2atbtUp0INnePX9Gi8bmRQfByVH6PglaMD/RcrKZxaX16H
zIxcyYTwawegxMjAVfVVcucvZJpARgo+1gTUhGiw7HVP57nVhQ+J/D10lRgtL+6q
vHyXilTWwKhoiSKh6NDGj9w2JIPSLyAns3VCVCT4z4DlmNTnGGZbBNZzKQ4Vtb8O
Yv+LNCMFVCwsiyadiKazCP9fl0WXPtBmNuqDpgQ8SeNFlEc3m/fmncTON9srCb0g
G8wPRMsbt7pm3N/BjIqnSpsryQJkUKGJhejKPO3xB7oH+/UGSFa1BX7uJjYmn9GU
/uxAwFNg1nkOTIFNLVpbtcRhMiVZsVWMY6n5m+Fy6hpJ0rOHCTlOcA+mZz2WGPeg
nzPyuT/4QGtxNa6ii2fIm0WvYBdCfQcF7vx0n1sudYA3wv4tVrdOMV7DrMHnX4ed
XIY34nlTUfyi5JNl15cwfMupIr73Fi0yM5VFWUrcnC9wR6Dv2AW3CgXhFu9l/w90
cwi7izH8JUS+LqD5fifooI38W7A9LEa2iOpms2nrXT23mg3tWnBIkRSpXBw8SwkV
dM2omP1t8Z/Y1h2xDRoU2pTQUJuOT6wpVm6T0Uj8x/bJpf1sL16v2F4QddaYvYop
uHq04sxhS9fBVEjh1LYVqeBQn6ZfNm+ZgvOeNRhAsBc/yFJz33WxC06GZkTgHKyM
V7pVzD+wGfsdxDyOl26mCo4614FP6iChnY0Zx9+MUfajQFCr5gpwzL+uvW87p4yN
Tj9u9owAaHk9XpAY9yWBk7nhtNWLkc4PZSE3PxPxHxsy40I5vq3BV7mrpbTEs0Rd
A4zcHv0MQCU0DLXRbZ9hG7i57JCl5WrfByTO1PhIYTBXq5ml3rnJi5P55MdkNVKU
hZZB+gbNF3jOi5cQ4xHkHahr/o6GmVYzuEO9x++0ukJFIOIhhCQ5kWQeRbXzTELh
SuWBPmpjQiPx0IL5tNOCkAm5Edkq6zHTn3uS4NnOyboyrP8Mfs3x5nZr12HTxFCV
YAAwk4fwbyyHh9vH80OYuhNpWIFRNpCBKwu8MFwkQVsYCZhskUP8bRB+LnBMmY92
mH3tpHimyKccJHCS9sQKkczyMKzSkfNOLuXCayR1OX0UsBmQK+lNVzoN1KNgHvl8
BWlCMSVOz9LiOM2rgriPg3vsAbLfNhp+ELDeWlLhyqGKOzctJKywx4Sqb7T0M/lZ
prbgAasN1MrHxdZ485NS4BdQsVA7S8uvzWchRjZvGqfdwpqzKniTSH+mIC04uN83
MjGD3c/NAofgqzMVC7eDkwJ78joWTMVef0+yu7gFZwy3+uZ0c2e2IJpB5kuDQ+F2
QiRHIcn04YlWSkEIz03uM1uT56lAUVBuavmxrH0ckhhiDSte82GAp/i2JPa6ksEd
gYM3Mifd1+CROLv0m2iN/mcqjZYWGpgbNrYTsOMiFyQcIWk74taeudlaUZvyJ2TN
6uM1jbvcCndz9J4Era7/mJ88tsHwGaI5QqqI08TaYFwBboo5Cla+N6U85zI2IaXC
376qFYRKHH2CGpnfpHaGZJEH6AXeLrOimCuZFuqg32v2re0AcD4t2JgHC8fX5uMd
fg4NCUvV1fX9sgJ0VJDb5a6eWC+LV7bLh+Y1rdi2NDKDJ/Lrd87ztfrhiXall+UH
1b8vU6sb13ETzEoyu32bWtyEC1gZCm/8AGYBWKLYRv6fGPYQs3LPmB5Rm9S6qmoK
cqjR2IOAlQ/G1WQPPDSbYRvuB8HtiHEctNstcWBjrgaicGjFVsS+rrcg8xrcekp9
JYnJv98A0xJ5BWpHkiRSJJEf2KgEc97MxSsIEHewPlvz4jTFLgOPVIhc/VIZZWnh
QlF26LQbm0riyYbgsA6EQ4IrzyWfQcOtTpWCzcvYZmxTGP7cIADQFNY3STKQVLbT
++NJNY5w4q45au4sNFUzJ9GMVbrIuc79L/9v5AWT0eOlBrl6MzmkSeJnQVndlGfS
UPGmq5jOjWMRA3C3KgIVlQ6MJJ+o4nAJVMD6uD7bZcDKzuAfmCN8YM7jOmjN4FUq
hBoiuWRlHv7US8uP3IEBmW7kWOc8AIsGcBzDuAOv18KelB1AIu12x48zOvyisxlE
CtNSfWPE3ohaRsQeMhDMI5StOU/DNyRc3Y+xQOg6E80+BnkYzQXwyXHIo6zGfhDD
ZLXhpsRBhEH9nMZkRlnAkXwvXXUtbehSmc1wOEZePw6oodbqu+NQ3lUEd0TnzRaY
eIVii75G0lVhy0MW7OTHW/XsdElhmG+RtJPU/Vm2LZ0kT0LyLj4KkSVxrmXfFD+H
PsqBSZl70up+rroM/LlLsZlTCwHrK0KsBT8NukX5Rqe+AUWqTG1A9aLacaPjmB24
Mh23Y8I9ozMZUSBpV44fqhtLNYebQ1OOZYLJ+nZZj4OiF+0UVj7jESom6OSGPwJx
J4UIu67nnave4jya6NxN9D+Tor2xum4qqsKgm1qaB0P5z4XUGu61Ds0Uoy/zZFCb
WuJ5SD8k1JTxpP/X85w2iN6yG0KUwIF/mix6OA4WtAg2GSFqI+ukj3OMGyiWdkMN
/z6D6HPX0J4Z5FHHR0BUKu6BuLbMXJGDEyEZs0OMIStFhLav45rbXsfNQ59CBKjf
Z9i5GZgh3bgSAHJRigWay35V7AJ8iNegIU/rPblEp3XHhyaRhIusCF17T57+JOv2
sVjWOPQZY9gbGZedk4v4UpDNbtUi2VFDDH58NDX8NmJ85mX0kzWE4MOVCUwFGCt5
dzZ6WgcuIMDHnb3u9p06WYibUSp1SqkuBjTYfCbOfCNEPfEFUZbV9TU0YckSaBSW
7kSR883kbiIpb+wYA3eMQUeZZZNqfF4N2fiWHB9sxAj7X/FN76ecPyUZ0AGOalXH
5IgRBQijrRpLXw8m0Pg+Gts950hQ/vo2zCgLPEMX77cj8/cqruknwawbz4L1uSjk
s0SUdS6+We+1gc0vwGdaQubxAT7VGqvmajerr5RJcssITcRhzli99haMbvhBcH3r
+WSBkGxH2dxA0jtGP//qmn+66NoubI0fTOE/p2QZa8J0WPRrLdg31RUORM/Cc7YG
OMmiaE1JpU6lZcZkDVnXquxTHDEj0aDdadoy29EShrvQ2kBAXBpj2dtXpJJrf16/
uAvsg61zU854+dlFq8taFLMZA1NjIyRVrtY81O9CRvqqBuR6JbA0qwdKdjwNx1AI
KmVmINl4of9hmiky5H6NAXccv9pfvKdz4AylCnj1IAY7w1AGUMSMYRAvRfw6FyrI
dk2juaClSSd/n+D5K5kxZlPsNiIfxR8mn/274SEbpweHz7UnjIdYAOVttta13nfC
Bkv++PkaHaFq8zu/d8zifQD4RuImXL6yIFgP2yx1jPS/qsb2A44jzCLwX5X7SvGw
pxugEZaJxZTEYUzWMWBtsBvjxesy0J8MJMyuCyRJ7tIQgoI+67OoPgmMOxOmf58M
PfhNvutD8wV78sQSaxdLbn3CHbFCy7X0XrVM6VdMugXE0uvvfZT23oqrYKxqjTdQ
VKuoTjALnV32Vha4k4ht6AiHQve94w77BExlTdBBjA84fBhALEpPgGmSnkkvZutD
Nv/RwHBR5vmjfYfgc5RYrcSB1lHBFSN3SqFf4/aMb9wklqnw9CVKd5Zc9JhQHJbB
yfUevKhtz3g8FSlPKAPV0Mfk7mEYs5ZOea32ASRtPrdKMzuCNb1X5eqp+Hm1C0DB
hVmyqEVGz687CM+bAQj4H4xMg9jNVyQe38uAxHtV11yskoVupEDxbVWB9m4oWB2x
eT4OM/Jr86Kc1dNjUihImrYWAQcpg2VF3C0s9UvY+lXK8nkgTMkdHawIAjJoVdCY
N3Cl8yNBqedVKg/MzBTFK5VcSM5dRrk0qKq6vHdQ0BzGSflMbiJMC7XhPZgSf0ke
Q00RKh+lti5OopRgt/T16axQb4ZSBnCc+EZHRC81mv+cw6JGvqgi7MBv2mXBdvDU
InngccCdD6Zrl6kysdYfxsJenqTOZNXAVxSL2gOL1dm1ASJis+D6CJkkOS9JlFVf
V5vllDG+hhpCcnXHD7HOa5Alz7B+1uj1w0tXlgkVD06/KsucQ51Ot/pwRxNUuWKf
5AButMZk0EEYZxOrIxcOaEqSL38B3XSV61vJk12fQwtj1CcwE3oC0r/6Z1bj0yWx
DFOWnFnVZy0eFGvc5wPeKFuOyaGTn5+I1lzv8u9smYAY9Jn+veFoZfU4qd4vDC3w
vyCEarXldFjlEkoo/HAyJwW/Z0Ut3J3q2SI+S2NCMGUHT2oZHlhhiCzJl8Kd8kUs
KyW+hTmE3gu2/DPmnCXGKMNVsv8A84q0HgO06s4U/L5qFu6cbPIVGTVplQbXXS9o
/SJgIgbywwkEYn1J7V6Bo43YyuZsuCPJ0AAhjFEPFieMdwQH7n2e+4hh3O6kx5De
nUbSfaWfhDkDjb9CAnGGq9xp3h7FwIaxvhWOG+YuzYx0Zn6JqONBikUwHroQCa8a
PKFBT/Derh9FJVdjRZjg2kS79kNtFAMcLIm8W7fqgJNTWvuaZP7yd1yJlR4hgrNa
8aa65XIMPNnzn+WBS7Oo57CuXtpausmw3Ps9/dEUcqZLWlUtuBYk4861Y9RB76sW
vN4HnWFHr3ThZrNhmPwLwxCGOIno7L51v3V2ABtfjNFAK8qq1Ar8VKWF1voQKy+c
JzLsNxgONaCquqB1SkG8hzz5g57b3bCHs3MNuNSjEiuGQQS5QNKQOb2HpK4Qu5tN
AMNqpPOPJyo2l1Ml5Naf6KEv4ZOM2XjOFTxhE7nXgGk+gG1bAazU0qtpLDkzOSrF
r3HZ8orwYsWT9aUICz3osaiwBGeF0zSpwOgz5B7z9REjiH65w0jsuwpgtYCMtReD
KmJOtLNcJJnWeadfRc97MoUYBMTjdvbSw4kY27Wm9LeZauYFqVXC7hfcNffCeT27
Ez54weObyPy05hZNXLiKnYzRrvwJzNaZE6Z/gZ/j1XEcs8t1c8cX7CRGj+VojPDk
pBbXcYFLSLuEQ6DhluVlArV4Obx+zaqrj6qOEJIrJIgCHb/JC8nn9s+XNWDJRddQ
5xDhH16v2y+5mnFeqTjM+HyML9ChD3pbvCCKuTtm4CmiiPMF4jwqUii8C0bDLd3c
8VEf/ptoofmfaCoxoFqmoCX/C3zJpaE81hRYh5AjBHcZdFt8LlINMgFaFMOdRFr2
12VMsDRfGCn69th0d6OA9hNxWD5L4efTdXc1uccaQtAUD2y6kEZtuCQHqhLlK2VS
SI4jqUR6X08dMf7ySxm+qt6B1+43e7HE9SEXQ1UapNfF1Szl0k5ET6kjIVh9d0oH
S9scFAbYi1Py8KL4LunQfiGtAo/cIKbN1J1QEV6Qw0lOWoh5//zHeFtw9Nnqgkac
i4x/Rx3bw34drcNRIfA4mzPB5U9ayXOeaBeLSWxwbtXe6xcHMdHaluKn8sCcnbFc
XCHyi12VXIZYWGwoe6sHL2EcM//oIGIMr9gN5D4RzLpOzAWvY2mY8dOMRxZ62ONI
SflByYic1oLeKm3duFqhF5wM5hSB8BeviDCd202B5ITsPB7QMENLjDyJsKa/Fk+6
OM390XT4MIQXpLjkdSehRg4pu40tsdLFi2MMpnKpR8dwgOrX8f5g/g7/6M2GNDOw
UnQst2+PAZ3DoMVwbovkX7YSWWz/dYSsKcJ5L86NC79dSlurnflLt1dfxAFTVo9n
ERFoywwWi8I/1xIE2aT69HZuWO5p/uf18LI2nIK/PA4YjzUuyUPb6xbWrd9BwRlX
`protect end_protected