`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 4560 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/9huKRhRMtvnNqb3Z+UU7TahEoHV+T8U3P3ufru7l1O
3DlgtZzb9QxCbOjthp9+wDkjygH0eUfDrEl1ovhZG60cncLmTqwCiyljeFK2Vlgt
oUEbe9T5e7/VxuqShH29JoUfE/91PQZM/1pQgjZHNpL2GtI6J7XQs8h3AtltkJR5
Q74Sm8aULmvAVnPw7u023dm93LWBF74ktq+5KQP+/IhfXY6ll7iU/n39ZMU4cK6u
KjQgo5eZSMaTcY7UNVQZgn0m/VivpBnuSpAVloB9eoNPqPKJXsibp4CIbp1/JbkO
bOTtb73q0UI7YE+dVsOUVoXRAL04i41GjRDjS62cCP7xYl7rspEFLPTA9w4e1GiS
y3kCuJKOJjV0yKBiCgg4FfBs9mwzDXsfnGO8egJgCBxaAMHPHvpzc6DrIOfUkUia
LMH3Bj5k8Oy7mO0ZCtIkepkuFbT75/we/T/52n0xvGvZQC4I1bp8+HOro2y76l0n
WdAVjGLPbO5qEIxzaH+XnMX6h3adlCp7vGRSimps/L5bCNo/FCgvloZvs2YkIhar
onigPo1s3A2Min3PDMSlEoVxTrw9EPTnUuBzBZZQ3fEDly/QS/loLthUiid8DP4E
A95yULyqyE2yvvY4IulMJO0iA4aD+1CghRTtInl3Oz2p3Rnvi2Sv9PsFVB3yBe+Y
SD85WrfYdkldzcekdz/hAYmu9Vg12Fvl/+4eyisxB4rOb6gtqUoBBObia/ev3cUY
TEL1VLbEltn5HX2/a3DYWdnMCdr8eIHGSepffaj0p5A9yI3RtP9hKa1tMmQdzp/I
bw5XEbCkwv46LMy6GqY46Bz6syZ+DIai2+T4hfbD7nopoE9+cbEO0DPxXDSLgq6Y
EmU4Sgu/sYfXfy+dYKeDR3WA/D2KO9Df8oPoIdZai9LcoUdRoCPDECFX1sFOzCwU
WzNHuaO29rE+3+UScfliqul/wnv79yy5+OGJVUDf8P8vQlexljHEKdLeW3xBVA8c
qVaxEiOdh2ywK4wEaztY1ja18+A75IPAXqlq8SEL++2yD1BX8QqS79vn3N4jWTUL
8CS9dKZgcjvCdlEMhPqSLyXh+Po97cQVqr8TfGha9wkWw79HPJf8D3qC0UFrpBrA
F14pGwh4eUKESiUEkA/A5R9E6Q0IyT1VSLkzh0B0941b/3hcbsv6R66C37juggcz
F3lE8DCZ6zHJzksEz0pKXkUikkAbiPb9NX0Wt1D2HHNnOU8jPATQ6H1Qin3hWA9m
T/4OSi4u7PyvxDejGaPupID6P5gJRaxVSVGuhQYWsax62elsKl2EkWyFG8Q6wkpe
orTQOCS7IZFdDIuvWwWJLmoKZ+n675YYFVNJM9IZALQYxTE0X8YN/KDUhYdzUWfU
bqOfjmvM2wvcwsBdkKzdgij7f9PgVe5RF87QZdwlmO8k5xpvEj6lnl6uxJQgqbkL
zahwKFqtMSMGuC3cOM7W+qALgxxNcqNZBniqjSC6VmebRi6wMrKh6xkwztu6h8E7
OqlClvXJcX58lWvt3DAnucYJER412zJ56NW5H1+3IqcS3ambp4qWSf2bqNO2x4V1
Srmmi2dHJL+u3fE1m9jv5Uqvqk7tJTgw4ERCb/bAHfYDrJJLYMc2rI6R21UNwSm3
+FjwXOQK8FIV3Fy9kOV4zjuHoSmpbJDxO9MR6HtcoAMMYrpaGrrNrIe5pxBxr7Xo
nyJBsz+yVOUyiv8r4kncD3ajrLZApPNSY6yXB1eiwy9HVoJSbx/4GRbZTwXcgWgN
O1iZ9e8yf6s3cCJTEiO+0kO2z3HbdEqzEIcBckNUfmGpWbh+HAabMyvAVYZXJQTu
Cqvkc+ADwvWghUt01boteFbOPZlpuRsNJI1Tp4/J5ZVbmttxy6iDXog9bi5tmKaD
+PDX//EaEvnMOYrXUR7WAsjaVQgKHhPtdqkH22vC22sVrYDLNuzfHXiMBW3GRUm/
2ygSTumfqqIN03hLshVFOMXv3ZxhicyuU5E2de5MkWxcOMutYaaIdRlfaH2nUChS
AeePixAqylQ8/Pv4w5mCODINtI689amnQ2H8BHEKmyLDgMTzTYHVsaCpwzkQtu6K
Q7Mltj3zbftq7w4Ejg/zU/ewQDXZJda11Gdy/fOiZEFOjHDFgHArPcumZcvvmAVr
vz5/oiqNfvw5DLReoxoESgkO31ZPaYjbsWwTOMuG1se32nIK/n2ExzZ7NFyjIQad
rnYZBEZj9pGoDsp7EEXvIOQr4CbgGrtO/lvsFSgq4igjUlPAc6rxFsoU2G/MXI0/
5u+UHpi4cqtavKRmJXLX4UyCXxqY0qfqzA0ab8JH/yvPv6X/cJluNXV9HeRQewzO
p4uYjEOfS/U8kxx/mMoQAclt3n6TKtCTeIhA5EvQQ+f4RDFsP3lnxH6M0TKUtDgW
BJMj+VP1fn0HQ1KiTEndNc21oBoC+STLWqG4B4+Lyibj8JIDR4DxHokR3K9JQxL+
Nnycw91A5mMQk31iCBe2ndmnTGuhTIN9wzlTMBNEmlKnzdFHs1Y8gBKiitUXEMEL
NuZNVxuFBsmfGfxQfbiVdsRV1r7ZNOeLE4jEhT9Wzhb5fdZAbJufkSVm8jMzyN06
yICnS0YVO+beYycKs4PubEsRYUzRt7WV01WNNm31GS6lNy4F/FNqKn2OIfgnBf+2
VyengZfmBw4jwE0huKgPhY083FINFpb6/ruJfkiKael0/WR687FPXsQR/JTYXKPS
F8HNc/nj38NERmCzZ4tOf3OQ1QnXA2Gcyn+hFl8jb8LA4eEtguRfOxlTTlDLL8Mc
715hrlFQN1VGXgE/ede3HJS4zmByD0TKDC3tAlWeMuznLdz0CtXVB4xVYMwtvmIW
3RdVAa2N4qowpNCgJmSi89mUNNTEkoEJvZBQ2pM3+RdbmPOvm0YcwNBSjF0nPCuX
w62xH9tt5oDcHSY2Z1G+rku39w73qLW5wJifcx0bG+u8q248ZvEhyEVdBFHiHHGM
mUwlsK7tZDJdwZ216zvdpGs7G/OC6M5Yk/966uCDF0stt4X5fDYjXg+NiXwP/Idm
6PfKI7gLiSLSCeey1odN2xXCEr1Vk9NoffDPKIqXWiktl8OUXJK5IFCJtG/Xa1Uv
1HVIJI3Lgnwk+VCE/+I6sHBsN1juh0qsibbRhBzD3sD/ihZs5NbtTONhEQvTuWDC
MMHaZfr9S52sJTkVVK+0MipvzW0r76UCiuUx87DOYGYBGsP5I3HJl5/4RfS8MnWv
NIoKl7H8x2VsK6rQCM7gu2wRH52mxVSt0BZxaYz4ippC+NFucs7oFF0+KwysNOf4
AELX1xv7cuavrFEgtNQlaf3dfCGD3IAzGQEcJdUI26fe2jscijGHXVXs6jpJJB6M
igpK7tIHgsDWmxOLn6KFIiQELWJyPo3sL+dLQYi56x8Aez0vk8gtoMQhL1EE34eu
zmCo0Z3BEFBu8KaKLq/I9RQoLchTvKP3fCEqIyptxQscMe1yM1+iEOCzZzhiwZgr
wcQYDLol3jaEapQK9cheTpO43aW8Rt0xWp6rpiFDTTsEH2+RAt9gwJjz6VbFWgiU
TsxAuJmIMJady68VOJ1C9CQBdkeCb1gIlJfMSOx0tLqSTnsN/Vl6Bk4FGJdgphNf
viZeECnRmwxY9Qp661H+IvrgaYICQrx/7UwgjLtXZP7AdTEfM904gR+p2vozg51B
ns4eh/eUmZOxL5U1cmITdu6f5rISmPdOUjJz34kMreSwqFVlior52LMCI5jJAnC1
7jfkOGONiAcSUwP/HdJgKBGZbF0vR67vQ0OR7mg4pxx6Ae69Fc0ggka6Z9qDh4X0
HJliiHo+YqyRXzGdQ+D+wL4XtyQSxdLRGhaq+7p6jnyoygdpNLcfxDS9aTFRwiW4
BNT7Y0wsOLBVdkXTMaUcfvwpql+XbSUOsbPHFS7hYcjCTRWrRL2FfrupevKl3prf
73LaYT+UoPxi/ck3iWLPd64NOcwaLVAarw0ysxz6GHRK/MxNhz/OmYiTlWGkntjl
6uyUPjN/iqS+eYhjEvdDaFRVG5sEIxuOv1MpQABKdTw7Wr6Hb4lcc4UlzJbS55Yj
u0B5qv5MhJNfc7/nndALxS45RAcoM4iZSHAtpIj5GqTug33d1OzjzIdmu0pfasnQ
PpxomPQFoH1P8pVViIOPvbbC9RxkptVbIJB/u6c/yrO1WEukX88F8egOBI6lLndE
Vh3+85iXDXX/ulyhuhC4D40d/VxX741r3+6Z83J4xlwQXXmPnjWycN879vUUJIV9
vZJMmkSGHoBW8Bt2MdLsTHm9+IMhmmRhoacRHkShPFiQxGbyoOiOu4jQQY0T1440
VOHaTG+ITP/Rs7oMKanKoTJXLVQuZQCvy3RiLv1Z2KmD56mRkhyPhjYgvE7JQnLT
QjZEx0ICCdsfQ1keEvE7tLtEpKOuPuTnMPMwbx7S+qoSBWkNKj8UZVwZcOQ7gQX3
AJaUyVp8V6pcv4+30VUQZLzayCH7iFYanAreRCUpcjgr+iQs1Xf9uOwHm3Sj3n6H
btOwp1SWs5s6hcgz0gK0gegA9n1tlpc8s44DDzTh6FxNAPhKxTDDROAZN03aLvnC
oIrG4/fNt7hwOv2UI6H/P1Fhi4ACFIfOSp7gtunQzqKnwJWxjksOkn/dOnudldJT
78q5HhxbQTPhmSapIkUsrau5JtnshDS06V5o3LHLjxtkALXbnIuYdPOg42onaVmM
JsrTMWfHz5c+Wsgr/DXE9QI9C4bUI7m0Rbv/IBvXQ7RdwZpYPjy2/SNQHCZJkWE4
MuS+DssQG70wcxETGDVR1BIxaFrlgE/dKRi8ziUhtsulUK5uhLKPXfgivV2p75Vr
Nza+IGj6SmeU8LXFvVMYZfFeBJxOI9q48+ppwMoBObN4xzvdbsuiF4i970NCAi5g
YMXvgeQYU8drwOx5lBeZM1DRGUbhXB0oeFD5VCvycDvnBr33gj2cdBiK1QlEmFdT
f3p2b/bhTP+0mAiNPh1c43DSrNQtTSITiJBq9wAHI2TmknhNz3nCqNhr3TutNm+7
81dAuH1QbwirK/diCGHyAGg+G3FUPiHkkM+MrXEygIs+WwIg/Vb5AQLTq3VOlm9Y
ElJqT6xzhpB8Py1KS1PfJm6TtHYJpqRIjhI3Ycfzj++zP3r3vee7n4eIPWVJ+H9Y
H3hCNPcmFZWO6Bo5EJCfx7Cesc7g4+GCSfGhObykBN3XhSSnwogwwk9cXvt7V7OT
AKK4a/3ZZZ3pK1penZXwLFf7yoc+AT5iDxaiDKjFYC7P2gV0Puj+A7HUpMYuLFQH
LsIpAc6BpTM/7V3Spf78Ohum8glq/KXhG26eN3GKOyNDLwo3Mlxvs/lLeGiCNDsB
HSUHYOTWkSX8j/7qh6DYq7tJnR0+OtXQgF9SyWd117TMGHabSDE44m+IQP6vyDlZ
Vq+x8qprNdxmVcCtmruKJQzNlV+0LsOTi+p0KR5Vo6oaQtuNXEXe2LMNxQkAJIkz
Ybf80noF2tWK3yff5s9k0mJoWl1MJgjywH5/m7q9yi+xbPag1izLFEy4oVHQ3A3Z
LpjeirLJhF0EaWIBW+8cGdT5gyXmdYNzacHssPofUppxBak+FUdYokN+taaMIw8M
O9ljolLFC5teldaAMko8HpLEGwgSD2sAkWk7z8iQurUpOfIys2bxVLWd61VQcGP7
jeqrzsPlmOVKKoJy6uUGSAAqCSVCe4UnNc0D0w4AFdgjt2v0i7C1bz2sBe70eBGO
eriSJWxD2kYd+h7Bh3/zAFi7iNQqIjUOOuTHZN7n5OIW/BI//aZkp5swcRaIZaPW
u136uQEXOqevTnYIyjDxQ2lp8agh4w6Pnf4EzSKJj1fy5X449Ml1QxJpMmjJX1k9
ACyN2a57IJjICTNLEYwFWefAGx02N+J6PU7PZFOBgjfwhxJ2dglrN1CSxGDLLyxs
2WKz83s393R41TVnhceL9T/93T0pqm9+niWyuQJ+a+aruS6OR1lhgn0NdJ/oH7N7
qQSoib8cYWvYY/8dZWj2eH/ALZ0UdXF79R4nLfEvJg6ILq/mtZ5zh7WoMpCjLMFx
`protect end_protected