`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 3456 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/9huKRhRMtvnNqb3Z+UU7TahEoHV+T8U3P3ufru7l1O
3DlgtZzb9QxCbOjthp9+wDkjygH0eUfDrEl1ovhZG62sV3it8TjPFt9YWXJrK945
AQYfRL+wuRZOrZIq9H4zg/h1A3fAXFqv4ToQyXZ2tnVd33syUPs8irx+BNw5QSmR
9tNx9LH06zrBJTqxmqhnfAsUwBydBGtLI9zhy3KV5H7ShWBBGYQYY9uqJ0jhL4Fg
C2N1Aci+IOTl9O4Rj8el1+FHeNUsWM1uAZorkYu9g3Vg45tp4vA7VUWs136V9q1T
b4JdgEQUAHUrxvJkwYVaRjei64PUKX9YnLXdY6I2IPm68EiyEgMBgRiCdWuZBsbs
HPN/u+m/jVocgLTuk63yU40F9tVhhtkOrAUDgtRJfZkF9kd43kzliTue1hkOYVxl
tlcLt+06kC70kO1KFAA0073eefGApWFnargaVa1s2Fspq0k+/GIsIvMeSNTKTK7w
RqUJ2fakj0mEQo7TfYmB66zqkvQVHurF4XcJecJsayLxAKAIMRoKE+LsQG8NYW7L
yCZjdr4bLtbkgVbgxFcOXW2AXhvXNgsyMlTm6yfKtbPawTckTOsZrb9lvzNpV/R7
pOYSPI0lTCB0M2/JXnsULEIB6fFlzpS6rFDVwCot7jvcwhZ1KudE/M9SmXYpSevT
iGhdCIDzAoCOriEB51BrlkfS8QI+OfAMrEyJBScaiXPBt0wVQt+m+IjWo7RF5tnH
AomwPbK4UDANwPrS5CegQDHwKUkj0fTQfiyRR5ydEBZcCFENuTN3QM5yGehOx2qU
QZSw6BweTanibFTQoW+hTLyby99H/A75uizNVBouexq6qgMcq/C3+6hesCrJ8LrK
0ZXF701hl+cwB5MmsEIkvKC9Ev1hSq8rMpzdgt7po351Usi4/t/VOdisZASfJJEa
yIJEzt/mgE8vTpErzv1Gfi089GrmSq5qt4tqC87pxFAVYx6snSmWbS+prfPw81WV
MrUx9xa7N9vctnKTpmJ1Bpzz7UlWn/Bkplt4ZFqCgNBA11q7gC338FibMNX9BhJC
qydRBr9gYiZzmY3tF0gPMqbKPoZYpCwRGhx4EkxNSbq3qlFdHAUky/Srsjl5xglx
+1oq8JDkc1P8WKY1I4qMye59TAj0KZrRE+ay1ViovF5dminH6I38xVPuGSwET6PC
S2/kzvDMhF1ORuL3PvoLQBjjCo0vuSnUYa4jjeb97MwXzwBOJ0I04NOprVa154Z7
zGGPphu5n3fFiLxIpB6dUP3LkQqEM4h6sx816b9QmJNkfp1XgPs36I+ZcaE+wakz
2bI1ZR+dbrichV2M2LxMt6ejDf2/1NChrF+wqD0jIRgcwXQDRGzvj6txzyOzoIgs
MIOJBbmNM8CLCHHFUBqT+9vKig1hfTQVWqqAHZP/qK0TH+ppaMyW8zkCXtCXMgKL
mwJew5tMqvwmbu4oXcK5xrJomuDL0c2uGvcrt9Xqz4c2gJ3RapSny9tp1zAApxJ2
EcuChE1GrKexYzWxT+pqeEjj2ferHLA8mnvS4UCr1V/cfJ7rRLosySLd+kkDnfEN
FhjZaYGQNXC3UjoiphzjYWBwX7AScPi7m4SJDhruFq41J7pMU+oZkHdtVVCG9uSC
w91ynRGBd/sLA0mfEeyt3TeVSCN4wk09+MOK+yqUq0kBV0OhLD0ekAAgatkehn9P
s6lXbYYRad5Lb9F5dCG/WxYH3qnx4yHwf6Ccb4t1kTrKb/gLiSCgukAWT/YWca29
FVI8mHHEJ1POb9rYD9lvXP6dUN0XCcg+zAye1a+D6JemMR/D8EyILI2y8x1+nNYI
k2jd/2pP6kRAVc7WTKPAzAueYgCEvlzERCstym78dSSG+is1tmJF05s7N0MNCCiH
waqPdE7p364jqhx3kNAOzLoI1xZrHxHOWS79DxUjCER5wNSBLN+5i+VVYlnLDdTb
TdEhTH1WWNc2ptrue8+aeERVzfd2AtSSShhFslLrE18S/wbg5O/ObpyHzUtlW5vT
a5mIsAZzSgz6itJrHyT3o32ad3ve+95dLRUt90EFcbMBlOHCyekObwHCuyBbqv+T
lcVhaOvhcZIhUOgp2S+CQ+DrbfXH7T8ojOdiMoYionabdY1mTMkoYCRgRfbWhl2v
FEWIYAP2h6JSXoF1QxoQX8ebiWR5wSJMBHTS7JQLTqokE85PY5R4Mlm1BpeE9yxn
kB6UHQYs+n0tEBl6qD4iHRrvG77DugDRUMCW1hK01JzaDkuuxtwwLjnEgcqPVgNH
khuYDxCDHIL4wcSN0/5fYEV0K+uX0UF9nCUeY8xQyQ3aKjBeLRTPScL4u6qWfZZ8
xzIxwRE849eCyEmBSu/XeBrKgEp8hcYDSTK4xF4yVzoWff53qAvBiuvROhVcDdIm
A676FyDFAdT8ZcSl77KY33hs6DRvYb/Maw8XuANcD76kdw7aQDfLFAzC8RUu0KjU
DWfAISR8Rb57AF503bVv2FJFyTkwQ1F4H7fJ4tddeRk2YeDbAIjMOvvUTw8ozqvZ
bHHv6CuLUzLXdg7L28WqYCxjiJrmFKqiOylFUUEL6Z9QoXDIQCrijH54qYFVw5nZ
cCnjA36udgVGP7FhJ+eNFvPXm3AxEqI0l3dGJBCVPKzqb7B+QFHK22vwiBuaQwlR
As84osQ9Qq2n8Fa++qhOG96NF2M/aif0VwLB0u+eX9Ah2UoObPGV5YaONlO3SL1W
yqHbSnsT/Hia0qx7KeqkREjpnRYb4j30T3uVAaGQjl0sGnnv0OA/WT12hpNoc4+Q
9fveavZzr8oEt9FtiSkrdLxPVUGCmSDWN8bg3etYWJzfDIHaeCY99buGBa0lKwwO
6Vc/8W03hBM6janJJZmXYHYAW2Vs6jtXF5bFLLn+uCEU7/ajj56Gt3RAgkuO2SvK
3Hi11VO33KIJQIJr6PvildscDb+3gbMeLb0ig8Ll8VJrA4RVzQmcyZxrZ+QwKbBA
oV/7NYci3Rb5hApWwBdZFqE9yHoLry4ERNYPl06Y2d8AVYE3HslDAiKIlCYWKiI1
1grT22v78YQCs6d6oSZg+YcMx4rUD+x6LG9ufJ5m3PIGbYreXeVXUO5DrA45HAzZ
qYleldp7KGtFsMWa2+D8q2emyYWJu/txtXwpesoCAT3vwgSBx5ByLAzlCOC9rPhS
1l3YQhgfm8Ilt1JmCfO34glBH+xMji4niI/lfJKrmJFmVHcQ8jMrkPktMLJN6k4W
YQq4vKxsp7fGbJaTbW1qoXSKS7ZzLf2u9sarC9wK0RzlEACuGdpk+qqT3yqseAyO
LlNLi1xnADQEhSapMAc1VaZtzR4HquCFERM0+JtVe2Lr37S/wDiKZ8veKDq3YMdB
mRoVzyYC3PLoT9f7/R9F5YB7o3OCrB8lS79hywQMt136IXgRU8T9dNnndLGpm46z
2sMabcBh8IsLLgCXy/rkMdBNMfdgTjVR2TVAwygBQ9ckzaa5+uNLzMPsH8l9MoMX
KbQcSCaB2z1A72Q4Ykmwm7PxHoTEF3kfEuJx/BtKjjjauke0Ce/eI3DBveSG4TpN
pPXydboZyPcq04DgCZycwlSoDFkZtH2iqmqB9FhKc5cqX/eOCGllaTA4Nmraw5kO
fjJ6EYo0msgzeGoBXoC4sM5U+f5R/OIIfGOh2hOZnWL1tZBqrzzjCV/uy6HJ0YpQ
FTpccTYwKxn1yiDt8mM6UN0BnVYRBpe8daQq5NExg8sxqPtlOIuW/zSL7Lqae5YL
F7HtyDrv/svoGZP8oJ5YinUIvuR0tlZ+u1M8t60Qk4DRdt3ozxfuq0Nk6HNPpSwa
F6BaKxfeWM5HtMOMVUQxoQdPEpkvXpv2piOZqg0fSvTpz3tioYEXddgSRouh6zEV
EBspjLoyUoenWsz0JQSql+s/HhQrTESS1B1ltP2zfC941eOW0ZdXAHi6svksUXkI
HYxmeVQGpvXn7emmBMNsc4J7xlRrezMVGe7GWCmial45c7oQs3OhT8DC1lG9whWY
O+EG1QOEpfm7iZ2ABOxWTpN5Bk1gkUppbYqa0h3mnzZ4Mwsm5Sf3Gf39/OWwscSP
pyWkBJX5yIjpofU2R5VPcHRSK+MO5Q38K4Z6ZSKkFaIpcWtHzibrQaPhpZ7IKlOF
/mPY3egR4Q4PWOjbRn6DtsLMRPvXeS+gf4VZtMq1EBXHgkoBScYpprLLP/I5ES6q
ClL3pqQFCK9ajhi80EyzvB0vuxwBMT6wTaFiDr7za7dIC/HSLAWhjLvlEkhEOYFt
j3m2n9If2+h81g7Heg85ZF5pIEJP+5viHJ0uuymx8TgbX+gEXDDLXCWH4/xWgaBI
vCrDeEpDxFJB8dhg3np2A86IrhHR2ANiPePMWc3nxRsH914DxULDk3nBgio85CAO
FExb4c8Ymrf0/hvtHWtY2a+RM7RaUA736v6O6lMS6HWM5k3OXk2jH6BZgxAx1ddp
ohZ78t82gWlMG1ehMZhlr9NC/U+AwYi5I7IXtnybfwXYPx1lrSYRTEJ0qjKAa0JP
YMQWG/yHtb+xDyrIE3picnU2TKdtPxpH6NamDnz+ytgFedl6fsjtveP8VDlb5n0H
`protect end_protected