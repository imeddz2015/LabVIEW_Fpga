`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 2448 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/59UwEX+aE7FohaWu0/8IpTj7mav863zUNIsgIH2BWb
Abd9opeuBjbGF/waQMI2vMJTwD1ie1YueHc3nSNpEh4OXp8P5ybZFY89uyGz3ztU
W1EsuUnchJoQgbHZ/sLbgtGRgsrAFn+ZoIeGN1d6RAF2wAESJmYP8zw+p00RvjZ5
G2ATm2jrAjm+J6bPpiDE3wSiqnk+EAkWLgqiGLUy46spyf2ygAnhzezOH0C+hAOh
kvyaXUfFnbbpmHz60lO42BTfyNyC415C5X4M0PTzeyfvTvE27So0ou6AWv+DukV5
xKnJhM7G05vabbzA7YNOEtr2C39DdM8MdComvByYoesyBluKBA+jkxljZdxkdJ4a
YkA5AcLO3+pPVptEPTD2nuJyEZv/duTBIovMwpm6mdjiAu3+NgF0YxVN9ZE3QPss
6AsJtc6WWRCx6KTwNKjdJZytNbewAO6i8FSdPQymkLe+iSTSeNaqMZlMnnoOxP2U
Dlr477+5j1lfEkywa4wtrVmDsJKMoDcy37jP7nw2uO2MZOzmJCwf0s1cxIO6bZVo
kZxH5M3N/repXRFEKw+2qFcbWlm9GuskZvn/SLYQN67v7DLRTrv5APwvJA2gPXF7
//MmrMX8X7hQh5pZ5wKem/CyuoC2rvbaIX4OkQdV690eu1XVXFxkaD64HQkoBIUg
r6wZTcJKHLxhIM8fzHNHluDyuwNj/4G2l9d1WodPj7tCaWbiU1h6Z8cxg97AvIAD
ffijDC1BuWhJSyc7lJrLnirrpp4MPY3qvk7g4ls1yBsoXoqErEWd0ZGwjujOlK7K
FgudD55LMk5XofcqiQt2u1inOfLtGq4MWl166XtMpjqOhrvP4jhcCKrClsfX36+/
dodaxwqRnMVp5nf557HKYGCmkbGt/Zyw/WJHsfvKq4mla+5pk/wtzZjbPfK87cX5
Mzh1ijangIn9kVYgTw4iYrOEyG0JI2dnSvzDwXA6s2M29isUJ8vGOa1+Lz16x5dq
W5Y3oHrIxRls5kX4J4wCGZVxRrdCv/AB/+RM20vqw2A9il/dQMa7utXnCPk2jOIi
mhVo4sI9x5YWAc17d6c4s+yQtCVO24Bu+d343rxGoZNxpOlDiJUSWkYYOw8m/VdL
YEUBqyqYYE+02whYLaD+qmh0Bs1WmNkS0K/C3C0piNY56vbT+QAhN1yM9GC6f5ut
FHQhOCF+Tn0k7lRDW8x2M6OAPKHnyacdBUDNAsz/Cb8ttLqXxXahhILzE7xVBhKS
wY4cWRx6zE5fpqAJvI5A0hedkGo1gtGNZrM2iXRfvsAshSqvJIdysrPGIVMuC/yc
+9T8MvbFDXtDJo1IyUKx7K0hr82+t2qmg7rJAqyKS0MK6flqRaAcymCekfzY9GMS
YaXLJ8ohIdJjleHI6cR3Mo4zsiSgKNfi0LEjTiw4IEQsBR1vrdKqyu1TVu/AHBHZ
AYPoFGvIYQ2IjxxdN4V5/Y6kDoo3NYbcvFxbfQBIHhfdtUxg7pixidM5gohQuo76
vdR8BFe+NZT35liYcPbkqHLXptWMlVoXKBVZhTg28JK70cI9fLs1V2myd7loRqwH
3872F7KyJxwQq+beNtYsrazzBtijiJnEJZNQ85k1AzcWGEKImnQZENUIrcFCeiya
ku0LeB9DnWGDsrQW/MsachUMNmTk0DkpTg5bqUFdIDwEauqB/iovSW3I/ssxgouF
ormnEh/QHJBx8sOclJ0ZHfmHID3BmNOQB/KoHTg2AKgziPw7JEjrm+AjTpVpXRzR
eJQNJiwRV04SwGhk16yQ2f5fdLfKhGzv95r5ClaZPC8tvu52n6Ba+8caVYXLq2RJ
wZ/l6R7dXX8ly0pt+ULhbCxWRcCdI548i1c6zTTZkVbeXyWXsmG0WPWHI383tAYb
wMyv8PRgd2/pbeP5iSKW1Ix1IAQ56JYOUDNEM0/X7ROX3Kz/+udDLAjyP+Y5sc2D
8EetfQnDTrSLy9S3iGHRGBivNoTguVK1CozikUV44G5Z+0Rur6Wx/x4NeDvHnVLd
Ks0znzbSs4DkS/sf+1GJAZpuO9LCoDuBV+qHILqKkQAd/ryp5pXrmxY7K9XNYG4i
hdWMwsWzHw2OY+t9QORreWJRQdZtyeBxti9jagYXE7stLRdNQIT+lyy6zML5lKjD
krxxK4PnCUCWIbfZIYNsRoa6Q/n6qU2JmPV4fHulADCLmSGAqENxaPt2GFTwvFZY
JbSfPtM0sveVFFBMsqIUKDDCRSPWM1WEfh5x5YUAMcpdtwz0qxB3m91v0fFHHb38
kzxQN5FNnUAfajAjalneQTXh9UuYkCaDIRAD4gLH4U/1Pm7p3W262x8q5ssUzoew
2kKYE/Mxbfhizxpyg3HKXDdSAs+dNtGD/hvpQe0rfqVP5ssPolwGh4HZEa3/k/1J
e4kBSB9s1MKV0UZHFh9C6RxytZt9LWK5Wk4wcAoMfwReeSAQGgSRxuWNP7tlQcBe
lWLd1TWUIV1pVFpAKwXiF5bymJRlxyhRfeD/izRvvQ/m9CdZxR5SjR2U3Y0FJTSh
VNOwY+3ayMtBt8TfgcDuz/OWBfr2pDXITKFZrTDHEskiVW/WFVCwV2BFjHlcD9vt
tsZ40+WKp9dEQ1DU9EU/8gD7+ESmf0qJDaJ7hRd96gwfNgjmjLDUU4vRHt3EaoOy
2hLUzqcv1SrCkL1vwHlmoKyjNyq2SEFPlXNw/ikkky3wYNII18fo9hgUZ3BBVvdw
EzYvxFTms8m0biv4iHPfe/26nfqn34O7S14Ems7GQmV5kd9jWdcnLww2iIy2qtXw
Wmac85RzUakYVevdQuUiWIE6q/ltiSkeK2gDvjh9j6Y19anC2XDYRLvn72HFMMkl
2YWQEzw/ohxkd9/NBd7BqE/N6EVckPaxqba6TpwjE7sD4sFaC+aILmTh52fdkPVz
/uEjWUebE5yBdF1DRrcezGsKo6m1wJCRSJXFJvmkRXoWvFB6dL+Hj3Ag9kv3IdsZ
WQsw3/qN6uLL9K7uHMyPfh2s9fVXYf3IipFmgW4iMlL35xjs56E8l/99cU6ElMeG
o6bQx8MEHCkJsSnf+b5r9eQbwMStTsYNMwVZvNUezHrPtg5SqHNGDd8N0yIGlJsW
oKSxD6rdWDgG+euk/1VqAqVw5d5ANlIbU/5GNWf7+9W8kb5eN92eEkm+xrKmnyXs
BgWO7ml+M0z/lhkKQP4hKdjG6cPrd4aWrrjvWiF6DEPI6dLOx562Jmpvi6sjry8I
`protect end_protected