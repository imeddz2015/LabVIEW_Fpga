`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 3472 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/9huKRhRMtvnNqb3Z+UU7TahEoHV+T8U3P3ufru7l1O
3DlgtZzb9QxCbOjthp9+wDkjygH0eUfDrEl1ovhZG61zQsk8sTLirEpRg6+Fxfgh
kIWhtkUUOm1OV7WHM0dv2kBSoruElQvXNh5YfiAz+D2VcaAFQ9nJHeLGVoj22YXG
okkh+gu/yTlkJGTuo/XtROoROIthxvSG4QjHQB+t+SWVXoPlbCHz7KavDC1gu21O
h7d2u0Y/MEJ9tEC/Rrnn3bp1IDh/4aCn68ul1igS9GdqzuSzkAAY582QzNpTWkC/
wrHQhFXSK6yMnWqmQPVNXuWkOU494yAUNLJVYH1KXCi+ohtBtEHPY2aniILCEI94
N5d2mXXNQrGc3yzrlTd+Kc1DRXVFxZ66FGguwzgH+RWr0ufcc+nTFU2qBbGOGor1
CerlQ70e5mTG3TmhWxFTZ7zgcWwQO5o0dPWP5L6h0XJajfzIeZbw2WqkMBcY1aEr
y5X55ZHqB0v5ndxJC9l/6vgxHhyrwHLbo5zetJLqX8Ppwb+8mXMs0bKMXe7xW6fL
6/a0hd7KT4UFg7QAB6590kxKJ9I10pJBcppIWGzZxrVLj5suJhL4L/9dq16HsG5Y
jtjfCQ85eeb3rue1GRS2F5/4CC930LJ4viGPx/uFhbY8tXVP6zCE1ISNX0dTTGNz
5rrRLFSOwRH3IRkGNW5brQYE3OoSB41SOFh4O7mDNsa3sw/xL2sj8pAmHnL9iJAi
ulbR84vJzGVC5bl41aJCjHT0oIDuNY8lQQHPCm999ZmqJlRmh/mQu+ARdwmKm/4C
wx6asYqVNlMR71k+01fE1QQCAEidyplwM9KhMjYlcyLzPJAjQJ1OsQwdd6IxnE9h
aPHmjtlgthA+3MtqOuMTDx2SV5O0sW5J+R003szghqEzAfPFW+TrIEhcAnVmV87U
WscnVynUvbeGtnEkyB7cQLttKzxqf4+9rmyrPEo+hexAyZlH4IqqXwQN9nDcLg9P
ibWbDNQSNnIyR5Vi/PEZFCarSWUWFh2l3dQ2h/UF7TU9YH8ERiXxEvw9+6X4kROk
frpFEuXfcLj5Bmc0HRkGbLB+p3t4vIUjqNzkFRKu2hJ3UCfGChVOD/avqvNHZ2tf
dzHdC9onsZum1Fpk9Rl6ydYJ6q6OWYsQcDCZCe9n5tfy69+aj5mTsFzwKUajOIZC
c7CO7H2RFh12t/f/7uioIaSc7Rt0w/Sgx8djEr7iFpTyZqybvy3GE/Z2Qsu91bE2
Op6jQFhW96w0rh4knIbXkQQZ5JOQU6B43v0Mll/lJGAMGKxvEs/JOHAFIXLORpgg
SujdNspjvN8nAPWAo/I2wItPiKPckyVoP0vpQgIzKFwcntqfhfk6UEehTxN9w3Ej
TObArSPhE64xisXMHnYaC4jdi2fb+o92TOQA0Mdu/YHFqv/gdwdzV119qnyYBOmq
iggKsDW5kJrvT1aC+WF60o9l5HOrYKzCIBq+SuUIDnpoE/m+mM4lbQxhMX+Vd6Yr
Rd3GOgTy3Sxn3BuM4DxMa3yOOPiVjBWyAwFk1lz/9+BazuuSfp/uk39O3xJMGeH/
4T5oLQ2+V522f6+k+PYilhAsKNobWRufzuvZFvjps0QtMv5i1vzaMuRblvel8VMU
UXvFQ0Dw6c9VlmFpYmjbkLBnAGEqHihQf7w0pLxgOBWrWr6ZB5wMZ9lT2rmUShg5
ieKJUWBcv1KXh2MulVqPrUGt6qfBWLSWv8dVzTh9X20yczB/q+c+WX2RAXb4hUf1
yXfSAsdbhPuCy5xEV+SrTWFdOY0Te8/1qYf8kOR3J1HhWrPO59N3w3E0QbbZXPX6
xFCGJD9JBPgac/f6qwTkc0D8C4lnfHJrCjvq5VdEYLFsgpT0xwyrJn/ZdmlLdFdz
sE7ot1EIImKZu9M1EpNsbDVoeO/3M0xgEBExc3k1tDOCR3s5oMiv+dMvA1d4grq4
GAEj++ihEZb2bnk6zUr+JyqLFljCGWbIv1AqeHE/0rbLSQKJuF9kbKoEr10VwzFc
wEedf4heI17RdHZLd+DQBu8P8xjj5lWArKAFTMZIgL7kjtuOBpYSUlXwoUCWassD
YsDM7XmstViRGPbwgtdvTZop0ugyT3Y8b53qf0C7aYd66LMubHD3quB+Z3P6JgaH
yfXmp0Gm6CeJ3QwRZ940es9wp7IudBoxppj08utCuPCE7UDMW5hFtkV31RtqU7Zz
DwYiUGTsXZNVcD+e6H3yhJ2E5DdAVjLY3aRhWFjrsIsT+QW2KehV7/vyPEFfjEvt
0fKquPbASLwnZWYSvyRE+I0CXDljun2FKdtKEC1q/F5jnORSCJfDj3XjAakQPhIU
GmvoykeCmuiouqdklxFpKM6lkEOCYWki9h5XHLFF0YYwEnNA+/1cgvn1qHp7Szr0
Y+k1DWAFr0FoPocpq3OjxtStGerC1taac2BSfg5K+pJYaJuNLBVUTj+21u2L2pqy
N5JjNObvMjcgnzAQLmXnLjuL0Rc6n1/GGdh3g7Hl40jpsYco2x5NHTHyZui61vQE
bf0ftHAvI2FNbIQLel1df97NmrE9ERgbONFbXTaYrw58bkQmLIqxilw6EMPixcHa
VhpWdFX7f1SOH0llY0vuN+X5Z61XBFN1AHIRQw4L+ya7ivI4CC66B2mXPH3RHlya
uPDii1/OAevhNO2Ib6Qo+DCh/KWqj+ELrzY5NU0MTSQ2m9/kcz+tUvqSVU6dVUo4
g5DBPnIbSwt7accHeHANn0aNgwxAq3AgMS4paz9VHiku8YGuTrOdm2/iPr+1Z8XJ
FbZDvzplvE9crSYc4+nETyP6Osgay0wL55RKPtaqclLNnZprvXXoquhSJUKDFD+m
CBzKXygsr51Bx3MiJp267kau1l3pjJLbDzzgSQEZ2f61RVffx7X/nsn7XwE6R1XE
eO+ERY8cdpQXC/Z7Yr8iy25EHaRKEaPWImLirIKeO7ulXSHM53I7S7HB3AP89I3D
DhSr0U2vjN8sr0rkBWWzZlMSEopXvhgprt+NzNdxmwtUU+Athoc7kElc5uP0aL6+
3/SSTTgLXCPJE+sjaZJhPahAlWB3H/mXDXbtOPIps3uwUQaTAF8xBXMfNTQlerTy
Q5bj0HJgqGixbyoBDAfUgyQPyufF9s32/IdHXRfqlKZbhH6z0HD4H2+We/i7ke7+
yODdvdAYL49aZWnF5ACwRaFiHZPtF0VH/z9E0RRUYSwWvVjEB7HqgwtX5NwvTRK4
/hIJay0VlnkAuVuQ3fx+ZanbTND867pDgc/Ozyv4HA51mndwd42+i8BOraE9F/Fx
DxDlR7h6mdN9ncV1+Z+zVovaWvku7i/WICQfIMDgbzyTp8fGtEbvw4F07v3kLhF8
lELa73TTGrVLNYYPykf9MZkD/H5/tzXojGt4kFkZ8r3FOt7Hdy/Ehw585oOZKDmc
xIOkQGHVciEhNgyoqJbX6VWIILYGqjyeTGJHpk4naEPFcLylAQP1q/o12GqLwffm
xvHHLQfzjsJnvah/mA8TNgaaxSBd8z7XkbBE3eFKlgfwjUCphhW1h2FK6tDmNXBj
hKOOCusszpkiyrkOhpodzUwVtWLsrmPT7TcuODZfS2/O2cl1aHDGwrqj6xk22BOe
fmHuEildqr3w78W53OOfEcyOjJe8WLtUuMlat6MVk7iRp3bIhxE1IX8ubLjf8bKi
TtZSW5jyIcLqbfWVTQpecRWIKwO+MdPVKchjamDBPUJ71+jNikEh6dAUUnRKuWrU
c/ahjHv27+S8Mnojl15JB/Btxfl+3kSmJI663Gblgx7YLsfRpaOUMGroFfu7JjF2
K3WCOqpuASYZtX9UlyXIsfd947C4cHK9Xe4LiscHaifzFOKzpCDycqU/ApEFmuqO
QuDH5SPStGs6mTyx/PQIcJkrJswkAgO+ct69bGU4VHopAoKnYI0qO1jSu+u1gVm/
KpsJKJjuk/wM6HLbG5JFGm+fcLRoeRaHUJjTYyNcFympfAYejrL/E8t0ulzT1Y6v
HBfdJ6uuR9ztqfBNtit4LfYLM6W+XZ5LZKF3SQz21jnr/0fVvCM/d/c2vhNnYSSB
MbtRH4jiYaAfH8py3GnUiU6SOkhVpn2ndZY8w1646oMOfYWCUdTxVF1O1vxiRnCJ
MSLRHBLVyTW+dFOA4INeFGR3PwsG7GS4opEcKv0KaBkM5U9ebQiSddGDZEjNvyFO
9CcqWFgwUGQ05qUhmFT8KbZpFIgv+rcxJ0+Bt4RRZT/FIM7b6Ka/Wi3T357XJJDA
dM6OyrIl/TQnhXOvDu0ZI2/JyrvhOVL7GrVqOBbUv8J7WhaNu/R45maExI44Anms
gHBIy/jh4a8WzeQTcG+yrVn/5q8Mli8Naf6hlk1lbS1HuV6OtSvGdNzivtvo9/hQ
N7p/zKO/8fPhccjTMBAC1r4Pm61pO15bStXhTTNr3o6jZbZE9o2HLYK0ovOwikIz
xnx8AmCtBRHCi4nCdbjExL6DofoDqG/G6DSGeE15xppp8VrTwb9PMQWpj48qdlx+
H1V7HUbb7qSpiH6/HePOsXcHzhV3i7PrssVsus21MqVj8flVf+rBhQpET3WulqOS
NSXtll37yE1oDkC9zBXIPA==
`protect end_protected