`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 25648 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/9huKRhRMtvnNqb3Z+UU7TahEoHV+T8U3P3ufru7l1O
3DlgtZzb9QxCbOjthp9+wDkjygH0eUfDrEl1ovhZG61GnRbgBekzs4BHMJR0xyyP
psNcbeCfolseU4wLZjiW2TsW8MTPFUaRrDjsRSJLWp9aDqCqFX46PsUESkMz+XJJ
j+71aWMDA5LPB296xFbEuEoiarHnYY+P7cjvg34qmszkdKrZWXoUJcPCdlfRPAZR
BMJElH9lJ9zcmPjDa2gYfBKKs6tRJ2k228Ro9K8BPrleyFDWSXsg773YHMwk0XFn
KbaEO8S7mwpbu6h7ZMapJFh9J27VsU3mCNIZQ6jzdBUOEV9n4swQpavITt+f9HQc
bq/brs5LNUMeQaU9dcQ7Oenyt2GVJfI80CR53MJMp4ZFNlpVh4zyM7xVcW8mFwCG
V+AfYDeXr2jexPaqPptWvGrxhBIQVy+VKAIV0E3VWio251P4Y+V5i7j2jloCk4GD
i4OOmrOvthFTprVXbP1M/APy6huyXiH8ODp2Ex5DsyjHG2UPEJT+u1GielyZK5O0
tlfbyVSo0PNYuUWg3Hwf5eEKIMHxD00S/fZIrE0jchpvZS0F9ouxeD5UjTMwaNBn
gdCTdA4mMrl9JfswQDP8LVWR35jq5aTOTOXpjtYAiYv8VJ2+UU6yKpLAEFrRL5RR
cFt2CEQ9Dgy2C/3U2uzw7LRbwF/eP/S2STRxbi++MCvf6xodLWULmqQY9O3OS5yT
CnXD1jcRB9GwrjznRPJVijqGu6qIDSKLuCe9VPvnPpzZlQJcQmomqSw1lsnc5ZtF
KP+ulvtrByWt4xPrAiV35H7vlKY9wlxQhRJCbNsBepIKqrz2JcbqGuPsyD3qxQRC
nVozxDyKXMZA9qN9rQ74O03GjJYov+4IWHiEfO/sKnpUSk0aZZKiGcmB3xyhAnDS
8TZyvnfXFdDW5xHQ9OG10zXe8+hNSMxWwyI+ip5NdJg9oOA7KDUSFVO/U8stTsHG
bdu/iOuWV4bHxnY8ccYSQg6MSvlHx7Z91x31unr/ndEQ7Ixbbzn4Z2vg4H0+3PBP
235BZHZXrndt6qph/oC9R2V5Kj80+y0q/rthJ1FPmg9kWi1waO58b96OYhS3d0Cj
tgP090OD2gROHvk+pR3oparQiiD2SR+RqjUvwT6Vl/UhTXIOXkH2rGWpRYaiRTKF
8ExtQgDivYKDxVA1/ozrO/cMIaRN4RsEGg7QLaxzWG7/9e/NmB+E+uujxrRymksS
JP0xUYIEw1E8cGPGF7RUFzO6ORI+EBaVK4e/2A8Dp48rL1KdNB5tNpMO1VDEyx6g
Ea3u1VtzL+JwrcHtExuCQBk5xQz5MsyCEh0j7vtX8KWxgXamgerCIvUGSFWNfxcV
NCwnzcXTo5sDIMr4s4j+WTn5VKId+nSuQueVsuXRxqZlfwi++zijK/nqX1DuZOtU
8qdE0Brs+TzfaUNMPdMHwMTmUdhNwJB+ottatX3gIhNiJ/2oQsPWLvuV00cydHBp
at5vo1PnZFnC3Bd3LI7SPWscIvfLIV8wvwwOfHVkWe3BFIyodctFKmPts7ypg9j+
+h+AxK0TKsw+g6I6WmAA+EYxlazxXe4qYCUJg7R5aIit6POem1AANyl5b0CwGhTN
1iXkjwwgwBMKaKg+zgva9mjp9t05d52In3qnjxbcE/AHpIpDBsl+HOti0QmpwHQ4
4AGz1zk7b+4X08Cktuu4TNsx0T8iwicbzOp4xdARm2yyFp6VYlzXQDiZ4Oun1Aja
/Vz8HrUlrnPX6K9I2lFX7JpNhTMqEpJGMVbeL/7xDKszJ1pmp01BmER8zNIEEs/n
J9wfLa3NsVKAAQLV3yWRrueGsPD6YSGtnTcif1KmpoyddRJ0TEELm12e8bzYjDmW
4zm3T3boBmqmdJo4gTyAedTS0qwdJglsO/T6L2OQ1qmohPT5xqyAAV9FLcHyXz31
9BCTS+Azg/+ZbziEuiyRc7MTfbnmX2jAJjBESK+GwRBV7odUFDUdNfl0uHC62Cf/
QJNn8Adh+euM1cd6yE8GSvmMuUWOApsHc0T/hjp8ONnHW1X4/LRgdrMBktGo31yp
d8YM/gDd/GYhuFi05+lpRf6/0gJgl8UlOfXyY1aUYnPbzt5gp4cwvECVs2Vw48Jf
eAx5/ybKxRvicYY0yP6QkVxv5MvP/SsmLCHfkj2HB+8tj8AO1tAWE/B/HmxuSsUj
T3Igt3Oc+MQ9nOg7HG0vVMVYx9C3gCY3Qd3qAyJYHWiOGLs2pS1oyhZo0Q6MvBN+
8d078OlrDgsGFfdyCGyS3xdHI+ldtVNGA1n+R59IwcwlvKrY9VaVKpg8NYJlxAHl
juUc61YavtCqu+7R6PiruIeZ9TG0cH9Tqlr7H47yDTECN2b32NlkbGY1tVo8ozKy
H1ylu6hdhf6YHlbVADP24joEIUxfgAKWsyS3YoU2Nl+cPP383tjQbGTre7Cagv5X
W2pF2lu72mHS7XtK0KIZFtuLlJtS9WIFEZyfs0mNzJ+w/2ai3xOSU8pXOCphTOQS
hcUJfI17OozmxCQei5T4BPU/YTYnQ87OjTCy4jK1EOezYRG099p81UxYNKhr1Mf4
SBtqVs0gSYmGBst0GQiMoJ06PUNY3TPhwEWCdinFe/5uRuqyL+CRqt1gUvP1rvfF
jKQIKs5NJzU1xFgUMRB66kYMfrQ/EJaZcjIHdMFO2xJwMZDqQsWw6U3+36ldnrdV
U4m4Zw+XKgEA3lYPUEVn8kyrFSm7dA1pqakFVSLV8aHikwdjpsS4zMVjlfKPvJjO
XUdfS4AocLVITo0xz0EPFT9uryztIMtFYE1NMP4Wt9TUBgzx3/Z4crZz1U59M5k9
M29KhYKC523BC8z+gXeUCq8awlylkg+na/TZSkeNn5pZai+2glAnrvJVpoZ3jPds
ieN8lJs+GTRdjO0EL1n8j/JPAz7Nv8YICgooKGA/tFC0S2zf1u9YDGgkAQDFdqI9
h+0DbWGdbCoSCpQY7reBVnQXGzKqwaqHAX9HFCzx8wI0fM9nBL1m9dLk44nEoa6O
3vBlxCGIXLNCUj/JEayK772+LiSley9FeywpDQL5Ls+Bn5ixdTOkdKfLv3Ot61Kj
KU1xJFKe3q1DVjVxAAwUuICu8eEe7hh/AbxtazAoz+KBy7F4j0B2KlqQZXWhEK2D
W/xYIB8zj+R34ArrCwITQRd/E0y+6eSoYmfga2O1h+Ob1a+gVSJaqEjgtI78d0Pk
j4MQSqLg4oW54naF3nq766P6SDcrCvKLofp0nR8F50JUyfPkfmVzLzbRR2+TOWNR
6r2pqNpConfX4QGWM8rKUwVDO2PprZYQiFbIcWFIkKmA2TJHIYY2hPN8eOE0cuVF
PalEO+a9ptWTGZ4tXUAi3pbNXnlABdv/aBW/50o89jvhsJ3tyKhwNQUM+MHDMGJH
nNCATQI+TQ2IOdTwQGV+jwO5vdm5RkYFO82rpkZeVzXDMyZer41tBRsy37E+H1dL
6KUL/1+NcG0kZlFbBxKrfjsCc35SENSOvQ2CnekNCexVQK1DLeaqKojdw77ao1Bv
382pZcpSS+LKGqcgTQhEi450fRUsplTNlHnL9DBUbtFq69NWnc2ZeIp+KlOT8zFm
pnRY7BtnaF9okEzHkxgtwLI8yoTnc30mLZ4cQJXChpmAWewxwNLuSA35j9pJrBsd
t7wuRd8IoEEHd5qjpf3ZQw0YDSMFb2nkFDUCXN+7UFf7DivHbffX6tpPPkBPKELc
S0o7YJQlPL2Lmeq4hiqtOIjC20D9kdJ7yUMA0IQVhC+76NmI8aN72U3A/ZB+GmUD
5EkWIdMwmAbjaz4L/zy7y2kZKHeppu6x4UH/GEar6LgEPqtFotyONbABaK4SkEPy
S+wsvUMIP8h/Y5nD5PMNpt8IMjjRf850OPiVE5EnZeduTLrPvdmM6uSNkNyq0b2/
tEZq8bFfUWRnsGegOOkFtocORYzP8kQW8GiVWEqzqtW7Xmqr11RijimBlpV+0W5A
LfxmaEr0lzrJE/L2/5qrNPzJFUYbSreaTSJu1aO62h1luJh+VMSA56QUukyuALq2
yoNex+p2b+CWI1OEANDr1lTgRCtt5M+maBt1WlLvmdoB0/sorWigmJXWUeZkjCae
2tQtztB7LfSjrZ8IENTDmoJL8lT+PKuNuWxakWAJ/SLtcRRaABQJ39rhB7gu1MP8
3hZ2vjIqJFW9nzk/QRNsZVRPuqW9PucdYOKCe6YDYO5S15+6trXaV535gSQOmOo/
dyiduUegecgJMEYhtmNKohT19mExUQIT72ehJcoBIAcVsdCjehuFF21MpCvmOakf
LjWFngiAbYzZlMJ+oiOwsjngM/mesObDiVj7WYwqRo/WwUs+CrgJCL3n4B3uy+WW
H7rN2hooYgJBkcR1y4TeQEynshiA6OXqwEi0HjOFx5bFJ1EqfVYfS3a01KcRgw4D
j0rai4VRO+rsjGE6PsSqv7az16sGOrbOG0DmqCXhDnv6mklo997kwUmdP/uWArP2
X7hUVmiCCVOhWCFwbkQRap+hvWYiCuBNksNrk850G08cI1S5hZKkCKlJxDk0Aj4E
GL6XUOomfnvgKYmUAnR90H0HL/UIJeeuIy9bKec1TX64t1ePZafCVOrRkXMfVJWE
w17IeoLwabKWutQQ5+VIHaVus2JPC7BrgdWSdh3759+krCFvJkU97CM6enOUM4eI
VkxvioXJ2wwVOPQiVmVdx5LPoQJ3uOcD2S9hmPFtPo2AX2kD1LVcl9ZMXQqWyWho
EYsLXGchqoRfmMHITD2EUefQOMl0pydwtMhcfM5ZwJDrkGIBXsxzrBbkZRRH4Csq
dCF8K7LceJx4tvzlp3XsgCWijEWWLqtWaUpBcNzjtSRQrDOjmwENxtDTwQ00K/Ey
GMPjt+tiFGI6Kc+z7fJiwGyXq1dbi7E6YvZc0GzKqleCTpvy4HHhbDa4RLzTCBKN
huAZjp3g5QjjQCfISAk2z1Efk5zFYg9ooacO1tfm/l1jI/7AerN699h1QtJt4EgS
KPlOvhGA9xqNKjsp/+DdJ43Vpy5b/Bp5uXgbjywn5W5S3UjNWdjSwt/hpKWMi6Na
q1an6t7Z1oeki/MUkfF4yQBAIeactwq8lm6s/gjysL2B1b8pIkgeFiiz526kFUfM
jHXYoImd1MGtLO+fjQG+yyTE6B13DaVFb+jTFaWgdxctT1sgMzt6umaZ49FjPDSs
Qe9ahm2tpB3X89mAkY4ix6zb1Wd53xFVL9lCsjYe+2g/DLY/llqnyIqncqQ54Fuz
l2vy0jJvzRwaPvIcyDtLB4EZNlLZId8IysKDvjzTckSw6bcl1T3N/4oEqkRo/bp7
3HlCTd0YJJVxWxKnYfkSTe113NWn8W5cV/7fAIsyqdbV+0X1CTFyf4e1OY+SD0Vf
rTIuek4AEMRVZVITehtkM2YfVY1XYJ8RbNvcbGX9nh9wW90/JCsgBPtNZWFjaHwS
25z/sHR+hKjKFn1xNx36un5iRDOd/P43EAs4EkoCdtuRBHsflXBxpSzDAWybwwGg
+eYEQ9Veq7jpOfcs5FycCK6gSS7KLVv7/j26Ny7QPCaHCtGq/O2VFALkDmnOmFza
rEuyuddFOnJ+rvadA1nGyzliwNU0LuAXmiloh6nwR3oQzAfQnzzdFLq0mIx3DQQB
X59xWvRT0HIw9u3Cez7Av3eK9+WbgShc+igYIcDJ/f7Y7xdZi8arQaZJ9L/G2KEz
dgjFfWr5VWCd/5koZgtg54hqs+fHxe0Mnc6DT4EgQJS7GtE2zFZ+35Bqd7O2Yv81
KcmDCaNKNndgCWmz05c+++43tdZfEXapt7rOZ5pKojiERfNtfAjhzhVYjsqhQ52p
jsouowJ2djqGY41p87GpZqCOSl/uoZMMnaZIJXyzpcxlXFl/6Dus5uIqiPrZK74y
IxYKy9IxSYKT+j7P1E7cqY9KkPX6N2l9GqKmBiR3NW7v87jpvIf0U0XyDkN88hYl
6ekiCWFF42X2wdocWQaJ1D6gcZ6P1RM1gm/LkGEKBkb4QdXuD4KZwm+v0wFq/mgG
JevqDyGBN7VDuBBf63SVgrVISBmaRejZ/nOEQEcUL8rV7QvzAwmwu2d0M+/sD8PT
LxcDk8ebW17YB9zuBGDnGczT7+qhkl20zSjh5zbB4JweykjocEvmoKAWOHnYl+tM
XWKvBNec3RCITRm6kXZMstmB/PSddZB0NrpNv8CFLXtg2tkq/MPIa9ezSW7/Ny9W
RTkuePLRC6BAYcsQ1Z0M5XRIYBYDNCmLrJsk5m6RyZIWdje9Fx7yy+ltxK2ZKlyt
otdX9VHyA7gVvvWCu11TKqhJsyQpXfRXfNTsAR1nnoSmrfnlpMxhEShBCqfBRORy
Mn6oTAXaw0jYADdiHiUr+59BsSZcWC/SUQ1yYbwfVTQkKpahh0NGaztLqVB44gqg
OoDE9oVFECJ4T47ZFihGVQ7ag3AkfmC0VeN1OQQqasonkclp7tHuKaSz+7dPNLBI
cqg8yMS9EvRE4dnGLCzyT6VL1M1fG+mrxWFNCf+qiazOaGVSxkjvGGXee4Fp2j4L
16q9rnWBB71X2KJbWep/bmewW8bueh7FsKDlF5v/CTZs/PEtwZwglN4JSD3xyNj0
y1OLT4z6SCe1MBYjJwX8MFtpANjz2hT9sqU1x8k/Sow9+LbQF40ksQOcZ8FjWpG+
7XYaVPZbfvoUBUZYsoyi4gq+dpu/YbUxTm+cda73F949MDpAdp8mOMEdKXQIE3GS
OJf+fqLZVQuVXnxapN2zmnAztX6fDu1UB/dqx6lsvhDUh5ts9vep5QPstplMf+/l
NheXrj5X5j6yJfnV6e3roCeDpPl4MiYtZF7kR+BNIXdXYG+lqme0MwHs6y/Y4x7Y
v0G2nB7QlBOeJAppsXXHM7jeiRWqRdJdodtANauzyyc/hqxvVEM6Fz6wBIAZFovE
mOheiTtnM7vvsIDqL/JoAoW3dHavLFpR4Bp4dG9AZWgogxR8SWnMd5bVyAwhY0P/
qT/h/NMmR+73kEwNm3hHWipTlfagGb9sG+wB7rlgHo9RSE4qzBul6ihE85Ej1hqN
wBWdmbg+juHSAUgJeDNJWYmYzIXzHPpDZU2hxi43CHlyHXJVOPLfP+RVbAg1l8PE
FCKg8YcCklajDg3Cb2zHLk0Yy0i/MJ7scT7RpYFDK+NPNZQLDGxqSR50Pn1821j1
5twuCGPEegGHsprOdNwcqxQpNBToHpPqILeU17dltpuxd+5MpuEhsqCcV6+yjAUx
mEIOofcxhmF8xr+ewwKXolOvHvcr5wGC7KIqVhqaMOQFzmcgArj6NcjlXKqJpWWR
vWoBJeIEblKgCEfwI4X5ZQh4oWZQNPJ/Qtoq/0/zMZ87A2iiwrsVbYpAOJB2JQxD
oMVi6fUbQmgn+1shfUgBB5QTJ5RjQxGwrO4nS9osnHzTsqE9zjGSj02ZWI0sSOyI
D+rNz1Z0IO+It+/3PUXz+BpST13uZ53+R7fmTSvxumfOp6z+9OklL06VckTHWhdk
UYf6SMvo3xlvhyP/kXiBuEsBAbXeDVZrbTX+hNk+dmaNwa5bjyWjzRQXRW8B4Ppj
HPOyBPEz8w3+dHTi+/EHPBP/r0mGEBLvIAqa+y/ph2ovC3XVqLq/Z0BpTqRWmnbL
bBt0Zz27QeaWKKzXGHckYJEOgynlAj98E4nNdn8KQ/3QdRqWjIXbphEoBt5OAJ9C
VQPMeNnsv3vvFCPPsVDOiPadl3MlfdEWTIa+rMRZwHTxgmW1HwSQKjrhe+f+0KKL
6U8WeUHBBt9hyUNK7UnlZDaZG79lloO0w8YYbGwvGFDhfBQGBWgTkWKUplhEmmkE
I1Wo1+siXG5eWt/jUMbAoGE450ltggeSA4mq9LbxjuS0biS8+SK6rTbKh3KDF9os
T/eRlBP8fwE+jwb10DNYgOQABdQewNuRVFy9wjiOGx8pbHmHbZ4wua6D5Gy7s4NV
cfMTbJNO9x9AoWJIoZtOGabTJIezAa8DD3OMjdEU+XhJw9zVDEqQy4k85lBUUK1z
jqMbe+abruY9L278CMVh/rzPun8Icu1HAjEAImajOsNMmKb2yStQIDlLnc6A6s+D
v0pAd8QWoWJB0cc0nkMKt7mLIetA2P+DYi74c8hD2zMQp2+BkjCnB3zZZFwBzSUE
yHEnrI+y7SVkS1C+lhwiJ9XIhQru7QLdVKEUxma2Xh0p9Go1VfF51RpYTa2DkafP
ew/fLXDcuIo87ppshBMWRGeyKN8eAY0EzsEEfuaqxrTzIivXYVCtQ+drvh0pNl5N
Rgyx+T4k7NIAGIR7dNKvjOc1lR30ifkxA4+z867MsVgvKWBxCKE8jBHpYAWLtjAS
3UsdYNH9fK/MqjHtzZp5hKrfbibk4ea6yZtRLfsQBzhZ7A8X69dIKAvw6QXmZQcR
WjNvbGrW+nzfxdDlAEqd0DuFtqnji68MwCI2BUKb0c0ucwz231p57qgpygHv07Ba
KX6BeA7xMc37elufim2jSln6DyUKeIjr74JdrVUF4A9zG3j3P2f5MFdEvygWhUeB
7s7CnwOrapZwSj97KlgxeFjGuq89fCp/8UT9VGA6AiWeJi0dPpDCDrdrAu8Cx/YV
ziO456Hb7Mp6jX+CoGoj0TNNjcxMSAhOAKLD3Ojh79nXunSLvjuW4UMBMXQ105Cw
PIYgLRewBYXHeFaj3VH4d5tLmU+J2hfkx1yo57mo+JaXHNWaOhuWs9AGSsBkRZo5
baDVqrczPCQ1xhTeG30qwNPt/Hy8AxvyrxyofUx1I+Umaqwdp5Uc1TTJT1u0Ndu5
wUtAcoiXKt9Sm0BxGOv9KmZLFEpRVEGqfmHieA+6CFbsy010swrmZ59eYNUbGwzS
p5qnlUIqSDEEGWYbpKBWrhi83mNmK/CvupwELA9GykVJuGI7yOTQ5Mgx5JwG20/F
s0bZZ0218ofZd8wSUBFtn+6oiZEJ3RGjp+r4qeCM5NH5FzhpgdCgUeLH8Gfhcdx2
CkKRTeBkbTMjt/cQe2lnfckdjYsJaQCO0mipZ7ek3kwTBCcmqaEaYyOh7uNLHuID
yHuP/jlRwXomzmt8JYch2hCcLiwc6QliGaDm/XTGzfebcKmHU30y05kKVa2fgL/6
0ekMv+X/H7UCaFWlUAU+wm+TSBb5rzL4nGxesL9YN8IrpJHKDXqZDwM61N5feZH2
UJfFVEQ4jdyM8ejVgzvv50QjvKoYo3XF1wqiD6ErGSSlL26KMi93HeOAaAGyaLIS
fThYB7awZ7AX7dBRztZ4zVOY9Zm2qGfQGMTDjd8/s+aIpIzsqird5c2fdT48q5+w
0TKWqeqgTLw0UiMSlx2Qhe/dN6VK9cijyhW68r5MxzYLdVQpPsrhnc5prbkZWV//
h5Vm13yUcnL9g+W0RQ4XgVO+eHQVXBddNcAdkjFNKv+jAwkONjLXq9z6C4TpgF88
AJYOZTi/nT4bgsRwZ6z0rG/bnxxMy/W0XszXgLTl4eVIJMyDShMOWFt3K3A73UtN
YI7aMmKB1+C6accdRqjUSBxKBuBchg37f2II4WTPR5H671LZJupdOnrOAs1v1nDF
ghQky4PnLbkcsdDOGLGC1OQl/1IcEwK6ST+psr7xoi3g7CjAs8zlG6YvbQk2Cnss
bXCskXKqekaOgdgiNfHO4Xj5FvW/uujrCzAeOZcM1Y6FfXBj+deGZIV0meekjhs6
RM4qbp6Kx8PYf85Hdj4Jp0lXQc+ZioaLrDFqJzbXTwWA6HnISwYXQNIkWjSpETwB
pDtw5WA8U5JdCJIE9jiRIOqiJ5NjqXyu/8/lS5RhAadgVtVlUlke9V6uwxLlLCLy
80LKe+ZSx5r3JBXs9NkArizyT26UtV+MzY7PeemPKRsNclU3Yw7rUmArfCfqY3UP
3acT0fn4pWta5dS6m9CopKZxwC+jNOcbLA2F7z+ORFkikMc5s1gr3S32MjhSwGUL
6k7t1ISP9HdQ72lDwZFueziQWFGc1sCW47GpEJsxoku7Q0we6scdBmSF6LTzt7FH
hs8ZgBXBCXKTcPHXpd8oWDuIsTNDpRwYG/ND6j+25YvYfxszo0sAtIx1w4KsmO28
y5E8YVfuaefFA9Du6KMIT6osvXH7i+wwx5zJn7FtoWVgQ+Bo8qZZ7Ey7SNRgOFYJ
nSTx55ZjiCEs8CpNQT4bxx+Vr5IAvShQtYlYk4vagP6nPjaVHxeXKzOccvi/ZmLO
pDZGS+Qf0VPl3g/0NPN2UtRicoUvctney0FYlPbCLydOc8hncdO8nmL3MzlgaJZM
nOVV+lSDSrQ7SXbiovlf8MPmBxNPVljIg/UZfxIUeNgKFuRUZ/eLBiWwj5MLNwpa
rciyUgiLsCY+T5TaYz/Sps4vXJ2hseMXgdiLhHy2Z6cofW4EC8z/RMlD3IBvdRUC
4+BN4pebKHy8+VgcRU80A3DmcRDfbIlE3brytc5QckD29GQ1qnFsw5Gvo9X8Usu4
YYB51sqUcgAFju6MCB9aYFTQ1gL3/OtQUOkAcnW+HmKketClesGvADE66l1fT35R
PH+pdqMU4m3sEBXMvmA/bW3lQ+uz4Ocp2EAy0xw0bj6gAQpT4iLLk80NWL6Jb9bN
EOfYsZDPXCaxQ3FZttLZlCRC+a3X3pJdP28Wtt4vX1fo+271vAHLOGkyhrv1YRMn
WG9bWbh2K6Zb8evlrziH5mKJCPvEgNX3BT6AB56cbIdx2KT+8SdTexfA2AR1z3zy
1aEqOomqbJD4P2mmqyS/WJqAJVeKzwO3L7dLFFDl5m4Unl4ZzJ4tKshyN9hbVV7q
/jkZPkT7p5rEV7nl9cS0MWhpRt7jan2ha016MYaTALLkLiVBh9zmh0CS/faAm240
8S4CGMOV5UFuT8CPOBhNfxZ+RWutecb0tXDI2lmz0bw6F/Ny6PymGiZocLChCwKa
TBu3m3oFKitjnowiXHrz2D7aziz9yy4p3cvUwtbko5aav8dzON0yF8+NIiHlse+g
nlGcAU1HzoY+m1HJ6rJSD6dWP0vglID/+VxNHmCiZasf/L1sg0Na7YdVSICckIX+
aJSRWQXpRnQP344MXJosC94Wf/P+xzVDBsDmikKq7zjTbB4+WuVYAzPiBdxdpqQK
g4/C1xgKG8EuQo7qR2XOkAX+DvnU7/YGRptfmEfQe5wmlDA0oXOa7+evdMS4aU4j
csrDfUSJuscyJllUc9/GRbSgCKbQJrXVaUx9fU9jbt5hD+FFA3KwMNGL5kAFmrGG
GPVt0hJ9EF7GchcFMZRtC8wYMGDaB4z7Oa3FGy4HWJf4bneqrumH/sZ/T9+lBbmV
4A+PRQWSYQR1cnK0efEDvxwPQSlv/JRRwz3j90Vo3s8xKTmcSLENeCwzSK+5fJdi
OteRn0ssQ+GgRMcKBdAlQE04uRJUZ04Kp3Vxy4adN0hDLyHbvla4NTmW2fZ5IBWX
VO1A9XdgnE8euwxZX1wKuh5hal7R7CgeZWCce+mrp0dMMxR1PxYvgvnh+QhfdyrO
tTNShjcjUKMMHfvPoYNhsXh44nDJyGsOwLx72KNOkZ9R/e49+bUZd8/gecaWMz30
MqLfkXvfA9NIqrcej6VQFpUVLl6ddXePLcNSJyxZk9gNz6LA0oNCnVGvh01tHUoO
qP88vIA0fGK5Zk0aVPN511QG6/O0z9Cg95e68j8Z802NZ6HwwDKzBd5fTxGX21yX
DxNiEYM082LSTTsgZgg9ROOHrFgKpJZTtcsuZKerCz7hgXMP96dUc9pYWSCtU5OH
/+sx9cmDXlYi5Nk5tsfduYm1rQ0uzNuH24kZp1WUvHg+nBdxEWhpEbhHEx91v9NE
PLM0gdFLugxV8wVYvNFQEcaEZkJlrZkvW2Sw6JxGFGvPuE+AEX29N3u79Y1S2czq
TN780Y8WPPxFGhVMEiutGTGyfJNYCqi7od1bgLeCJoTvPo3Bj4E27LISRI16MfM6
Awx5MDyVDpQoqQFeqTXZBJ6iOi8qeZlXRTMCgmkGlPFhcS7mhlwSmRpYpsx5MqV1
khHcuK4w49wTpwCQsIBgSMSBFe5YUP5HvqBLzTFoCYOLUXHgoFhMBmyUGnttJlbk
spOKmwE+LJYc02auW0SlijEHnliBL7y3/erJqid+u2EBhKrTeYe59IPNzdpbUa8a
uOjWcnKdi4uQ8c3fzmoQCqvEwzHQaE88gXZhWXarwjEdTyU44AD1H4jA8o4ehA75
CHODETfo1Jq9Z+LFVdihLc0c+ghV6KEABlcD2xP2+p2i9ltMOIcAgED73WASaMs2
uN485WYWnYjr30aBcsnaMODN2UgFpq+rJWD+5vZRzQ7IERLy/r6elUunYxviNBvt
4eq4KQeg+/HJDsYt1HDHXxhiNJS2HWdwci73ChsirASCcrROBwfvAqRitbAYpXbp
Hg3GnvV6s7Rus8X6ggfgtCTTSlgkFOBmsBJ4DzfEOko391UhSgl2EMgxq5WdRdJL
KnDyrs15r+HGUZkxmtVm9iHiiRT/rDYfiu4R6YbT+uKPdSqvcOU9moD776MiwIJJ
7Oq+0BFFJ5135ToKPOPGVmzeJzpoZ4Q5UyiTtM3t3JBfb+0WaVUjl28eDNqwP06B
CgRR2fPmFJpD5XkX2woWDCu/Cma83hlmSlGS/SDleK1VzMImgjGYXqp+uNkypiVP
16j7yO9vcHSKHPLqiARPaK2qgjAHXlOmf1cvD7gde/nTZMid+yMITNeOJb4JN0Iq
Jkah0fdKSz9jgEYDY8YL1neOnL4QKYkggqwlSbAIAxyRzmsx7Ho81GclzaijOKrW
8XQjzWak2XxVrB9O8qcAqsbWA5uNVXd2ksfjIZNNwrDXq0PQcQP0J3UZVdNAM+GH
faqFJKeTk5wDcwsFv/WwYsNOyLAF7rW0AahExFF+0YlIMlh4PVYzW4vTwFTVnN5S
IRtqcxKG0I9xsbMiAZbofakE7++OviA620RGWTU8v9MeModQCSIu3vN4Xd4HcNCR
uxlgRR2k49k0yD6mPcIAHuRlMp65vl2XNWfHLcxU7261wdMBv5Yu35ii07gnPu3E
518hIkcAomw8RttXYsZWOJcuKMbyk97qwaF+3nEsAowtojsHJBStOdRnKrICcV/P
lAf0p7BqJuzqZ1s73o5XDiYMpLDcCHcaN4rEFJeU76W70Gw3SnzCPADn6ub4VoUH
m2XSFe/VjTM84ls7FY3gc0NHKZz0MooGOwFQSZ6GI0+Mw6Ct5ZMWXlq23rW8Qp4+
KVVUdgq3TLrRwhlV2SRJi5FPnC/fUeovS381EhEjOu7suUY3cW/I8riuzQWHdnBV
6t21iQLKV3oEXCe67O/X9blG2PsEbQjeWk2ZU5eSSTWkbhDoFXX0h+SontCWALLF
SRmmnJIhUJkb3NTDRrvWcMLDovIEItQYUFYubxH/S02HN/AdCAm74I5BfNjbGz5E
vArU8aiLuan5u2x9tJQfKzpbhlzcz3r8TE00onJy/yRAMyOwYE4wZ0fdkeWR9qO/
PJkaoGr1l1Y1w+M9omEYHq0+VwVUBn5e8ojW8+8M0fHc8HomoYuU/6Q474oIRuDz
gu3XH0K9lGVRpGo1lkWQAZprhv3I+K/lPsUoLIJCQJJQ0vQUVE52r1uMcG56x1hS
zxOYOrKbCuLU4VWDJnibuaOzZRUVoFAZuo6cyo538o4eXkTQ/vOnIvCJq3onPRpQ
2ChQgWGe/7VJwwRGFVmBfadvy+wR+pSz3CboRSLZGkmHfzgCrGhsEZFucubM1oW+
Zo99gG+N8E7IezQmF/9Ps0bnwF7ptuv+ylikyRt38RZWAPYS1qu/mR6M+tZ6mWzW
8KZkKupAElaoYqf+i6ghe4rZfLcZYk5/ZPvAeniq9alQXuTuanFpjlZw86kQm7j+
KCBQd0CHYYueptEEIW2QERk7j+C33kDqtfxTf5y7V2siGrGi9OLyujWRezcgwZSt
6XG+asHSVu5eGvKZu+oSh905KcqWMlJ6mVbR8n2qORuUCP8UE8wLtI1RhbaSg23N
ULX0NK28AtAU6pSuZEVaPGyvrGvZZ3kRR5QRac3DKbFaEU+vW1idkNTWzGHpMr9/
AmlY9il+44OD7ny07RnAqWg2zfIgP5gMOCsb7xZlmxyYWl3NjjNGv/Cl0iTlZWQw
Ov5DWYI46etBZThWOIglJBxAlf3or/yCtpgKA33PyZ8qeGUu6HlsaGbA4y9zpmmn
F+LEl0tLnk1FiUp7169lLdDEr9qJQyUf2yT0iKfP/8v5A6fgUBa1ONfwxKH8iY2c
TaUL1ScPCT1va8C/hjGe0wD75/bXiAENyMJxtyf9M1gT/V6M68azOinEOjaMARUS
TuTpIE1k/sk1U7/PPaPcsKnSHcBQC7ea2Elv5Zxo/C4jYnCP0LpNce6u67w943cM
j1aguqsVwL2YO4Ps5Al382Z37ebI6IyV+Hu/FBpAZI5kueOtspjlJjqPgTzgSMGb
AGEkVi4bP+5yeOsNtDAw1WeY0uVvmn9yck+OsvgfNiSRno7kfki+YbGZBlXfHDeP
qLs3w0Zrl80Jq32/KOZ4bT4ViCkr/B8sy1Ls7668GwjINI8DBBmgtZEeZcXouVpd
Lueqwcx84logEbdATY6CkIa+z1bhFePEBWGlNPVL0eIBiE9WMrpxwMymH9GuTD49
bRo9I+FLEQ6Pk2qMqiii4IzclmAtRboCPXJscUPqup7YDmf0gBVL8lSVWgNDwT0f
N4A4pL4fh0+0oBmX0cF15JC4OJNV2MONQx2PIpEA4zGsym71C8akx24aIcIv376W
dSuH1LXU7A4RnZcMB4uiG3xAeyLVPDxYjh8x5gI8gLvhQje7KqMTIottxeI9j5pu
PH2GetHFuOrQQo7Nq83HA8uc+JuCrj1FNblJmAwURov0fQpORIPnJXefdOCrQcXx
6zuvERhwf6SSnve+WwhZHGZP5WSvYT6WKOIsrNsuhtmD+Jdmbrut5eVlA8rrwdLD
3EWifmx/o/LBRT9sILDUtPHcuvPLWBBJSDm/vwdY+2hsHMevcCSRoaF+ItvIbvI/
S8x2J2gBlTjoigxHeDsF1wPjYoLhcjzc6M8dnLpYhy5mcTZqFgA9tbMWFZy4N4Yf
eYZaK86UAx9HzNDgKT3q2liO4LQnMUaOSkJpGifpdzQk6FANBs4f57+vhg2fxT7E
5J7mLk4sGsl/te1RerXPTLAls7PEl1wBElpUjtzRkVerN4p3NemmiX6jlQMOJ6Y2
2Wp6T08VfEds6aCPYBbDAKofOX6DejYcXfP1rZh7DbAri3HlcXus708LG29/DrYY
+l9sADEyazwWZme4zM78RVXO5WxZqwVeOM0R/sd5lRF2g0I0cwRHrXrJLGOYgomh
PQPOirWHpHn0hj0dPST72zXEklJlU/fYTcHjMbT+rfWSQSErXpXJP8s3xR7joOqG
orZeVLOI5XFXNMwKwmuHY3+RFl5tqSi9p+b9VHmKzA98zzvO2o+snPsGabRwrYdm
jb5rATTSclbk9gAsq9wGd6bxXxaw9wFZ0HkgJBY2keZ+iOQmWKB9oxNNG9DqbeKF
rW9/1swVORJI5o0wVkeradJyImaC6d7tUS7tcIF7EnmMULsuWSnU0UiqkjGkz4P8
2+GoOWQDgTv6Q2Mi5ApRjavLXrYq0QEGMtSN1eisNfofmHPrJOCnJJ2LDk0vn8lR
/t8NZjKk+HP8qHNby2UPOfDx2lPasS88jUvB60GaKqvx2Z3me0pBAZ0r07NeZar9
VTjRWBjgD8wVwDQAtYyBFZ2SmeyC4Va8r6rbU7/tpWiaX17vT4MytkCf3fFAXd8N
xxNKgnX66uzqgYs8sfUe+9krvOV/fVyBIOcrWfYMKK39fm7XLOImrguutZ7jsz5T
8ehwkjd7QXgP1+1Z4UgN/xkIXlC7EtG26a6pOEpkYEMyAoxaW0Txr7PUs0SiPrEF
c6iY8cx1OBHHKlcAxGdzlz1GbFI/EV9ykiCNjIJMxKtOEdtFBY55vXHErFLIgo5P
rbIyGL8wDsAgFbZ4ub04WMvkEO/LlK5SZITHbNrvoNq2HcXwumNXexkZTT8qE3N9
qcbqCEbPlOkHQqapYzhpQexnwoGIdHKsnrCFSKywyPwj2dIqfGb1EN3q5CGBNNvB
eqgcv05QYCajXZatNM2UxKtY/qmuV8xfjJLlLittLgReXQFpbACWd+aVvvIJgVzx
fS4QeK49nnPJOqulJeS8rRB/Mc/jvM+jEKOJWcjE8/rmlIeTkPvqrh8GW/ej1iCv
FUKAlC0ouDVy/8UrEe1mOf/iWc6pAzQyk9oEytw2enz5sTUUfoIYYKyRdXizCW6U
2C0RQSTPRRhTIdGbgbxG8nKACk0wxA4wRsIlyKFBFM41fnNyrUwRLEkph4++2Di6
X/aY0jLjWJzVrjc9AwIGlh1e7/1xVyA0aw5Upb3z59bScVvTUbZBXV8KRh6HcPor
lOwUW6t1kfxk/uiw1xoTfeoY1ju8FKpeqgBkg74hFc3Kdxy+gzuN8QOAGCvBIF+Y
/47CBIKZPRr0RF9JlA+2p/9ibYNQMjgr6XO+G3g4wFX70LW+xlcGktBoUpaRD1RL
lErv15OxEvKLZVQHOrNG4atW03dgbCpWVSWW0wQOJtDPNBdhBRVnFhCbZTBjRVYT
E3GgNldc1WlNAkYx0LugPFG1O5r7o0mfOo5X1CLW+by2RMW5EfukB2heWl8OwewC
B8N3Jt/q27FIZFHTvzoP08GN1Xw6Mm0AkdkfQvkgCiAfEKRPROHzYFm2QsSqhNQC
AQQrJr1sNPZ0uUBMhFiz/GB+Kb89AfUpa/UJDIk/M3HTpik9X/09HFoyPLVzKrdC
niTFcrDp+8Zm8wuzLY0DR570vtplgy+ksF1uyma0gt7GE53sXZMZTABs6l/gXE2D
YjSS3Nk9YW6GORJqjEzD2NIHr2+rOCY+VVe3IzoAl6OyRdCNWK7BHyTegQeYF3V9
grR1Fg9TlSwEGbB3noiIqje1OkjqmmL3qKQx0nKB45bOW30ACMLxxHSmhl0UBzd3
IDgWWBjUYixL3K+ZccldIUIOhXVpfsEmtJuE363vtTfixKHILgAvmLXdHv2OVVpk
2CKTXl6Fv1rySXBah6pXMngB732OLxc2E+Ak6fckeIF6X//ofQ0++0MftULdKTyg
Z7guvErUEc3rWOjAOPoJpOJ2VsuHDuaejQVcK3LEbABLm+df6IW/NfCw8HmN9UAz
YIgoS4b4NAqhouYWBs1ivaoJ9X/rFby2207Cec+OSWeOwEi8hmqUS7KMqBKAq9MR
oVkLNjvfu1gz2CZprox+w28nLGyCl42wWuxc8WJruTAj/pah4OT8/XnXp2B45EJ9
tKyPa4oos3gsNZ2/xksgcmkP16K8XB/MdPDQLs5TCtlqynEqyfvr9ergwKtjD7Hp
nlR/6VB3Ym2MvgBoIMrlw7kusnce3uirkh/jyV14p3RS88e0ozCc+s/4wTiXNhnt
C1p8CXOjI/G1Ae56pUKwgMi6Ucag51bREcL2ro3PTb2hii8YRPnQ/oJxFI552r7q
tKrFOIifDNr4tMjaWRjt18bYSRnK43UrZ0r86YW5OiA31WX2k2JnVfhh/z7CWlPu
e0uyNfz1P8B840PtIBOBdIEVcHyoKt4xY5+1xpKBDEELzsXt9o+RHaFte/Z2OjyS
olOFFmMrHOhTMnpRQnNr21HJfdi+Yef4LaaDo+sDYrJuoRFZg97A9I0xMCDfZi2z
ijc+34QqI8xL0uq4xpL9ybHTy8Iv30NehSc4lRrO7yHoLrWZeN810Am1e9gbKkVA
jGSKeS1aRBAbNuWPuIsrDq8+gu40n+3vNh4fOmZao5sEzTVuHxTEascVYR5FUdJ5
IiNDBuEj/drdqhofUa77BnFcI1gTiv3AJCvRMvvp06yXlmM9xNm6w3VzQ8u/kE80
m5zF7GdYrAZ6AwLhE6bJ0C3HBek209y/iz5U8IAkjp8rXkDzJ/v0SmeLzYQ3jcfO
c/xvVG+UiOCFo9f9sNgjfv7Q/9md/FwMIgn/kSOH3Se+VVa0a/wOamnIcTo2QDFQ
KC9rcfKM0slOEAmLuhO/bZxULCylCHbDjGCf0MIBmgUgVouoqk79vqdCmgoTwv/4
o2WF660kpV26bY3KT2HqZzpAw91zhs8DVcDJ7163W1mE1XJbqEJFBGoUSeIjz+SJ
W1iF/9uZkXqONdjDTZhyWeOF9TxdqGfvkn04JQXoBhY2JUcllfys1C704PiKyBpD
n500f7eHBUuBbjyFIvLjSHCZ8B9IbdiZsHsjkaPvRFD8r6wVZdW19ChgtV9cCR+N
jBu2ZHkj7Ui8Cyh2s2ZCl81eaOJWCJtzj2LeaNuDfPmbAoBOet86BK9O2Te1Ryg0
wOfZ4FAIPvMjATXNOlXTFBWFv5SvUvasazIl/iNBLYwjhUcIcbd21lc+86B78ejz
E8WK+qajuCZlOZmBheJjJuytH9PK21Z3bDkicc6k+zsDuzIXjQKAap9spx+GFZT8
qcnIYdWdagR1mzNhYDD55jqZT22g0ZKkEB7cyHyWVq2ZCB+OG6yU1yd3P4iZqkA2
GdOCcWh5UatCJDlx+9C+abaw6yu2O0CUVAJx3BkTjqlC+/uv79JnL0xUADNS/Dpi
SxmBVXUKmqjyn8FKYM3FazIkT7/3dcQXgcJ1PbBM5pUvsIrTrT0BAHWBbCnaqtE0
LKRh8V6jQZRFwpIuG5gs512T0f7OPU05OShM9vJU0KjCZWyb/jFjbNmaoiYoXY2s
IiD2JjkouHd1CVE8zrjdDajiEpQ5fD+5svAaFXQTkr6ATSYgkuyTryESsDRqqoHu
1qW7JTMEYEgAwzWm8rBPCDfaIDFlYnnSsN8mLvoWqeq+S129Fb6iVQTczXRFOkjJ
z9MEOnY6iMVk5GjHyGltJEyR3ijtpF07da69hQ2tNWgrZIp2HfDCmKbmR+byjZsN
R+CWrrAL4sr1MwNNXtWAppIp9+8n8xGVDi6JgWvigdJzSgovW0zrFWFeT3bbsBVv
l98blQ42I1jSv2Csd8qoAdI+sOob5ln+E80jvnwpdwjdF1OReA6SSDnCTc4yHBvG
ivsd8gQ4VI7hMkChWMDUjYZlEc9LrbD1LiRGxwgqAeFAMRjBHObdKRos9t1q1dEb
vGJKIBsIlUTNCuKPksbhLhabyGAE06N/lr/58qfEoMGFZErcTru+gvy4LbmTdmQG
U9hIU4xXgtyPeT1azGAKXIZJIEnUqfznbnuXLdxX6zGoBIID6Q2nXFK/wFL/vZu2
ajQM3KGHfdXojtbXx6S+u0/etvDCp8GxxfsMcPBd4EIfAScjqGF1WGNAE/qUagzC
f4Sy0oh8uVfYcMka9c1tj/sbXRHEn/eqp2sDYOwBzX62/n+R6lbojVF+SDJKuglX
NLnVGppXLrnKqhRNDUnyp2WHlhBXvWxnch+00OM4himRMWVsSmc1czj+ALzdP1Oa
VZqg+7dsvt8+dsMvofIthLPYXuIj9kzLFNzzP5sj624Bg63rVP5V4+LQfBjU0oJT
530VcRmBffTp549PQgwjH4G2YdFSvrDSwjWEKGZC3Mj2MREEWJxA0SSoMAg3xYw9
2yDUwcT9xuNRahGepFo1piLcH6UiIejJl7rL56SwJMCVd4vj9i0OP9yO8TAduZOc
A3i8hSU0bbI1hc909GqbGnEv0P/zyyJg7IUvI8oMzRoScfLiMhDBhXw7jwftYpvC
3JkznXCoFOfDyvv8fooM9NuRycH6yCQlVPmE6kVGQpeXaW3AzMAiPLdTDwUAiDcp
SJcEXsmk4IMHf0kxs/nABX3QR8WIe02JYsX/Q4shzHqiYbQe6z9UDG2wOHyqnvQl
2eNl5pDeJqGYDuh4I1o8mmeHy1UvPn5TDZW2dEQiICVUmHLDZLzt8++JURNLQuFb
BzVNgQimgZdzxnfAVVg7EmfhdsoRN1CWBFpYDzAhjbBbLgTrGdHtNtK8xV6SKTZj
JBOXFfvM8KzWJoChpxM4WZs+tdV/DhGf/INl9WpMimhsla6TX6DC0DAoUI+jLf+Q
EiPrq/QrJhwJkfpsFJJv/ANg0FwtH2LPSTmlw04XxLuHjMHvQW9IsPwmw9kmW0It
zk7sn/xDo4HsBNIh7oEZEFkyLEF/cTUrMXzSldsyoq9PKvKtfC/J+Mr/zn/XzGRU
mBQWt0zD4a+Q+K04Fnvw4osaml680Z9oD3vuVvJbfktQ85leOJbUzuCUvfxqRjw2
i8LWSbi7GEH/lJJr0D9sK9i0pOSt8Jw3nS+XZbhAwXY4jjTBZoh3pd4K4bX0ff8W
GBVb8hpTUDPENtOIwXZhld4fV4NvZywRbmCWvi+duOkfvbtCyv6nTeBsidkqY29b
R32aeuswEDM1uCTNsu0oZKqNuwDN9TXTz16ZMqzn13oCyCQ/Dc12CeBzl+ew41fH
FjZP2UMXqIUEjDVxkHS4pokbhbu8njxz/ifs6dYAjHJNv8b4jNO5YG5kkYlMAhwp
7+zzCey3z2EPmUhmNuktKv3qX+nx+SdY1H6MtTrLYLdq/D4kVaI4H7//phGJrEdg
iZm2ucaIhUm+2m9Kp04uli8A+xE3CligfUIBu9XnOqG6vthUtBd5/XR29758Fob4
V4kgJSUvwxoWjh41F16LTBPa6zxDZ91ZpP7Qguzm0V4BSSBv6jz0LuHd3qOfSKUz
VFRoYY+HUNMLbadIaUnHgjBU/pjmsS0olSfldeC9yq0M7QkZiO+1ufeuZXSUzFis
aN+L2/aBnrG4K1ORcXOLK38xCxMejdbRA8BxeTVsB1vp33UgNEeayUGKw8llZZdK
jrsvZiwzD7HFZ8y2UHk8i/37MswKIjRzhgx86fZlDs5aHY2AuzkgHooHSeooRKyZ
FTPdXZuGpgVc2teQSN45Q9+nYTFcqw66PtUjQGO0W0ovIkWa0wk4izzABSq7w55j
+xfrvgeTiWiDjaHgYJxpN/McU/YQ3IM94kKr1hF1f2OSxccgPxUF4lZvLsGrWP5I
hj4jOYi8H2ix4iOVi7jhoB8p49GmmkuDFwHze5XlJpSPirZDXIjRaAjtQTSum6FQ
AYu8LYGs32Y8MVldEld38fC21bxqhdw18ZntE3cI4GBE7Dw+42oKzq+M0SXzxtWT
QQxPsYDtjfF0qc1GBjIa2k28w1HQbnGKfTuVXtT3HcyAy1GeRaFHgXG0IQfXMamd
YINXhr/rGdFU1M9ON5wX5i+D18e3zAa5ySnKQf0UxfAs7sjKx/A5s2FYTg+XB4AH
ZVn43NGVrP9RWmbzPvw3ELMxBnfSSzrXqJVcO1li+em4Nf59qilek4v5RwthzUay
U88D56cZOoDtUBgUw2X0LPrBBhpoaT3xQTLHPd61XZvqNQBestTl7SxuoJL0VKxl
o3H+QGFnfkgXlRRNPR0QI0bZdrxC8nTWbMAN7ElMVMDnB/1ypemmNDuKb2X9U+7D
2YQbdwi1UxihXrLsolpg0PK9gMZclNCcP9TwBuSVhd8kCtx8HKdsV9YtMziqQ1+T
BrsbDaClQMcMM6XdmBh7WjtKV0DTA0mW4/l90Aonzhzq7jj3WMq9+tLrytgSYmQy
t/UDfq6WiZ6hvqLFYLtfRxCAX+Z42++HzxuL3L0QF3U9sC0qRecmWKKN/sAT4srg
XxHP4fXzRcns6cdjVKS6pDmJCRG0rGPqDjx24kZmP6gDP05M/Klxb2+XiZnDcFDt
MUJCQ0Gu1IfUFP5DwTP4ZOTJL8d5oERdxej9BTchOemeLKTlXWFS04RqX3T5i7jz
yAMjWXerqxJwAp4HteqHEG8kCt7b+HASmHDGymX/Yo2fQWvJHXJoLwa8CCND4zjj
jLRJG3GCorp06+IxTEkbHMdapMk1VBOZpQFtL5b0krGMpDQsS8vS4iALaK95ZJbz
vSpwHEHkr5IjD3/K4JQ+bz2Sg8k+y3Gm5XmaNq1OVbfiTfcCc1NJrd2ci5Gk78n8
Fa6QOT8zJjM7y0wmYVB1nDxC/O4/ZpTRH3jfpfkpD/2FZsdpaY5yD0ZOeONeArxi
tYMcVjCo68gIx0If8gO1wzYwht188+/M4xcuBBdsXWs6QvUAApiwzRF4CIE/1NK2
BD2w4S2ant75JoN2G9he8G03xMbF257Ty5OT0/EjFXCX58YHg5DFoFgPR2gZx/7+
PW0XJ+KtUPA1ZpbLJJdewiJseDxLp+tHMG4gkz+dkg0xazCIgPRWD6hL0V9gUmS4
I5F4ZxnA+CLCSZNQSqmvm6LZ4uy2xNY0iCLXa8auO9Vm38wT4SiDB83AU2Chnf7V
VcljMqksQ4GuXX8wsdaJfWVCQW92rz13jcy119eVky3hcnR8tXj1Ev1Ne96MnPID
JH7kRmu14K7GJGes9bIyCHzfylLpmnpN0ohRoMuCZxee0CGVI2fGdSE1/WizYsUw
aZaX28cpkT89Zg0b4lMLFvGfvvoE8pZKzK/0asHqD/Z98HeU3pLqFwFH5TvujDHi
L4TDI9KhBc60ntarzpOO3T1QFK3YfEuxZoe1sLqI37fRmsQaPY5r2BArfCki/cyS
MYBe0C5ZTpkiXUsUQu6Kx15K0AlWzuCpizWbxewgTrcGehaCjgYPOH+E6G7Cv09d
bjb4rGw1a7Bd1fj44g3Yh4Px1qOoYB4iHNVMt78O/ZSHZfr+RTZCxPrLgPBbBlEk
aASkvuIcqV+NLEdDyXE59bsalagGjZ1T0WxRmXoZOcMynz665hsSjbCLWtbibqYu
YIkq80oN+01ynyEoeJsLyoHSCHeAVTdGXdgC0rcv7Oa6bTdkBoWWmmy0WfNYebmO
VPr2XSV+pgxrvIQK03rNgsVZUOvgHHbPS4Lgi9bLuUtd5m0LcmK+vIwRGtox1+o0
ACfxMZBfW5G+O+KzXldEeHNxxjmlXYMK55zsW886kujdjY7p4dYr69dRT0+teVIr
fTscW/ci2gPsPMwT39ZjgfqIS4cDNQ1GOVEKbTe1LAPwGpKR2+s3JZmdOHJ1XApl
B8f7jFHYhen8odb8s/943wJm2PI88E9QojS58yiCdN/51elcYZI6Y5dCjU5t8+sF
pdlmbYZWi/FU7wtnVzhi8N4d7ifdeV5yvIeRQ5fDKghS5fkNvaeBlEfjyb6v8org
+vIOxS9cOnvVEfWRu9YxzG/UYne7WGTDx6Xrpb/fACW+UWBJv/hqAFiBWhM1Wj0R
RrI4BiA2Nqa44Mjq86FiQGUwTR1i4JFMf8et8UcKzd1RYq9Pvo4+Fe5OqORyjQBa
pwfL7fgL+rwcv/L9iyFjQt4vy+NavwRQ/Qf/8vhy1AsjvUHrBFzB4fRQjzHYdOAB
fqrNszUXYyRCVpE8eQjtvQMZvLUyRZtEg7znhfKGTxi6+h9PHCZP3ob6JRjyZ7e3
t4JqDZQw/WQVKbX90nkcsetTQ6kKEOt/Sy7wJb16jjdxIkXe2VSXb+TMLePh08FP
Ov2URv1QFrwntisAX2HKbaHhuw+OTLxVNdvntu4jLngGS/HBxwe9b28Bc6wjsMhj
tYbpd75bQYrO9s+aVbr/obNtWPxLT9UM3e8bxLx8hiHG8J6Nz/nTyA7peGqHUOOY
GGLGbkaxwPNxxkL2ojL0frP3sgRsMEv588DVRKfzJdtZMsCXv8iCu7M+/aIzKmK0
c/1vrvdQ2/+ali7LMfANL+jXrkJJmq1goSFdx+Fe2dSjoCmxGa7tcRggjMHZ3B2t
g80sKKDOudyUHpuzOoNuvh9uy1U31TcGIL6xbLSEvJfWv1WNLXPFxJ8Yrfii+YIc
6TZTUncRxAjiJYXmhwSGu+cGR7cEysybTgw/3Snp1H5SvdamegRUyT+QdrVRQE0n
aSKM7qP2EfgVQbkRgyGD5JVFZus/2xyV7Lzj5gd+QtsMhjWWHlP92TTzYoLh226V
uJiGPYtwI/9+tTysjvcbhnvFT2pGvLfr82NMBlSmMUUb8ci+cTB+yYQht6pweHKC
Zfr2m8RTqywGstlNZfHvODtTLIZpU010K6jIodcd0rD7M68zS4lfCALkdBihyFIW
HoY5BMcEFI3Br3GSnSLDon5IHMc8KvKYmnIuBItlzOS+CEu+tpLv475lmM6bfVJG
Wk5xCe57gDCOZMJQ38SKZ0MpVqncTxL+hZH/U9AR4GV4UsQizt/l0dixIk9BOyoA
ugcjo9q5cTOtSd3NfH0bilBB4j7HeVewlj+4cJKZQkRbsj/mk9bN8ojRFRcd1miR
s6iPTPDJHJYMBy0qyH6ZzIofp0pc/A75bYF1zlMIpxK3GgCmRwDAUcsGxpECpe9l
WtuJpCGNhVO+ctTMzevGxapuzGGuOsjXWb7DVY1JZX05yCVmOVYKwuBnfs/JCHPb
EOcImb7RRYPIGHHv81WEUEMYScDB9JNE5KphrR60sVDNd9NLZcI6+acaGu+L5f0n
1tDIsNbmpWv8cJmw4PhGduwxSku5ohhNLxBXdTqk0BK3DWWqe04vLrTivfOvKNYo
KF4SxpzmacbB4Dz46vxPTLfqIEe1iqTOZZscxtcyklUQchh5RA3+xKPIw6W64xY9
iUDlVIKNfsVweRLyoCwkNDqQ899a7ZdgqZGCcwljTWCxRpJt4N4sO48IjPXw8TNz
/QmGtkb8deHrd6zrjzyyjjU2FJ1UZLJQAq1r6plZLucWitG6YxIHXW+h6dKAs1JZ
WnjaPWYcbYZky8lYCrDdILURKiGmKkYDYmCZ2iN55Fx9VleF3Y7wSTMkbuPOY2e8
GZ4un5KizNWz4Sake02xGwD9mI6hz00SOeMtYq0AFvf4MhjbxXNxyKUHOuEk3RVy
BPX0SBwajG3M0MVtI1eBhn1A8FfaedG9es3SPrmFC2/7ldYxd9u5aZEvyDbzZySD
AOuRSUPMNKxEBvz5l4h2R//YOZqkQthraYW42h3tTjIPhb6FoRj8QAvff1Rcr4YS
+sJaAY2OlVgFXlpBB1zRfLddDCXDlbpUw/L0QkW65TnNySnViCzrZ2ao+H/2QEBA
/FZtCdI5syQ6vJPGpCEhb0iyN/pkmqsdrFnKetgZfDrGP52GCzjwAzeLN/2ghGWS
U6mhBkpgVwnzpr0LWUTir7170LjrVTfFqIKwWvgM0y55zoC6yA1ncQPaljKutxe2
R0Yqz4OSHpLkeYQ2TiGdkHMgMp6eUioOyXJ30Rel11+T96dCJ4fdLswr2tGHEEon
BzkHtsTmqyvumaXFWWe7v7t7wuEKf8z39Qxu8x7V7SuG4LTYRCnYqmogMtoq3rYx
drrEHLt3+NBHfImVNkvPMTKTKI8DUf0PoB51i0K13bsoH+QuZwpLR4CRjMHWmhQb
ibObHWlkXB3h8ozNQFhWisPpKX5ufLjQWwZcariPZa08NhDFuNJVbEJsmy+dCDgU
jbEmtbgEKc3pPZY9MpC8Nx8rGn7RuEoOW/D/cPQ8BkjRASs+Awa6dTGiHCoPFGxM
QWEhdHm7tmLBmpofIb1+q4nGKr24/RP9vuCllwrOlnIqouM2ap7OdRRilA5nyuyG
T16qHbWjZJHslRrkkwmUYHiQXzQtYQEKm3BpSvFUPB4sSkq0mtiJZCAci1ZEbpAr
9uSqYQqMysFdCOwGTj+Mg68LieWgQHgBEJ5DjtkUc8acwzCa2TtboqmdXmtPUrtM
BCgjmfEUOyUvIQrZYPyjufpaUyso8yym8rJt6S0/sA9QT4AWgCzWMO7D/5np4aeW
SLEbxq9E1oqEpNZXB1XipcrmUh/enBrByXaNm5tvQWWvVTlG1M6l0g5Z72UzMu4e
60w2XrLLBPYgUppqcJb6lsDtTPdyykGkK6mFGTfyMHxEcwNvKGyCZOg/Dam1Nkl6
OJC4C2GD6ocYuYuzzz24yHaQqRDRNecbWuV5OnsFndbbhXN5yEbGXdZSbicRrfi5
tRQu4CAJMr6CnvMcLEnbGVy46bSyuOGxjDlBfqpz3Vo8gVbCsVZ9SSg/PudQTGCC
x1Un7C2u4t/yHv8GYUAvHcy6Z9+WXVs7R7UYpczGm4WxGC8sNbbhRxqLRBJ5IiTx
1Tveg62Vgcye6FQ/hRpQ7z0N1yThaWS0mV8rvcApAnXPSsEKhAwP+chioQn4rxW2
L+iRG+1hagRIFGDKpbQvGLMu2mRbRTp5o3kwLBcN+Grn71C0UQpKCHIwxvMQjXL5
KMFRcMGg+cDTKwSro45s/hUWSAj12HnYBqmdsJ8WnxGphv/NcaobvEa9tCroa214
RxH0FQfKt07FVlGqHlJ9iHJzSJ5UWkuscGnB+Buq2MTfb6p+ETZ1RW+XVnoWGnkM
osQgRxjT9X5WU3FERQQWsdDXRGRv6hE/OStIv5VS9ypTRC73IzNQP0NPKMu31Tuw
2zlcsVAVMucTjuF4MkxF/5nyhYaEW/tSW1ZRQ3KB5OlOCJJy13V5K3mwP7ahwi8w
RUL0rl67C/awL8hXZmSpJJSk3235ez2j45zHUxiP1XWcyBApAnUsAiAt2o+HKJLx
UwRshVS60E5CNWXWxYOlJKfP+uGdM5dntSbZfijf4Da08Y6ZdvIcvy8ffFIKqknW
0nhXaLYY09bWZ+pMFFhxl0cAD2rEKsR7KyLym/t3p/T08fNRFaCGELLSRTR+T/rS
4mt8IbPiJrwmfRyDeTL/G3izR7TP6HNrvoEmlGIucmP+PBZkuuye6LSLoB5Nindq
DoXouDbZu1oDJxnc9zLe4JP4G6GZ53PmxtGk3yB8L5vL406+qG3UsOo9onCpF8ll
bAs9dReFpREThpTuovdEE54eFykwbWN6H9hRG+5K0BZbQ6sIF2a6Mb/oc3aWzxIH
xgMatLsNoCSYEUPLaRCwdOnSDf7fRU+AL38XI1fn3+1K3uU/8MDHZwj9tbgy3t55
JK9QD2dxXYvuDjDHQYKZxyBUTwlfRt2qx8+aOGvpuKXlo5X08+Shwo98RyhyEBr4
xak51vJDce87ttV7EPMD+bsHFMS1PnfxmzZlq/dq5HpcATjpW7q9i0nrAyaWZ4qq
aR6P7ZOs0DE8FYa8ur7iE5Z+dF3Ao1K0ae6YTEJDZQfJZl3N0KopDAc6CiwoB8zv
vW9TGaATRhqiTxqe1+IVU8+6GlIG950b1QzC6KEXqMtZmWypwTROVhVET5jt40PW
o2wIG2hskz1rUFMobexRruyAxYGmatKGLtnMI0oywZJY89Ho0XrS2eB5+Z4SMYxF
iWv+Ns7rKxgqMLfVi/ETzPgdMzXNcI426acIIWaOxwaVmmCONk1qTu35wqUoOKqd
wju86SPqgSaRGNGob0dRDdJdprAc+uiu/arOcykwdsPIlrH+8o1D0UmVU5a81cqz
A6/7fz38SK56qbcvxqXzrlVdR9kQ87bKtWPjBomunsQm+yW1FWfXwSJoiszrjh8W
+0QNuXyQUKL5BstTlXLXzQ9DQeDrplL42rGVW2HvUxZ+eqaTdUKamxlmK+ljlCFT
zyhnZm6w+paU90lmAKVYsSTfTNNmWrkOZpJvZ28Bq+B6n9ppRpRIuHtdnaNV9uus
mb+36D2S4Mce89I/SXxIDvlYzngozjh3jjwALPcZD7pubwBFqyPRQTE1TEzEIqAW
4JcwLCF+vSJUaZqEyIiv0WrqdAslIziSFgLPpkLteQQL0B/9C1ZJ4dJBy9GgWdL+
sUGvTVlGBkVaPXJx3fQkSyB5xIhvVUnH+DPv/Hk/zzm4LGzoArkKFl8XlRPne132
jNUckn+c0ns6e+ZVvBZ/e0pHykigVyG7b322ciivRHaSpEAuEUQDpDGMioeVYZ3k
H411F1nh/SwmYmwXr4mhwdqGuoB8/gOUDcEFSIO1BjQCgmZukSiKZ31UFFC4p0b0
KMoOI/lMBq4IQyuYZeHi5cchMFVxPaq3wHEMujW8Jx7ZNXJZMnaiRqg5gek0zvGR
Jr3r64+MDko2JMoRMCONK/0ls7H20pgH2D0Mj6gZydHa0KH0f7N5Ul4kZJ4B6paR
wnllUA9s45rMFceZvmexKsSN9dXRaEt8ANI+vbFwHIKYbJnRZVEZUsP+DDF4M6gy
RPLd71PWpiRA/HgQL8YrdEzPs/bvH+t5C0yPmmPPTAZLq6LoU934Y5OKYzJapkLs
/df2rengsLOEHpPsxbUQ9rZMvbvtGoNXntcRLbXjzpJ1EYrLT8e2bwJmhsPcOpfW
BRVfnQS2w4p4Cox1wfqpcHQ3VoSc0BA8ALS1QsDqjpJpgmlMzBJ7p+ATEyAGNKXC
9wTW4lMlBXLIQ7QVWQueQXH8cnDXJ3d/toBQmRG25ydWQ0Rdgsb6ttnz8Tj5O9x7
Mkmna2K6usjfCT1SlFWds9DnEGvGm+92HMwFKPW79pTzozNFkmQHkzggXZKcB7my
85K9AqqvxoaJXFT4zXBi28JMVydZv33ghzsG6H4V4gMDrf0REb0KR8TL7sa+kh7X
vttaRrF2ID0PgYUuHtzAuyIpLGzpigrPCTYWmdLqb+bUwQO0Kday4umfgmWi42nQ
dITSbHNArUqxy4Gom+5k8uci3fbLIcsX1tspN0kpLMzM6yJ/IXrrvWqPZa2TZflM
YubsurTx5vpwvnBG05XEL7zDF9NLn3cinB3pDoo3Cs/MBNKLWoumQtdNgkSbjJh0
Hn4NFvRN0HEwelOit9WwFE9SJgiRKYt9WSP9D4vk8OxzR9aJ63SisLhj+UhVxAZB
7lPYOhMArMyXIC84+mJs8uvS13RnXuYiU9hZVJnxnEbhmCXEbdhMhPOJqa1HzRnT
oszlierQo9LKC1EeP4MaChZiSJDBoBXUA/ci5Ibxv5XcjfZxtlXAkpbze0zoI3sh
7c0oeZkA1TruBjFubgDt34e7lllEqXjdvSUOh1BoSlkWvK1UVuDm5BNFOfM70Z4D
gX+Y1JuzyBV3pNoiOy3umh2GCN4Evn8RaJBU5gTqNQ2bk0kZc17PO6Egvl2pWb6X
i5tZcdXg/VYrhK15JJjxXq5sXbVmVspzDrOwtHwj/RzYyGqfGnZ6OD8gHjYM9eN3
LiS40v2rfREbq7YQixu2UhkEBF96iFuqgbOsbektNaDRmZZEMdjN+4W/nVa8p9QQ
KolWTJ2udzLYilOF4Pi0VGkAVk+X+HaPOtrhFQe2VF0SrE/pZSCK3C+Qh7mf9fhx
/kq2ONTw+7h8gazVeKWLxxkO/ojFvyJ4unS4H2lX1b8Ir4xCbli0X47bTdPe4ikC
sbozWa3FlpBhSdfJHXRr5AmOjpRPQa2N/l0N9wSy4FETFqvHE3BKX12Ut+NZw1xR
qpnUpixSs4lzYLbRKLHL59cgOxv+Fqo/BzkYQHFgtldD/PnZMaWKtEDrjiu+LdUQ
D6kvHqqLoDqRXJR9AIJMsNACiU/QZx402CfCa8HPUrj9Gt72NHJOavgcyMfFymg1
PD+wu67Af5VLn5N6U282Sf1On2E01RxDElYz4NYzfock2Mubn/OxSfsqLPghHW8R
xCpSpA/QyhjKfduDkGDKao6TXrKjFuupzSwjFUgZ1pEppaFehyDM7jPJzwSgJQ4V
StgyqGw+vm13cT7Sj2NfX5qJi2/vDGV7r/j5J+xSpT6Fbtk2F3YyDX0G+6FnXnYZ
pBb3Ia2O/9uGV/Y6NVaEHuw0nifbZxGbJp9yYpWc4Ro9cRtyyXhFnwWoGxR9nbim
8Gl+KyQ80soOEggQ6u2DmAEM8/Pl8GFS9j8lNxfO1iIHIOB9Ll/NzIlXGAXbe7OE
8r9zRx7z23i47CjHZRYQ7VMrqu3nks2Rrl5vp7k89FoU+QotkZN9LNj6X0jGN9Ua
5kH8Bfn5YnJzb9cKa3jqKE/OykvEGvIJ6O5z3RbMWQSZJbaYXepOOLxkmwM289rw
Kb4wXUDsHAtrQyiH8xV794ikSBUuS7eAexjIr3BW2gIkVwvGIcz711QUS4JE7sfl
LC4gpxCxneMB4zJH8DGvfxGq7gTq6x4fd7sjEThOCnve/NfmoFtoBPNB1TANA2V1
h20qDrLafapDay2O+0cBvKHaB8PPgU0QDlFIWZi/yzjg2rU+XT/kYJg5ox0PHaU3
zZHZt/YlZnPJhcIWG/ZC84rdPaCUZWqJx6FN76KpGgOLswk+gNO0e9JDUXi7X7oW
NQJj3lBvNIscDk/8ctTuNReZhjNYibO5zb4ScBPPTRF+zMIwBW4M7vxUDWhwV0ma
KsmGyokHytKQuBZMryVU7gxUKKTgBIbcxuBOfYq+kKd7p3dg9/5jta9Lo+uflJkL
wx3fretigDsaJ/4yPYf+xkP81vc+QEwNVA1XvGFccrF0QjnNyiJHJD7k5wqvJNlR
iYbwZmo8SuVIe947bJFj7j92W7JjtzweNgKxaDbJfHPD0JG/J1Dil9sN8rn3VR0a
ZpEmdCo8Hzu038qvltMRF7F4YLGXKGTq2YSWfgUNqaeInbY0DgMijIZ4H5XrnkET
Vufe26JP5QK+8ftzf5jozDVdKnWzJtYJoweDC9PaQVtB5LIRaoB5TYUx3OmH43Tb
3g5LtaQ8i42GwMcYzKYjyekhVOmkLhtLeKYJiJFgLciyAPO7JjWmIQ8hNJM8PDHg
uT/c1wN8jbCZzrT87o8smO1R0aorqSQlnABaYUKgYnNFwhtAMiJp/5kf4VtwS1/H
o2dcAjBupX1uAN1hNvZjb0F2mwq3aF02m41ksZ6iKimTZoRu6LJVS7PYI3OfuJYB
93cW7DcU2id+IhRW1lmkdKrGNpZk2vGL7hbmZAaHHpPYp7iBTS9h1pSVgrMuP5qv
E8ijQ8uMgCdmI8AehzLFZ3Lfsb1pdWaplPRHT6h4H6jJiCsbVudh1rMM2BsoQCi5
EJ9DVSlw82KHTJOn+t082ee1ax4AS30AV1L0caxmE2Ew114uDJtrrLiR7e0zIoYL
IRjeootcyGOputEzz0wOBwzTsEMhhdeJhkds4AX7i5OSruUPCDFL+NFwIPgwhFga
SQ5FIlDLHYS9TTGArAZMPrUM14/nSkUGPs6184PUT5yycawilGDmSpbE/dLhAyMj
BrDc77bLEsXm4VNYI2ELCBWM9MBL/jTDrPUIbGWap/Mwar+RygZtuWUQKcmdBSIG
FzAJVdPhIGn/yoRKHI1582FVEI+M09hTVS7rnYi/pzHPPt597OVoDhpS6FcY7RjW
Tmr2PMlzA0lY1Uvv8Gp7ywNhZ0t9nBEWatGgpLpdRkiuMzMrv7NMZgMIbYwqQOG2
iDynIcldVAgfitnDLshM7rglwlCm4keX70jvp1NhTjlHz0zZnu7ayovYlP12t2k6
TCRYeCrGC/urYBje9vYOveAaAS8GKtlgopiPQgfEVUri9DKr99UlEShcm32AykN0
n5mG+8vS+PBgyFoPM+mjSOZzvshmtDYTE/P1c+XA/9/2QwqxwiZSI4Afnhhkr24q
I8yDDivUWynwDwae0ob0p6H/1zwEJPujobgim/g4BdQxdaP41PcvsLE23hL1AJiB
aablIXYmr+o3K4BRWg52V2KHkq6Q8RgJk4+gqJk4cLuRS3Pzo0zsGoYU9gTOqmAs
xgeI5nGXP/ufB+a7gm1EqADCllygAo4FzdfNWgeNNc2elw7WK47bwVaE2Pp/Gv2s
Lt0cpdfKD5Ab1na+jy1tiGoup5w84KhzfqVG9D16/9qIKfQEhw836fR0CJhqUQ6X
71xIwKKuj3h46wAwYkjrB20c7El6KbU6B1iKdups4rs2ZH5ltrBRpYRxopjvBy9A
JgQgZTNMoU4cCbbbfrfMO4P+izI2bBXBjlgMdl7+U6/b5j2Y44+8mg47iP6aG+97
s3AFfQHLkgzcaTfwaR2gqL2TTBRY9FRRsC0yqy78xKszddQ7PumgtgfvRwgvLzIj
dby+VhPSZw5f+c4i5beW4LxrfKumF6nuIKKzoruTVylq0V33NY8bqUbynLvhFU5t
aNVzmsdH7Uzc3UpNubjD1NsQLJgNZl3tu1UVdQHw5fXi2d5ME+Sm3vkdP1hl7/BF
g6/1Jc4YdKBkr3gh4twDiYCS2xlJozjKvKg8WdP5e6twwNQ2D1LicyNtDCV9Y0gy
2ZGlue0ELu7ZHT/vPQUS59V74D4y/KocGwuS5daLUtLSajNCfFqf3+/JYIKQ1O8A
EpYWpGOedissEYEpblrvD0rYPh041rHAd0HfYeHmBOBZUdTQa+BU5AMt/idKrvCA
PBG/Gzjb55hmFmC19fiQ0NgzBV98gbdy12hRWpPr1y+/y+RnDXJB+6iRoxRBo2l8
SyJsq9qxyTTO1Dvhb3x8C/KF4TUY2WyJbEjvesyVIt0E9JHJHe7L9UUYSV4PdKcF
UoqIo0PtPY3RdHnEdQy47K8Du1NwHYw1t2/kZObz4TdumP3FIeV+HCsIQYkSBpZ8
H/KhDfiC2UsB/JeXMPi5/G7gi8Bnj6tjJRQN+1F2BY1kzT+M5SylVh3lhTm5PlSn
3mll7jiyp4Dzs+kcH0acS2SW5I3CzFg9gKuNpIEDi4PevRrmfkQWSmQn0FqCZCBX
VK8eZ7Nt+NyBUiu/Y6xsrvgfyQavRGYO/xUEwHQD69M1k4IqeL1n6etAZpLn5qg/
jrl4g2uXGkdUSjnSdrxObXaKbzZ/wFMSgqGpfxy7+95O4QxrrmEF4wnHfiCCyWLQ
57287t44ce/M0Zt6AQ+xpmdxROPjX2C+Rj3ZmW0vci1IID4PG3jwIdXNLzFMMQLF
BefwFjN8+zsU3uoe4P+3ap+vJQJshow4KgzqaK0P1TSr0XS9RkWDSPFeLskpHKoj
YG/Xl9E2JMVqMZ3J06VE2poZ8s+Pp14YWMacbg43UiukaZtJT80MDsY32E/aIsHV
4o+lRVH3NfS+AwmuBbQVuw1Lk/Hi+Rc74cX/GXKpLqfaT6tkjrWBeznT0xUiNZMo
nNMPqTGEAxW7ztRZXnkpzQwDHhGRc6Si2fpv6OXsd6RgOvxuWeeTHDfbam9EzxbK
SaS8j1fu8g84WOex/NmA7pzJmzXp1aEN3M17Q4sDwXu3HSzr95jyN2HcWE1N+7aB
4zz8AJiHeIMeR3IipH76rNIRPa3HQklHJOm1P0NDk7b4LFiEGu7huXairtj1Ixqg
vJ3acuGZj+1ySmjlpHh9TngbbsdnP9eDZ3S5kE7dZFZKDednoU/rfwwYdbxMoNZd
Wnh7/qVaK+lb1fzWTzqsvsYXwWqJF2MQpHPHusLmMCTDQ8QwKefwAzv5BtuJtwGg
vxVz4O48MgaBLW/1QU6CPfrw9E/GMYAEIQcaH5qJfDNWFjPA16OeihtRrD8VzihL
R8plA6Seubfx3ty4nTjFZfNvBnmQAtbLL6cmWInl8Em4WUOe2y4xZho6qRNWkw1i
xwNHZsdpq/zU67h52/N0Vi8p0c7A8ZvM4NbloabalPBGGqvt+8tEBazueKY6nAiG
NlahIKLZacMFAWOP/gSjUOcME/k42csQl1+O6N9zY74lJqxd08EPq++Ss1ExIIpT
07Jqtc5KY1xi9UYhQHGaWiagk3PtZDAo2eIcmiAzXPPckh9VjTl1Q6J3g/NycTVb
1AwwBrufA1eF626xL5tEE/mV1v/0fxJwrbwavfjUECTzwVwgSnq+cr8Klv+W2nrA
zWA+yOHTnMezBevUZEF4xnIfM047xsh0MENMAb8HTurmdYR7dUQGtVJtx71nDX3s
yWcb2a32ZF97Hsq0PHtur+FcDlmEQ1URKQVq3+02hVg1WJb/pgUoZhBTWnJ1uIpQ
cnbRwKVykKjw/HV5yPad6kInjRuFb0ML7eqS/OceXGLQEpIR9v8GSka48QfLZs4a
VMBJSzd92mYYM+/eDi3GzB8m8EPpsa8VS1phQO0NTSZ/Uw2heb0Z8QRzLG4qiX2Z
Yq2DYg41GKzH0AQSroWkGbxYIkVNR3k9aATvt2KMspn4SDpCXhdHep6JS9k8TmHs
OzoVTsIe0Me//DjLMv6gRmCs+qANrTZL+c2Rmp+1LUfv5bXC/S+GHsuqkZpqemf0
Ia7/6qozmLEFUk1DbUJJd2jT8EA/A/zqPgb3xWoD8PxefmjLWP54UJW5PyFNW30v
v1CaHlet/icZhGH5TKNbnOfa7mdmeD86ojzdgwZOqedTm0dGriA4snrbcgTLz48T
qr9TPUi6KgK39EvYSG0Tiy7usR1x2/3VEyG7wtxb5qesz96WBgLm3czDvsm1eahM
6j1ldDf7b4hg6wZGQ6KLOF5b9xuKLtd1ivVrXWKtSY6i/glnltUfCeuYa1Kut4wd
B4xeMJ2DXFaeiMFDCs5Ja8ooStSzm+eOmPm6dRf1WyfrNWTIrAvoISyWoWt3pvSI
K+h2g2UT4V3XqsKlXEWJmA==
`protect end_protected