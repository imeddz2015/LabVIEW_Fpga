`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 20736 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/59UwEX+aE7FohaWu0/8IpTj7mav863zUNIsgIH2BWb
Abd9opeuBjbGF/waQMI2vMJTwD1ie1YueHc3nSNpEh4OXp8P5ybZFY89uyGz3ztU
W1EsuUnchJoQgbHZ/sLbgtGRgsrAFn+ZoIeGN1d6RAF2wAESJmYP8zw+p00RvjZ5
pBGEHX7wooDexzkaqKS5G8Gwg3yBAOPmiSYdPIEVAIHLnId8yNkOgdoCI2eKMHsl
b7X02XURMawCiPLIjo4I1J5bRGtj/EO6/ue8C+WvM/ceULi/PV/RWhPj5zvxXBtz
e2GaDSvE3Dy4xNZSqbbJueGFuTxWEEVHHkvlwlULmVKwYFu2q2w4BFxdsmb9NzxG
CKcjal9cfPiaPOpK+mrB4Qt6nKEZd4cgOU4744ird3T7t82mZ7yD2/ex6Qe29+ss
HS+1ukvdwoMiKb+HkmE9YT7JFxlpO/sy4psECcYzBDugu1sw1GuLK9nzpmWdHq2P
3HKSTqhQWUzwI8T5QxgzJ1jhdjgCRIl7I8ua79NGS4AhGYnLDvIyR32OATl6Qv1G
OboGfG/zQPNUp/3pjjyodsacPudtgpKCen3keq2tfRFk8FHbzAXEJDIoMCdV9HKG
hCUg3id0nmYNnWP5z2tkk39y+fI9xoGmuc1PKvsFFT8BKHTSOAJ129FvHkL89FMh
0z3dIl+6N6hq4+nru1Lv6APFk4l9ttoc2JU81fHvxkJzJm16V+tCbKbiPa0d+ao9
KSIIwrxjsWYHa71T5MKI9oDqSe36Kb2OW5tR9yrEAzYTkmEh6ajE+bsgErjC0HBp
0gwoswgf5FBQweEzvu5zGiyaP+ZbzQDSaJ8Dp/Bx3zJw/MFK3F9Adp8WuFkCjFYK
wM759lenzMKBrvKA75tR2RfFkn+OEMVE3qLh13XFKekdKjGHSv3v1Zr4X9fIZYDF
Bp411lu/KQfLgJEF27392Xu6MFp8kM/VR7rd0RrEkmkqeewisajDkDtdQVsAJC1D
mpHUChrx/F9od61FFYeCH5cWrvGKt6zlTxIzjvIfuhdYVndAitNfh7jRJBXzTGe2
4JKpZnny4YiJCv21bBm2oKkt0fWSkQAnQ7VXiAioVSANRYGUhhEK7rHm0LjUEU5U
izdn0sGIHP5cFQr/u0sXRSpwmD/pNnYk/rz0SiVplCLT93iQUQawIzSFFdA5Ql9h
+3i6g9P4uJoveMBVzLdIPgpduISmtl+N2RHOFWKqQnHT8QECOlLVyNkZGKXPaSu+
cIOkvheptO+u+KoYjJnUPMr9h+IfRcsloUyev2vJqqdFWxCzzdt0WVED4+KyT0DV
MTb2DbHksr4us5JFQv6PjtT0LE/j2kRKKg36y4eQbsEqmFUEwysIiUnWC4of5sLZ
QCjHKz9q9unYsOktkoSMTqvZwp9JL44pn/CPyD6w/4T/KQ2k9XLtNvYEhTMQVUir
JTyTgZnnET4AD6hj59IJ6qu4zWm3AFouSuiZRw6akevKY88WJDeEE+ddpyRyCzVO
0QH/78LvmVulRLqOOiiLY/E9bA4ShDkz4Rlob7Vx3rfk0FpoeXOnBz3pkcR/Lhyh
NWDpV+PGQyaNha5k1UhLTsvnulTg6HiJOoWTe4IMAwqsnL6UI0MihIIK8XIL5O1S
rI9PGOD8DSJpLbNeswmCdJlM0OsQn3OTrCJbjRCYxOYCNA6FcNC8Op7m8SF7I6Yv
duxTgVgjhwetVQwGj/JzK7cU/yERP2xmjP81n7ae+ag3vrEgVzqfzc8FgdujVzTe
MrIW0/e7r6grRpDu6KBcKLwwbG52/38QrxSvfrofjg3DPEibFqHU9heuXU/ZkFot
fRxuShYsQbwKAivniZzRzxvn1feyPTPueTw81O5h1I0iDjE27DypGrgEMTiuszcz
/1i2vnSg+/IhiTya6mQjQxSQXozst3cFIUQnkaw5IgwzeSWjOwgYHQFTunGSV37/
Tlqp378Cfym9cDy+YHClaeeololBSD2IMTwiFHZlFfVNtXukE9In3LVE20wZfxUY
nzdqbv8g8nuIaR5UQax/Bi1jz1aTre1BzvHPW+5Lg/ALAotTEPi/pPCHRybISB8Z
sn/v8aoEZUNyGKw3yQ1dEG3LDFdBL6c8mCOvJ3reWAxrVnAcVI8150TyonUyYq91
EBVAsbWwTFgmOCQA31W3ZUGkZJvUc6dlVPFBjtrTiei5z75kmbxBVF4lMAOVGk1a
HRkYbfhRIh8AMep5OFVZ2cObLIwultwymi6osNlRbIKPN9Fc5cEzTJbMWCv7+cLt
bMhfuQ63RBa8tyOdE+zhwizzR6YFCDpJYwFgpgMxVbYkwlPnJvJkEuwEHKbvUhmz
PbpJxWaOlrvkjl5fH/doC+WuD1TSnLSJF95CQgeHXT0ud8T9saAkyXFfxeJHuz85
oDTuRx8MT5kk3qTzalYkhqdlZr436j2T7V/4A0wcoNGWXFBoc60qApPmqQajAtJV
Fj65PGTp1bITaUOAF29+WbD2VDDZrKzn4Z/qJ6B6K2laV8kvhkK3jT0MzX4miAZu
CBC6A0UYigNARHEpuxc5brdeC1abpru9kkB4PWUYdGmgGVAbYT0OFrr3N/4NF5xX
N4z/Cxb6Ju+ny5ENnRnaBwrCeGV/McLk93VvdUUGouOlUBf9nSmefU10ZHx7AVNl
A5nYgn/hwcWNVcJoVBJxpvWuHJ3RyeVZIzL900AkGsWjo5/LXyAN+G5IP5py8gsY
W8ujMTiD2tKjFa0X68dammGMxejAttotcNrkTVO9ir55qCvo2U2GGUZt/9+I/qFG
QF2gZvPbgZldFpOzeoK66fnkyzUgiQuNCu72HczX/fP+6dPhBDDeKd5//iJ10b7G
LX+ZtXhnGNGjhvwTf7R2Fa0o8Y3QUc2YfhCM/ipYIHPg/zQyHV0q3Ag1MSoy8h8O
LVp9f6GYpaGgeHbW6QlHk0A3cO3BPajN0psKOuc8mkhJjY6nWHeHs/YIiDrTVBnp
2Xsv0e9eO+vWNYuTCTwK5+hZHlqmx7G10cEdjolNzktviuuXcm4GZPNcLmLq92n8
8uoD8CzT4gxeI1oJg47/cQNX4nioh3ObL1/AqDVSpM695DWUaOYudbfrVYMZ1BBL
PfV+YNsdFQWCIGF52hOKcacWgvw4+HEQT4pxfw8x3WbowwaecGjpRD/v6HDJ2WED
piaTDKNOW5IlRAAbGpsTzq5mt96eXyFp0l+9WNE616L+lHBm4iZlpX3E6DdENrh4
8PF0WiQWsSRJE1Gkz6a9QEyb1OgaJswi4zrj6VOUPJzfbHpdHobGNcyMCk1rR3bd
KDbD81RfLDTph47i0hRmWh90L5FBMKfgF+sLfXISV2gFu+SnjNTLWxTvNcNaAI70
LxaMVX0dsMhMGZ9uofis++o21T0TI8JdujKk92Cwz8vdbUiHAYh/4B7BDW4T0Sqf
0RrjsWxKQ6P/3YPkUTHA6ZT0m7N7I522t0i5AdVrKv0alUu+mTzXaLBW+eshdec3
Fo1cIY1ClanZyXWa1WLFgh/QYjXskLb1z7GBtMhemcMWOf54VvBCxVRrTMuBlm0b
QHKYuSFQ3np+wTuV9Sb1JmTCf0vnHViQU0xQyTWesKXmrev/LNQwagCcXy+ebl5m
haSFofmt2pg9Bj9WJhYVJ4/MMWk/Vwv2pWYKXO47axng/5Mz3J8rcXedIEuh+uPH
CJTqrlEIYQw5UJh7D0mt/pIXBin8p/KcyjYZP0XAxPW+8F35d1l6SFTOG0xgbZph
NKzvfOCS/FxXB1hyufzMZsw+XfihyI5dx7JGFr9yKUKoIE1Nlt9/uEo7KSmecoBm
O7k3TXp1cu4Rf5UUftfqPN9heNM1pXCb++AL8wA432ZiH2gTyasjq6JzC53CCBtb
l/d4R4B2EMehMa06CMYFTOVyWBB1C9jseBs4GO3Bgef4P2ymutzcMIXqVc9CMCnq
OwHF2qcrnBczZ8ojfBAjYMLTi7sMcypAqJShKr8LNV6N+xuTzw6tWze+haRdv4EP
OcuGtQ0rKi7YqVXkaNINaYUWzPAY47gsj5Mq8qlMBecY9cA0hkPez8/6gIwJ8sS0
kfznP1H1Suwt9CfGt3Svrahgj2bLKArJNJu8PpBc5lZkPgz/g44xwClMavor8WxI
gYx3WsbUnWF9sjbDEp38lplt5LdFl2CXm73NSjSEHYDCksXs4iIguqZo7jpHKQ2l
GQzvIKFDYrdFUi+muabS97jn1Qg5lUvd6MmYLVnKYUX3EeaPs4hyRGllIdWh9G83
LDhke+4WcF0cc954T/CzKo4A9gv/v1VZhEZ0wvqJhUhVXsLyK7wsH968YBasGvGg
WlOugz/xeM8732rBRgkJzKS8XncDhIq2+85LCEtaRDeZvYXdUvlWE6e5DkYM8mqJ
vbB+CVWlsui+b+fD6lUS/jVnuwWRygWeV5MGuCT153n0Kcxb33PYjmKFekmrfW5j
c7fTAR5n8+IYTho9QqEldbIE5D2iAGmpnIGcJwNIwew8DUovnhXwpeMFioX3wlUV
w30fAQ82VOafyRLGgCAMsS4FGVqVhc+MQztZWubiRa/HDZidFFHRgNxpJg3hd9Dt
vm6tjulBifDrPv9c1AoZQO7QJT+qS/5xlahomIwyJtZoUsONgEm8sWJCaZwI22QS
D0wVU6o4XgKCW/LNQW0p8fL4dYcPL7w+1Rvqbg7uVTPp1lby5EXhxUjDYzdrXadx
H9w/ZaYYENKjwPK6HpSK4IXLRpCRijVUxziK/fWTFFOYcg1SQx9yVFpye96uw4pb
iMe0xXyxYzrcnA8WK2oa1D0v3SFwf7iF6a+19SiMOPKNqSTeBpJ/ebpvFhpPHJtX
Zz0Gnu3e8y1Toh8DB0bLBk6/C7xowmg5ZppX2HccqHHNxmSC7FLS7kCNKmcyu84L
k0iQW92tEGiiTBLojlFX/HA1pTfOUVk83ehw3i+vJwZZ2LCB3aMSaKhXzuJgvcNg
VsvCox7899+ZqCb7MHuOJkpacNk3adM/4roGEnXPiLXWeFhZUe/DABecqbWv7TDU
PK0tBGqKyu80xTED9fHNKvbGWiFgFD/kOmFid2adtczP6iqq4RoKnESilRnEGW3G
tGuiCmsRgtJN1mJbsN3ztHMMv1nArILWfWtZ4jEPn1UySbp07jrvQsCYfdvDM6gv
Pi0cXC+sE4Z4B+pajejg0amTXlsJL6cif9nCAECI7Uc04PgjfJXLp0dgL82BGq+8
qsbvc3FdNiHmU7OgMO4XxJs3T4U/7UrJXjZy+aVJtliCSZqWD1hUrOkVqPWxpREr
gLMONF6ujsKn+QFVi+UbOcq1Zbvx+5yVO/oLjbD1d+sWtKyxyXHl/9Gndwo0uWdH
MHkaA/rTOW6XoVeJOHYrklwcsJDom40L0RbLPvLguWaoIf00/yRq2Z1iNPwEXvhx
xl/yd42/3wOqa06tjiznAb2IHyYAqVdFmktOlnnUxdXUxslz2ACnFP/PtjCgTKHl
3W0CVhkJD8BB/GDrpaHa7VRJbCaJWPbzdKrdWchzNEv+xC7oZCnl+uZiO25Ruud1
HHQGpt5yEdYYwlFx7DS/Z8ly3mcAA7IQzo8/8hnebgZPbU3aeDUmvXbgx7d2jIj2
HVlbWF84fm4IEilqN5Np0VQ1Q+TdIEPfXkLoxs3tfoy8xmooH4eMLs6GlpoMWeWP
Dmc8zOJ+04jwViPjU4GF9COWOF8IvQ9QXtzrTRBz1lgY4eSubVz1rPY5T5VCzjzL
BxxGLb6wvVqq6FDPrNzPxIy7/iy5lN2k789w+ycGNlw1v+IBs/RUoFyfCN/ake9w
/DYVLgOMNVC/LSEyWgjtZaTTqaxnTcfbPCBuSCtxHG55GXhb8uaaN5u7zWe23pzl
jWvZxvmsSdOrL7OAR9Xrv2mdonGwzbyYkLR+WYXId3HuD2WwA07kU6dL6UdXT8ny
Db0RzvNbxschupnLA/U/EaRQATPZQlbzX7YQXgU5oKT/T3h0vrxLs78Yh8knH19B
iR0zKXqwXZnYBO1XaEz+bFqK0lOlpson9uWA0zrWXnBpp436Y1sESfWOOdoWKVXZ
uriCau54Szwi4L1TO/K5UihFt9gKrC6AbJIJdd7gJaDiJ4CaaL5LaC6mEctlJiSE
PDNj/AD4AWSWkiKfl+ibWPT6dGTimguB9cMBqlWXATB7ToKEPCoZvVcmpbfZMkZl
x8uPgp7DVMdl27KQYmMN5QG260ODnKJsVGcE/43GkklQ16inqcNh+RqM4eNpKxCS
EMBsKaWD2jG3pErkI0tGVwkpuTP9EPqbO9+ONvxuTko6leRk8WahwtHWJUhIfvCI
aqMvbBObB3VhbvYeka5eY9LbZf6TGjmgd90NinpPMV4msxEJUdY6Z1jb1voCjR1t
wTyUhJubiwcBf4E7ZlanVQGbZfwkGrac6k+kNSs6Q2XYMKzx2NjFG7kFx6KNsyl+
LjJR9Ex7nwMaRv1Z8ai3hNhr1djuZ1DKDQ9WPb4k7lmC1/GRxb81QUR0SVYcMnne
csN0MsaXy403YsJh9FUd908GwvoSMb5yHOz4NS723QcFIX1ueWJrQQlrhpBwpL+m
c4moKkpTnQT5ycd+aWXKdYXzMnpO7NKWdVWmmq0qg07M7PRJKOmL25WolXzR25gg
F1wgXgeVNBfQfdB75Zp9cbaKPNpDsWOBQLontq6H2eeVEyAqOAowjuK1QE/GWk3t
mJYKFpoUcfwsMPv5OVJuRrjxN60wVyIFejWuMi7qiMtEtivE9IChxguCaQjwQxym
+HB5nZx8tB1LW6L7fE7Klfu6y/M2NzXAyzeQdDznh3iUEaFCy3BgFesqbH+gr8xk
3ONp0ohGNheQi9Um3wNePAg0orRe1LTNaPdA26bqdPcOv39JPrThxDGP/sQcgESF
Y2yr4AGY1WugwunFqVmn7ZglJJxOICzyGg7XsECdR54Ki3QqjB6cs1iGvIBI7NSZ
hMSNEjCk3Kqk73KiPTrX5bTlmdLLVaeDvUwNzctqI2uWozoWjog2CQL2rRA1IIyP
2tpojrjVnPDVnLp2BUslASMRSfqYQ7/IHeKFOONn3dtwkMpO7c7KbMmCRIddJhQO
/GTq8WoMaGaoi9c9Rtx9rnOMyZvmUvV+S/K5/VL+xhFFnFSxPIatVJ8220fvtRMN
8JcH8G4lGyDdWseGzITUwD7qah/zNNg1VgY4uklKrsMQJ2XwSq6v6e6pBqioOQdf
r2YOkFg+2RFMsqJOBU1e8DtU1YXv1cUFhRTGma+QNVFf/Lmp3HPBNOVPcTPfo1f+
k93vKECZHXle3UcrzXMp7OyWaLRYpJnMTeYxET5tkNT1akYlscswYn1axuOU5Liu
9wZgGVQZ+ydCvZ+FNx/HRYwSKHSoAXajybjHJvyQmVkFGviqlXfV5qjscua+NsLK
CDVXHDP+f+JSGAsAhPE2SFjOH8dqDZkki9fomjppcybhrfCpSK5B0zsfF5pe7/Ir
O6iuGBgY2kJUQoHXin8rUrFX2bL2zR0dIQIm/yUy/khNNCUp8R0+vcLsFzB+Q66Z
OEJLn6aBTOc7UXJK8io3LPs3ZRUwUQh5FgLZisbvOstwP6b2a4e2M+c29IFU71Nx
+fqgknx6VEehIJpOscjb8yNSz1Wb3/F0ZxkD3JO81zpNlO5IVjej8lGUyLgxB1pn
JWjx1ho5FY4HnfYA3wdemNKvPqIqSg6nt7XHF5BATuRtLxutwuapfDQ+gV4Zq2+6
jH59KM2pa9HFVXZv5Wrlr8nQWsfRGOlURXJwXNayqMcE2Kw8Db+zl8zjWc6ZVoyX
9hjoAI8UQWFj6vpRgrl0UDvSwFVjxXctatTlvuwtpI94DC484dHTJpG952KCWlFS
nJuy7xKKO56p8K1z25KjJ318yDcVAK1UA6DLIIm0aSOYJTwPwuEVBR5KCekbJLOd
9NguzfrIzP4XvKAxdzIcVggHc10XODvUjVD32zObbVcYMo0N23W3pbeuggkXJxS1
JQzJEUTEXAG5S53BE3vxeDriziUhyKtRLB4bXaoIamOxFe4PB59oxpquW6+rDHkW
Nptuymqn3wvuUHl8JqcXj+gl+fgzeUp/5b65RoAFViX1OgisRlSZXx3XkeFnkzmD
9e2atHrvr3bBBSRDL2946gp+j9FAQHRlyxjBq9Dh+fB3G2YoXMPGQYEwqTuXwW2D
4DT8RzePlM9Vnys3I3M7t+dIpHOJlmT+Vy9SA9vyp+s9/B9v85x7Ald8tgfyF0FE
X3TDmgpGcCXAytDj3XSY93Nw5+wUxmSdFlPIDtG+D6/WVvpwa8xKm9Ea2pa89nkp
aMJn3EYygzuY77F49VQ5oY4m24zgRnh7qjIkydsLPPPnLE+K3Po0EjdwSBDZhljr
eYlG3d/YOhyh3Sesh4bcztPPl3Jz3d+3P0NR2GZIwXFrlIkUWhLNckjUEb8vjIhq
ohsrDUUvjsYke+bVWcfMr9SMShWUKJep4RHsRaDrhGHX7PYndON2ekGHrfuGkImo
vcGJ8BfJDBOZqlA+sULldhzPaUTmxOH8vxW6BAuHIb/JDwwbgGfS9ZqMULtTw+ef
Vx7wKovCO9GLFfIB7+AsO1gsJysEYwRiNWQMX358RbjwYHEM5JZuMgreP2SnLrhF
oVEZ160zDHRvMXglrrK+LdsFmSggh/plC4PIcTlLSl6eRCJ7S/Z5/HUMIFmtVwL+
zkMWb0oobTNU3Muq3tPu/ItSpuIsYzmIibAbRH/QKXQ30kgwIHdonE45zIZLQwJZ
BGiHIaFvE0omLaKKrRgW3ZDjMhjRnJD4ScVbROAZjkhOZfj22IKd6lDef8HfEYKu
+b14+AdnVMhOmoE47qoyZOU9fQsVPtMH7T6dTrzlYnbRFgCV2BIl4uLLY/zFhMJt
MzewtB03tOD2XxOaG+1S18WaF/fRZvZ7upoOzlxG8IRJ45rLP3kqAyg7RfIEyY0e
85C4uafVqNoHat3LMz+YsVigDQBGmwWS58IktYLqF9kKKqfUb0FKJA8nlpijuoxr
hu0w3PG2Fr4oxXf13/qfW8VjifRvtd+4i1XAkbI8kDidf/xNZoq62GgRPsOjQUr0
X3tvFakFdrnO8V/muI2Bd23WqdepoELiIyO4wG+3ym7W0ZUnb/cKm/jjuyMpahJ4
o1kL9EMv6t1Tx9dO6Y15mW/EQLr8UKTsD1K7LO2dg/WZo/hjIBD50+3ZGK7o8CsH
YJO9f6hx1j6jNRkn2MFPgFgt2aPB3mSQgtQYQfGmyVjyMGNqVYcc7j+mIDwGuC1k
giMSghF8K9LCiIdLkbKBVJMQVsUloroORz+Pd5sPenaSdMbdbkjg2T36tq7A4fqm
+Bsf/nqb7CZpttXMQe5/YlIHCTX5v9xmcEEGRSkRrzDOBle8erEeMCOKMb8X9kv0
MJwiwAj2cmjqWbFXyHRes2FmzSTn15YFkodavpaD42egDRBo19s5y4RHYwSz0nTQ
xmmBP1JnSNc9+y2HaTTUFRElt/mfYh4ANoj+m/FyG5gIX6sP9ZOpIwUS3AvND0tT
XFza5w9UtvE3eLz5LFit+IifXE82Q7vhoeNzpV6HbEx4b0mrOhFgoopcgm5TyPxg
7TfuHYszAFnhAT51fHCZLIjaJ4rE3UBkkdIMTAD2M7zJM2m0yTxoKoR9vj3AHPZh
hF3YvqAUDdWu0/HB3owFZlu3djSb7p7MzEDa8SpBFDHC9+ZkAkFkHhvvyEuzcLNQ
12Z/VVixAefpSw2dGn2ySXWE4eQ3soy3skIexqz5A46oEenxOcTwQph9BAiy0gt1
OFIrbc6Fe2OSnVjOD5BC+qwEOripx2FF5B4t9Vv0zpiBpA9GnsG5FPE4YoJ4ahF4
d+8nZxlbY5Oq57EGKBuGNwiejVo8BNMnX8txmn/Exu+obnEQfTXeGl+1kjpkrrMT
naA3EOvtlUQPJ/esbq73/P/Dvc8vfGuxJIeiHW8KlBNS6/duvapB8v4bq71SVv2X
o8yaPVzZs/qy0NxdlVMCKuVS2oLZ7avI8E4Lsko//LYOPcQIwEXj4aMkuYNInY3w
JJ5rJgehSqhAepLrHMVQuVyscDELRlV6PjK+Tp/7yPV/ZNnrqnt2sQjlnVsc7L4O
f4XZtyhOiPvT8ojp+MAhwLSntARlsTw1m02DvwRWaxO8MP2ZIDhlepRdkVZCj+yc
aPtmnFCEeCocuuzUz80QfxwUKNXC7l2dp6bF9DgokVLRlNu3fR5PWY4AR9sqDx5z
n5MGoq1ZqxZTuQXhhUIZvgml3GguFFZTWBARYpNlGkOazQuLvEWJyD0SyqhNEDeD
8Oi8TvFQsoyQ0qB/n2odsTlAbw5rjkMtWmZo63bwvees8MInIeo/G9aPGfO76dPo
XIiYkDJeUbZ8chpGLn2y1RFNkDkR93ZJJBxUggg9iRTz7C9u2K+wprTQ9V6vC7Sj
rtZXJpkmJM1s0C2EE9pNIM0zs8FDIyvEzkjtpwOPbcBuqInry8IHmyK8r9/5hUFU
/9R1PdWFp16VvoKjHzNlaK0HAu4Qiq6udphToQTKjr0uy3BZ0HL1lm3wAXrSSV+f
BL0wWXUU37CJpAmx9RoKBY2q7t0dpaSsfG6hLxrc+YvFww0jeZQn0eiw4idwXzbd
LNOMNEgoci5BvSkhrikGkupiKgMZZHkikipZ+rY2subJeHEu69Un8k9j6iCekTWr
hmPgKzZuWXXI5ZNtfpwRa0qU3ztxbXY5IDdMnwk5ndiz6cD9EkPs0i31mphzOmpQ
bdHLMxgnLWT0zgpma9M3vA9JoPsWpTWalJRXixkU1xP+6ZTJoImseVvRo2DsdSU8
ClKtF+BROSvSQ4lcwcXC8Jko/744Xm+g3U/C1AbptUVhWg97GYOX3VSVaD31xrzS
umSRKW74ebekhQlPOlt7RykvfPeVp3bsAODhGfCHS0YvAhfizHe9pctr+CbTTJ8n
T2fjVvKNSeZeCkWga7hqqLXSGCGADWN3UxsUTe48rIPg0j5tpev936L7lphb6yKG
Jvo/kCT/QGs4e5slZJDXiOY0elE93GMFX/1I5vC95f42jtinECgVVdRBzj+ujDeO
g8yaJl+n0vYGxXFpIRLX1ZIqWYf+i3ErEFf9B2WrYCy+1Q7/yrbo1WM8MfO6agLh
ESRbHEguZHOEwyFYm+oNddf0Xcw4Uygr21BqaOfFD6MzqTxKcbUS07H2ROBK9OzM
HRo9pz8AYLodaYJGcf239kl5RtE1OrbLq2ZydTTDp2zej9uM0asHkrPN8mXiN9oK
KsiXuxbHauFDXOvLPCHnhuG3oZXq8TLyZQuE27YYEMP+eKKaLzq7mWUpgQSgeh04
bdSO0FWUQFjtJyNeVJTFV4+AgXkZRI5t082BM3QwvfcKoVwInV6AVMDSk4E2ccir
mdpgNM38lnB/TslYH+bvUACc1xeREK0yU1DFpSIYKY193kIML7qikBwHqGDlWVmg
qi/Kwlq82mObzZeLQR+uH0HaqiZmeXMJh1yVLz4CDC0vyJwGroSosa+YzN1KESu7
v+yB1/hOja44/oW+rVZjxfbhfwCHc7Cz5eF4aaeXWMPfZzI2g40LYXDemxk6iJVo
Rd2ES2jWjzCODXqeM8SgZF8hy52HEYaOUZxyHSf3UA/bkSHbLh3BrF+55COS1Slk
JxFQ9szp0I6+YcnGio4iM0bSPTw0KDoobvvu0YOjUcQdzfCe7iyBzcj2ysd08FoP
QkmHv/0U59schsmMlrei6USTCSzYcmsoQOhYGRbaCEVOC299Ov9/A2Loz3vHeIRw
L1IPKJFqi3819Pp7jBCyaDAOitHDEdxTE+/0zv3nZWLXoywQBSiwDpo3/4XsPjZi
LCVDdycasUDBNWweFEwS4W8h+r46nVc2eddQIt7VAYkiA/T1RX7McUPTAbV0w4Ow
RpZ8RU3SIK8miHwfVIHtuEMGeGQ7h83+0Gc0QH055zvjn56pl1XY/lSK5dqEXZSv
gQ8P/8ATX6II4K9mXQp6X0hWbnXsz39u7yJBlWsMxuBUyggebFvKa2k0OgYptqst
cZ+nceV6fkW4Dl/OpcIRDbwEB0/fruppRpI7xIZGnQnC2mvmbDcPBVNATykVb44p
4CuesHD1xljgTaJtoDifXoNJoMFrHDidn5jz37vWC191otplUUyDBkfrF9c3nndZ
7+Auklkfl79a95i1kp8cwouwpCco1FqfoGSuBOgrsC0QQCum2Smx+ImVcwCNmwAp
6FVtfvq3uW/KadxP5cjh2TrIetIw6oMHLOZSd45aDZAc5vnETkrwQzZByTNYh9/T
FoylORxKvCKKk2XbeKFQMaGKAtSr/u/BECbrg8xKSoFD9leeLwHjqsF5qXBpSkuR
L7tQJBrPSe0L9OSjFqzSvK7JzZaVB0q/NUGCALkWmbrqLZhuyC88+o+P//8FCsNt
ZTsRDFg4zqMXfZNKdFgHaQeXszR55KvuLH5b1Ddh+24sR6fs2X1RcccXrVJQ27/T
m1JMNi57DttYVaxKfAbb9YlhzM0JAQHL0kO4FP++hMByHJ7VT0lNmCVBWrZ0C2FK
oFrvG65XFM1sPzRUq95Hb9qBkIwx/CuF0Gu0SMXHHnMS7DnKEbjbOiBpBl00laVt
1pL+m2Oeb4hTBRyXMaNigk/bZkyU5gx5DK+oPSdHmgwNXQa/v8+7tiwC6SEB9OPM
/c+7ABlQHltVFu3FFKXFKkcVjTdhXRGfhOrjLe643oGmiR2BguMS54AnQB1tpesT
BLWRU4B8JI43Z6jkZv7ARy7cU62tmKiRrU1HG1708I6GrMExY/Mt9y7/nONEaCFs
o/MJDG56t9T1GTCMY6yOtXQK5jOfceWZBzu9a9WNRvvq8FUKHP9sn8p3O2nBn+LF
0fWA6LgpAHB6BOTdh2I2yGD9XdwEIZp2DBfoqALOXelgVxT1LJCTJyQ4kpKKTH7s
NPSBr3EEWc2UiZ+ffNee/gMayyunroe1lU4f4dKYwjDbkCErShgAp/iXrqE9ufOy
ywCnwKSj/CLuEIbEPJ7aRHYztJurqu+3pELGrwabAsF5XWrrKqnktjkcXXSThTtt
jDu0YJGfOCO4yQRL4vA1/OTffx1Q3RDdCkv2r1vkG7EHszoV5x6P4bxrp6mmzeSv
N0A8zcGOdslbzW2D99fz7LTt+FLlkmJgxAzi3kXhDjkv8wApgZfeFt6l5LmjIRFC
dzJi4K4ZMSsoLEN3Yysm9p7WugmW8XlrrbHfHlfYYkZErp0bMk4tmoAqTzjRP9L8
kg5meombn8+ZKaNWw4pbLQ3EKd2AT5N9wCr0Vk1nMxbUHcu/ajKiKudaRiIAFfLI
O4mITFb2Gw3l5WIORYKcG/TrS1MhDduSRs1XHt+MTyBFcC14cOZK9w/5Xn7xlACi
MQ1JeM8Hbhr8vd5hNsK0p6vkD7E5C75yYOMBNnMfo570oITDL53euQbav5FoLFNw
YogXdonTGSWSaGiy4Q4pfkH5xKpYoSy7OOMfW8KV3Cydp2dQyLx77uzXFiAK0gDW
Bp0UsAGvJvv5epMwKKamYPxSg2B2wAuYkTQaL5SpWkJ/4rU8sqbftnRhl40viVl+
D/W6G7ZKN4YfCjgGX3uNc+U2sOFBaRdRrx2rkLiAa2lcVkex+CBD/+QnOJoAv4+/
hEEIMfhMoR7KbY35+scUdGFQ61U3pk5oRt68h/CJHn1ME2VdSBxYwty5OKVrhi47
yzVmKmgQamqSLlno4ptB1cR+aLkih0bfKwcFYc9NSDtbCFwrqeCToEcthmBvRzjH
fPolpW4jaA2Q3fbny8KRsL8Vullsc8Qgwyc65QgncBBhgz8SFbSWtOtCwbathsfl
1IWoXDVwtLWwW4ogS3wM1I9uqvhesc9Xk3VAqj+yyPA8t22DfXCg0GFiN8oNtEk/
4VM0xlJ/uyt4JPZalFAoqyhiBGE+Zdtdkp1UUiq/gYAuTmFPC+VKpyLTiRNVkjdl
cTsRYlhvcSFduEFTC5O1zGSlemLHFBuSp9Vemqh21H9Z3xP+dFbLAmLWeYVb9ZaF
voZLhp2GUKjudo14wwZeE1GFAo0dr6RGQlSUORXcIFYhkBOrjE/CDdPUPd9FF6cH
Lk++K1pxvFcI5RbMDIvyyUp41QZJqvq1eBfEFdvFFp9RNMAUn2SSgy7AW/XvgLt5
sS0tt9X6j83yn9PMcZaTZpXIY0osEIuo3N+b05A85hHmn/rndEoFh92d4H1VjXaK
HurYAH2OpidwU+8HlINy2JOBrv9ABF+5nA37Q2d6MF/P/lHGYZqFNOyWVnxSurSs
cOQ/8IxfKotW1Z9edAEMuEYl08pHNcgmzkGHDy7saGkki/yqH++mm4B0XJ+LRnnZ
gPhjEvGeiL+2bOI2wFIvNYpq4e/tHCtFgS8oredEaeE2ixRzeyOMeASVhEJfquJB
9HEkHCHVI6HHEIlYrpDFYHvaPQp8CDHoApDp8RGsMwhUlxpdKgtZteV5iiRKFv8s
NR+4308c2/8x7BYajnDe6+Ys6MvWg2q8cmXKov4mgb9B8kRMM8w+wGc74XsdSE2P
SnXxRv5jZ8bbrZr3sqK5lCo+Hgs4lT3Co/1nqXmRTKAyEP9CEb1WOqeeI1rXFUQA
uVbhmAD+QCebFcFXM71/rRC2VhfSBOGZLFHxAkL5z70T+j/unMdG6RtfeQ3w0nPH
LTxBvuSik2gn8TcA+1mmQh3jotuz/NekKuj68Ak4A80u3toFu7hwuFLjtbBgqLQv
KuFi3i+qNUCw2Xll/aTWvENdp8rq6qKlJPDgUS/oLVN7/FhieGRcuSyWN394s91L
aXkJmkZWPpxFdQqDF0YaiJ82cJ8y9pFHKxdfn+JPl8tbY5Sv1Xy6hbifHWftcrTL
yeEUTlFR6ofHOyZK+VoNRZDO6PCECzrFk12VGv1VJAptmVwZHVpeDPzcWJsryFkR
RmNHJlhjvLi2a7gCN1JmM60rqj1ORJW4f4rf8Gzy35PWLDo4kS8gXdQDKjE/31Rs
vUZz9LzSUHeM7ULUNvGzFessFP03YDeVVQrrb37Qb5TjPOR2nv4mWez3sJTMQcSV
ZwpOLW/qj+9nJPSxVRfy+9EHvaDEA4JScXV/nj+35bNW+y+I4gZKn4us9CFEVpFs
NQvcq88skx0ap/uDL/O6x+HOZBT7HgsM0FtUjQmEKfcFpkDaUpXHWQp6wS2PJqy4
ErXBGSUaOkmWqk3j2fbSB6CoJp5AM6yO2HHDTWUvCWV5gD8Ei3FEzfXbalYrFxgs
dcBMnf9qGyHesOo/2QsQc/ybZOvgjk7Qa9oce7cs7kKwG37DAECMpF9hhJzM5H5u
OimNXRBV9Zilj9uYHtY/iVZlu3AYg/Om7q41J1/EI0ZGP132qTfofM6czlxnehJp
rPc4QOcb640+ZKqVb0qN9e1Jb1KjQbYy5Of7J2vpL9yi3D5of7HTYV1ztSdycg06
0+QLWXSznoirbW/KDtxlR90QMFZYUkOZFuQVcE56BYYSqLUAotPCL/uV1XhBh4YD
Mor36WmcphMlghpHXc5NtxNc1xAXQfH8j2vSDFF/xQJT7t2M/fa31u+v8I21kWEb
EiIYPbgeqb/ik17ge1bTF9J93aUp23ae0fAHFAt3B2c244arS7VV67GdqoG4wPl7
v2s82+yGaoHtdl8QmSIYLvpm6UMuWOrTSZNqSwxwXvjJVoI4D58W26NHasHtHEJJ
DqA2Z3+aMMlG0HboOPNR3gZKQe5ePOE0kmAIzpU/4U1X/9o3fSlqDO4cjB7+IM4g
ZjbQYCLZ1nste2pycKUfPaYUPJHSB4ZiAYvsTKAtvjyYNzoz9TipHBHBOwqrU4rp
CzDAkAdUUnXsG61izIwcPlelBDCiPsQP0hIoFNdJ6DBF5LqBFNIq8PGRUGt9PFqg
Vx6+ZZgBBineNlJuFOLEkg/1YvCIHCV4897rBrD7eekZwmrPil9L0b7IxamlohIm
pFEuiGAkCxwwI5Ntouzo1ZJOCl9u0qtKRBELkyNkwQCNliMmM4BzRv8911KPzq2Y
XQLh4FAAa+Tizz4uk6nlDgr9ZGaI49069Ndv9ly0umi/KKiJnBuqutjhBKNa5vcC
2yaeo7PZi0fzy6x/47e7W37Rm1urnOwvEt4JRRgKXNGne/LZ/GGuN29kcC54KtQJ
n7azsOplOLHbeFX9DtguHvg8fedimfnpXiK7QUGrpR1/QjVnEIJ58BrvGdl4qGQv
XygA4VExha7EPCjGPNUCsHQdIa7MYrmqzAVdDeP5YQR5wxrRjM3l4rj+NeWs4Kbr
rZqbSiROTOV8eW9bkJZMvbRvNOZu0gh6ybx84Tzjtck/kxHk5N+dTTVd6oGnNA8G
kDPM5+UMnxiaODvH5wbp/qRuuYR5MPmdyr+tB1nJ+Mlfq7sFG8sCaagvm/pz8M/h
NAeMTrC8qMQY2BY1r17y3SdIytkaJQYHApdv4119NZvQ/NFu4TR+KXK22UfILZtl
Z+evbuqvJ3rS1QYUL7XM6H+3OMegjbB/5xbaiYk2Ob4BNcSO/xzZ9B/hsOChwG+O
FX0LOakZq114pyMdH3/xCfKVcIvD8E1E3kgZtPO1bIgPj68QaAiSus+RbfzFnc5A
8sDSiWlpS1X1c/N1XnABEO3KweQquY2oXgcIpD0Q7lGbXHvSIHPmUvtP4nGZqZN4
QAaFCYTjS2l3BheXY0t1l7DKGHg4wcXZJ6F+7NNFdRivCsusWrBxSxRu9TfS7wl2
Nry7lga47psYfVInnsoewZQ4eIgaO/xlbIxF9a8vo9jIyANb63MNbtazrY9+AG1O
8CV3/l8XBCe4QrPLcKgjiskmNbhx/M7UTBOjWVQXZIsx/geQJx/U49PlFvleBP3U
0Ps3Snn4EjZGLd3wR7sSIoaq0salAgZDO4XFCwlv5xw64NC3MKCHgwekhdP6Io4h
VJbQVC/4lF+kScdffsi9KUOPl2pKMBiONpucvLO3dSX6fMd1OZJ1HqZFsa5RJ1rK
I3EOTtEUzWMhvCEBjRU2eecEIkb9YlGl9AEmg7V/0xsT573broOWynzG1+s7tRdD
cVenh6PUCEIg7HuJaC9wS3rbcOAwEbflBqw8C2lnln/9CCoSIOONc//W9slEyq71
6+JNWWvjOUEAcSx6rqStwTNEBQdhng/69v3zYtoAoCxNcyYkrJq7amv6qGiEfUMD
A6UMsGuBqIpXHjdxXxhHBLonWrktcElMyYp9/y1VW0I32xKhdTem0ZdcSmFq+D2e
EMq+ZFWGXlr5LpPfFyKUGzzW/ecAA0S1Ufor8qesZAQtmu7pbGwSiAdIOSGP6nYF
iqYA8jETRQBndxGUEkphnSkC092CpoxrJ6Y6C854GYQcjNPRXsl1xmA/GY213NX2
XSn4RWxu6Q5k6E8Aq58zjNaB+RIhH3dFGQbXvSyyLxCBrgrq9QQigIRkfQ+H3gol
Lnz8ycdo33BGh58hN6rgBHbO7R39JvYyUjOOCTBBtEhx4s/P5MELmEM66XI09nov
VrQINXCBuEOwHZ5FXHhnl0PsSUG2bhmN1LmQw8Cgsiln1eNqbQOs0PUMXdHKvmlx
I7e7nOla2FW+2SGuW7qsZvnBbGuVnn1H1hhs7Rjx1fsCS4fQRGyZwj9P/TlZIUEK
13R3ufrYceDuz91TMpdFSknWinse56aVbCqTtDQPBji4NTuvnNNFaX+og0jFeeNc
s9Oy2ja0crLU9LzCwnjR086ClwrGkMbpsFDNbFXxs58bwwy0CIMMywajVgtqSxKt
334o6vQu/PFtTf/7+epy2E5L6aoubPMmmiLr9GzkhkD/794DtD2zdsB27QUB8z/B
jNksQrwcSiYPUPTImlitgztUkI8R3hAtzi7EcfoRAWkIsaMGbgTy4dwLbrFEL+8u
YFN9vLGQGJPrWm78XJu7hQ2it/wT0EQDLqIhPlxRKR3bNAPJ0BdQRXAyASXmSgnL
U7rAi/qzDrFJ5kv9EDU9SZKzDALkm1T7i7nD8OCvel9h81AGcnggMN9xpF1hgJKM
oJGBO2k+nP3KatDgClISP8tofSrscfCV7Zd7LOyazZIbvbOjeEVVFQxF85iMYkpS
r+Ze+l7VTiwo2we8qP1Vh0BIb+0nwWyTKggiGXTpI4pnU1Ytq6mFCjVoKqT16ygj
jXj2gkhQBR6I9wszvkXrZyqUfj50C865+heII9HG65lCFXijm7RSlD43r8jKHkoz
a1wqsKFO/2jRMf44iaYYPS47krGosreDA06Zv6Hq5n41ZlRYy0cLSjNq4kb5LNo/
rUiESjsQ4qfy2ldBWcbENiiAqAIe8OF++l93PZlwlKpo/UWaa/wEQ9QCV9lPooG2
XqDRdShqyV0k7Fy71f8TeWf/nvLR1IMi6Xf63AEz5GlIEtpnHLsWme6eb0wm/Fey
j384szM970pWDjPC8CcB0ohFEWK+iO/2NtQCFCVhpeLyeZAcSB/0knZN2HlE6IrZ
k/Ko1CT72WqFE2opOeYluw/VEg8GDBpUTcqEwPM8NbfclKS77jHwYTEj7G0c3iV5
gChWtZUIOmjbE7AIQtYcMNJFXexqsW2qzTokcyo54Ats2wcrzxKbpRDOrzxmwKmW
/nwyM4aMBkjHkCxSbsq/iplqD6lsVQKEZpe4uMViWZTMIxuUtnR6a64W4IIf4Oix
xJm3qKTTYcMyo+Esf9s4N0rdgm8B+CTbDEVh/0VIz6M0BxdLRoai4PGXxj68DmAR
DBNHMkkdXVhq0qfHNJ4vkDaSvT2b2ZvB4FDl1cLQuwBetfEJZK6L5a5DW/CPh+hj
/0Q8Uxe5qZHME/JxN8X+gK3Ds8GIPWM5uOKjSu161GvzNO8vci25HzZr3pVe1nH9
vQkKeXKFT/ZXDKLdcyKzX62KGAt0XRyYL5ovIhOCrTttHHKpRRovN5xLcBZRH+AD
8vn+qZKS34V33XgtPro1RnpoENwoQgTtKbRVHpu6kI1ii6V5SHafqyJX6foPiahn
gWfBgBu6rIK1JN7rC0OG8MegS4z4LnaN8WM1QHE8/F5g+G2jZyWCt+4zBLwuOUqo
eifYDwqPUYU3kNi/zHRII4GpK9kG7gWR3PmFcGYSjga6FIJ7Zw1iL3+k9esz8OJG
JQPjONoMPPJq8HoX1VvhB4lkvugJDi8pMPEmE2eGct921pO0n1WpmjdkN27kqWa9
6XYSUmp7R47JHR6rthNTl+wKq5hxZ6MbBcu2OMdyQKQVFgM1oiOZRtqCweN8TwuN
YPDTZM5Kl5mfc6pHJaEyfYhR3Qmva9sRzWprGPUggQpif9v02Ga7xHpf2fw17i4c
GEhP1CchooQlA5quvxNW0zDpdzdQt95noBqmoWZOIPbKn/sgR3+8A9sRJzIVAxWt
JFmDfUgadDTWEFhJT48I2DRyjzfwOzPQ6OayhrsaOkyRWPMJvEwsLav5hUNlHfId
25xg3ExbzWuNL5LhjkXHITTEHG01b17CR2nCLK1engR3Qk6on6KNOfLOqkGNnywm
wxEP6O/lfZuMW28RBUhypbwNRdCywTwZu8HklxA3+B/12BJVhQiBCLAAJvFBwVh0
CoHkLXIHxER2AGE9DF62Kci1UEiArt4fsqL1Pb6Qgs//dYCBuCpv3oHTCc2Nf0C9
s33qfq5lrqJJc68SAYFUJ6zeINzZm6jFumr8E+TjMZL6s8uDZ4ODCvufbtH3qMoK
TuBIyRtEImV/lPRJ3AxTsNJ/XMZEWOnS0llU3lwZLDT50DB4R+LmVZq21gDh+Bkn
GHj80zMNeHBpNi3aNxPml8wFgYGxJiUopoJ2woxicQhuJEKO2zlELmu4CUYIKsee
FWUkm5HODEbL4XA7+FglXRNgjWQDyjn1v0gZiALeltpcHUhIAgIlp9j8JaA5Fvru
QfpMpJZPOZH4wJiUXPxbCZSwHzVx9utvgzjLX6YcDbo1QANaFFYMUfTimFVLvGe/
BxVmTWvoaybNhcW+r+m2cfWV3gLtHoFahxPlsIXlBEVPZXMHiswtV0LlSPjIHnbW
fl8xGm/NpU15qCg9X37ATzszTOx5TP15U50GmtjIVqoeXgLdJ929OZ+Drm1TB1yP
Zn1++QQQC6Mv8ChQiLP/vCbXsAFSuXf88mlGUWdmanqqy68mJqRvhjPAlRzYNa2i
rgPvkgM0uPyct37hQkVBD5kQ4aWnbPjhg/ioJCp4qJlqljp7x/GZkBp2+tM+qBky
fYOiPswges0u/2zdJ4Q7WQvEfFCfVxBwZ58EkwGak3FTiR18ID/otKV96CABgZFb
zwhG78f5zwCLdHR0g0dZe99stdqbYqH/DGvSG3sgmAg0jrNIp3Ps9TzoydlnrOrQ
+Rrq1nK5ML/E2k40ZAJedE53fqD9Rl5lO4gph5mWH4JCNiOyJylkkWjbyGXxOJSj
ifabvuhy4cSmr0i3Fh79jwY6S6P4Wyw+hPnLP0bJsN9VvvQw0pj0SnHfrcJ4yn7l
fgUJSfYv3YenW0wrUtjK7/0zhvM7i8T709mPDlDmKZlGidCDKdVwIbYUzUdc++zY
oAdndh7fZ9vFPnT0sGblT7d9jn6vXxm7NMVdA3zvPXXyvMx5+yDqNXLCPa1L3Anl
4NDMIs1qsWwXBrfhiWq5uGR8dD0x//cgUKaOZvtnyq7JKHcwyNi/a9TKVKLp2BNY
FGQjUfZDElvMVO2bI7QafysxMjI1u0uMB5gC43+j4uXuCHAIQig8WGWDtzSHsihA
YFL3Jcb3+5ShHeKP8/0HnF3qGUHlmVsJRiEOpYh98gpUeIghF0DpH3xWG7b2pelz
62rZlRDLrf6Op9SCrefC4/xJCscA3ZNW1niZz1uqPUSmFvNl3YTmajJfZQnkVfKz
9vUqzwYI5is2P+mXrilbANZzyyAB5vhkQu9HdOXO6YGQ8iWF3SHL0A7G4Dj2E2us
VpvVhHaqJ4c0xlcTKAIXsNxNfVHmEcZmL7RSaCTkmiSgqD8Uu1L7L6i3LiV0TjIK
J5l0+4KB6y+YmEdKMnJOAapQ4s1Fhx6deJ94e0fLv+a08ISqNOqnqLatqKES5eXI
UZmlyycUlPPOzm3k1mMQZ351CaWVOFXtcmvv34qh2vz97g6vF+AytN7D/HVaQOdg
3sLIszIBGse7MRMjRTVO1D4WVMWpFKSH3J/PE3YgjiWJQBqV/W1QQLOGYf73S7Mu
nu17c6wQ7sJRkgJTyxmG94J3vyTXXJBesSghzK13u4g9op8B1mzLO7q/GByVtmOC
Fhp6R4Si7Z/YWmfy+ii7/mXgHFVBblvTYOZz9bZtt9fywzzEWKcmQ+fZFHRk9yv9
XLIERyrKtzshD4htU5UxRT4VwprGeI+4xFrPlkhB24ZuzMeoHPt+UfdWA6ZS+iT0
rCh9vybpCRqTv0sMZUD7af5cNMnfudypxA06ul71uvHLd2NS6QBfKclwRpw1hJBP
d39xBZKMiLSlOUoj0pO7FZivX7KmXsSug4TuVlh/I6KwT9/Tsv3zvedn3q0POMWz
LmIizWd0c39/Bh/9nZGYA1khNPcFgZYQqr+E5RgZ2QhT7CM5lzzNaYSr8iq6ALDm
QAul6M0jijgRt8OwJu85d+vpDi1FYXVll9JIlpnAcQx1OuPYnb231QAPKCRgmXoB
gf1FHJmaoOdQGzlq3WiNpqWEOYiwzFxN8lvJJRnq2tM1FhlR9GdByWa5XMh2p7Kt
jf4EU3vZLHrZAuOXHRS6ksz9K8jRzD2cMM6sMF6xUNSA2HY6grA4wAQDS911GzSi
cf/xJNB4bluiwPynOduMeMdv2TuitFbn4PS/lctXTLm4wsf94H8pqWUYyeU7c/D6
jbUenzOOWX0jFrsVUMpJ64lhWAnn1NYcIb/PenOqu2LqNSVWk0GYcSVMgFc8duGm
zFrcEjHwLEIFL8teRyhCmX0Quam7zwdTLDMNgO3C306lipC7RGXIb6WvWsPfCQy0
JSqzeiyqZ5jQRTOmPT7Er67ovikmh+JOCEocqA6fjXuzaTVaS83WfTi1se4eGAmM
0IfiP8Y451nydrt4OldxQjirtc5Bh36LAaXGuLvW7899G6LzyJL1W0Ksv9LBnPGw
05KoUHaw78pvRimYVUOkbTo0kCqdA/4XqNO5mvMvtgQkkk7csmUovxVq5onDvI4C
u+ClfQEjTgGpaobWRn4ybOcmhOOVAnIhb/EYXQzzDYXOm/xrASNB4ykQtDAXXY4l
UgvAUKjKGYeaunLjUpH5NHkYEBCTzL68+Z+TYCdoUs0/ewMOwdwWXhy6SsDLYeqD
WeD7hdGd/h5eE24kezkBmRRT6/fJX6JymMpkCvbXvYeinf4a5VC9V/5jBw+jLZ1P
9YfYj/baaIQQmg+qxuJ9ytizE/4qv/Jd5vCtjh2vyLQeLkCQgxDSjn3DyEsAMoYy
RoBhJO4Y9Yb+Ad0uH5ZxbJWAhP0mYm42cyREQz25fWYneYHvXxKVs1RCEkZaOgkt
k5kE3TR8YXNJehAndhqGbANlmdEzZxC6I4T1FC4BsGzR/aY9XG9Vy2c1d2Nt94nI
fqoAWMucBYqMdECTmfMlom3wJ9q2vy+A9+w6drqSlVibIDQVAlqpPmYsgbKXjcNh
PXqy70w5mJfaz78n1u794YSTOBCz0yv00oHv053yyl9F0JdI58vtDxjCBq+Uqs2m
TO1Z2TUfnRd1o+TApingJsuFOb2c15ppGp0TYb6j+zpPz/cy9SOhZiWj09z9dZaf
9R8jNjsLTL4r4xgUI3q/AejKp8xTLQ4u7XdTPsPJjefWVNDLWtQMt8eB+f0G9Esx
wf0E/Ofsnr4cv1edbwZoYCVVHITveg8CvlYl/Gp7d0jkQXEitx9Mv+rI0I9XX5Tw
Tf3fBJ539Jq26vzXjdBoSY32aISGjj64OuqGykK6MEF0XIn2clrfZLMIAGNBsBY1
4JhGexCsdQNuZ0DiJ55VvPYMZGvVVdC8sPw0E48seyWxYyGGfNiw7lLY6V5s2daJ
FUSNaQOimZS6cXmZmvbGXMEn0OQ+WdjZzvC/qPQb9T8nQFhxCqkriFfzFUfEHqx+
iJrHAHIB6ryz15xq5Wx3AiCZq4UeESAhArjn5bNVEXn4teDsBh+OUZo4oR7/RLNR
MbpTBOdQq/nyGRzoKD8blgtsdNW+niwl+MXaFQ0wQOEfzO02HxKwIBwyU1tlObVF
gpoLaSlYyRGb7IYZfrG3dIJvooJt+oKs8XSrMhKp1rjOwcuRFxaaMW1OQD+YgRaj
ZfD55lLdduiAxkGnsvlxirZilY++fr5MOZon8faTfTC7/k5sU8UIr6meeprwKoGO
Pq4a1PoYZx/C/pTNNlSRshP1uptAsyPEiFFNdFJVNoVoV6zzoHbDcJiYqEp/AWEU
j7sfKbod3KpB4dNxSwph6sozJR5Z9iM8R+V4p7Mh2CVbkmJUgMBB7OnzP+lOG868
dQ9IuMljnZi7qCafOX6uRgfwV3pANl+FY8xbZxThe1aIYbKCvzYRMLNcBSMR8i1C
n2W6yB32DZs2J9yu1vAjBLmR+sQglj4xjSK9XVMetZSaS5Xa+VvGKYq96veHNI0+
pKUyeJc3qhSQyxXW/AJKGxoIG5Kvjw8+7T0n0zhV9mGOkcYT4vONyrKnxUvGQsBf
WTDPadASNLIJKsLTBKuEii4md5LYneFOaRW+a42AorprRHE5QikFE8xGZHECd6ci
6c6Rc9QYWcivI9DLs+TPtjgtwXFHQjlg0Dnls1Q31AOf8oIlS8WJAnNUvkhLMCri
f6udMtGTe1/rDfBhFjgNnb54eni3rbIpbTnm6UuZAD2gBooKruwpAqZF2eY8wqEZ
LqJUe48ELsIc+jQMmlWvxZHFulTxcEtR+CbJVuSYfBTaPYYp1ZbbP6P0/j9aiPok
SnMv/n8ILTdRwTzxpg+gyfUvJ2q/w1kky0XK8OrHUVVtHUNESROlv8yRqWnS7RmM
quSVxMep3/GUq1sLIYQMlU2LZFyB2JxT94cjAkLItgDaSxtZpIs6PR7rTOJLAXMP
KfmnfbGXe6QVVsoOxuBjiuA9Ox8MBUU49STJoSrMIWg9oH6GJR0zATsTvC/CZRBq
kgr45daG5njMEtFbYBrH8dDYxtO0kJzJfKp7/uiP99XV/sdIyR16VeRSDN0Ancza
YKCWIns9wIjWYinUlgnYhuFt1ZUFjIj8QwRe5W63UGj3avWnTXckAWe/SGXQcN3A
bCbB4yclHI+Wlm+Xo6uaW03hlLjJ1uygACgfxJQnqagb+yRaQ7zLuDVPvLlYvwHF
aeVPEHyLypWrUDRCGOEwBOI2jx/1E2jgJKvzzRfnprpLGYhJr1zGFh5UaZ6Qt007
CqIENzZkw7pMp5MJaBYHttVGDZ5UaSNuAqmxrMJ9uIdEelx/hPUSTpvZhlnULuoM
L/Lx96UTw8gQvmLgQ8Oh8iV87M6hjgSUInRNxrCH9PqXuh34+HS9NkkBKqmJj7Ko
gNwZLvs2l9OTT+b67k6YC/Ijh7fh7UkX18RnE6Al4JmFLv2aiYx/CZbpGD4kv0MB
XcqAtsPXx7n70HImKuqr8Ep9v4DEH/tGj+29uN0cCdRDPzNCYsscmwi0pgDsGiDZ
zljH2HSV6cQ3mjJCKlK/R3NsH45H+9VUcsKYs0UfoQ2Izm9MxeDtj69HcYcOiv9U
t4L2Y8gNChSyOYolxSmU2KqxYY7X5uXCdyM+9VAIESz1OIaJeNWeqUQlerVthGuJ
YpgFrKmkpbcqzP1YX7mavyIlDJOLDtckxyQ3klsqkFf1ntYUQRg+q7A3zESchhPd
aqYmlQj7iq/y7XviLcOPpexqdroiqOXQhyMnhjnGwU99p7aLK2d9ncB+sHz+AzlP
yRrorLAkMiFDcQ6b+NLNodwhW4Yd44hSiKTHBCEKFK/vOZ8Qjji+0yd5HMXne3S3
u+RZ9yZh0nvodbg2AZq5O9IuiC1tlipD1Wa+lVMBRPBCiCdi1Cr4mbdD+aT1EHIc
Vba5Y1gCaAoSKaFgyHbCrpCijupR0bgRRsxv8dWENnlh2H0+cm8mVYSzCxD8YNwv
LQc0SXGWftbT/rM+E1sSVTpWMF0n++k2ndfBQzkErLxupOoxR/yeuMZPtZudalNv
BVGu3vlAmfEjoRu66Zvtj50T1P5Qb2OdNjzVzWD3HyJWXrHWKz9IX4JdtCD640yj
60bB3+iOysSo7mifLAH5sLWG12uSvHN//wcjaUK00mn81cNZDbfH2xHnD689JvXK
Ln31BQg4TLapM2G4OvWruWgjjOrBug+a0lC3U9el8XNwjTAItKTsqbh6KgBwty+Z
aLBya6C5CjWAOqhMxYT+7bg5HG+Sn5oKDyM7QIECyHfDUtXs7xTdKoNDqhKgXesi
kYC+dQfnbjgEmm211irYSVi0LlqTK9EV8wTuQJSwNg7uP2DAl3QUjwMgSOBmU7yK
XWrvKCKwTcPSgFr6i8lrUcF2bjKNragOECK/86EoyBaucII112hahilrZgnq0Ga+
SBTkoVQN/LybzDHtZC6Q+YlHsG20mooKFdL4JLG+a21mVBPBSmMM0Uh3ChTjadGT
8OtFU/ZqjJGbeufRR70RUq7hyiJTngb79/kh08eGcGWWtoXhvl/mLBrIaxYls4qx
Z1S9VRuBJsENBaU9qy1+5fi10wF5SbA+HdAfY3ARNpczcuETayqt4KSfJWEw09fB
0/U8h+bBLfKHRq+Pat7/BqxYkRSFVmJ4I7yqfUqQejB4QRp2fwV/7fmBunHp4btU
n1glpXak6eNQdgnMneioJTXen3fEu+M2FsCF3LahLOFgYGOUthLnFPBW2HL2bzTO
C9oYDay6SQzb1PBpdItCzJWbzjoOKTVBwPHEUOmajoxdlLglDXR5qIHr5XMVco7m
rHtmXfQSWcV3WbKoARd8vYrnyBe32EL+K3DHOqB5nX1omNDCBBhlj8p939hj2N4l
etFtNUqsH25jISK4GfsTBEOLp6K0iXJ3Ae6j3Xr5sJU3CPwVYVsxB7Ztb/ydPv7N
em4coo7ch1LcmSAJzuIfhr4AO9aU32/a1P6tBkRGWZned5B7GcnTtF6r2QNa4R3c
dhKHZ0hETwadJOF7NSgw1tPNVi7snQHE3rfpvgE2z1wtUyayG/+iUoTRO3sZkzp9
4y0LUrPjeWIuWJzmwXrF7xBXu5Wh2PW9xi/GjZTThajKv4rR/ZqMzR16Pof/k2va
PBPA93Evj6G9xYluEsjGQqtAbK0Ah//PkpBncR44BAtCTOla2b9NOoOpYRJWYKWZ
PYxmB/afEbvcl/M+q+XgE1RFO7Su9yj1R0vPKgXhwIPIM4vbMO2Ld3/aezIRMqnt
bEYQiYgnUzFGJUh0MCfZRaHmF5u+ZAgJy8sJzXszRHoaEZwF9iYbvrxC866FiSuH
445O2BOvMUSbwspb3QkaEXmHdxAIDA2qBYot3jVeQCBe7hngos6WPO7WCeyDr1Uz
SdShqwgci44isy4z0fXx7Tdp+zNbVu+CPJrtFRb52xhEExrmBg6WOkdD445w726e
0VuXrnYouGrWAqqLwnh96BZMH7FVzzsr9eTwY9Lsd2EtMl3EAxHL6o96rZstFqnQ
bEvKnlhnuBx0YEAJ7X3JAvm56pDtthpb7V8Ei+YRsUvwpCiuCr9lqAanOfPb4nq5
UsW0QC9BZYPnBPJQdSUUSkT7vT0XgCFYjMxp/xmL0QTLw2Aj9Fb4vZhvxmb00hMF
xk7S/rsnjQdNo4JKURuCSBFiLiZsvBCctA4ZqacTbFVASGeYeAA1H3ybHNr8LYhs
/xgMK3cHVBhiwBS6Dv9lwBCtzrsRcsgjERhQtPBN3t+KRZd4Ys7dv/FVc7drB5Cq
wIZMTXhcOrDFnebff2NadqkU+qRU9zZKmiSSlfMPMplk3hPCiKDMdy+CRyL9OzPr
xq1L86fzmwsOBJxxNclWiemQ/EZlXFrLisbzDRxoi0davzehB4SQN0IGQKp/kDB4
WfpAQXraGVbvRUZn6Oye4z5E6aplfIwkyXDQX4N0zURVh0x9WgGNaf1Pyf2y0tSV
oZyagKDl/lbTzQhA4AQ1FueGoTUapt8+9P5N5888vtdrW6GFjDs9ut3sVq8VJuRD
HlYLmhhxggH4xS/KHUir1mlgeMS/1pURf0rCWJVV+ynwVgpFr+BKqO5TRB4O4LYQ
spm+WlN3n4vR9QMX8sJ0GIGce88R6ufMILBCy2lmufEQuopFgVSwerowsNSHpM1c
/66iieC+eJlxWUnOZuCLX9p5XeOIsiSRJ82anUvnvMxb9sDHMRgh6wRsRy27c6oG
JuwscVf+Rq3A5eb1HdF8FqPpXc0wMCzncgFQ8LsRxXG9HuJTQSXfcp1J7Iw210sO
tTu5EusYMEznbk+r0ucOR1gAqFRx0lr1E1orS7Mw0wOEEdXHXCLCc0eow26RLjtG
2UumSvpQMHQyPvI1kzpnzroBzAtwhExPmQ0tgKz39Y13x7ILaTVXLBu3U0PTwPP8
KSIj94vDoym60U/xre7M/JKJmj71WiC8WJPQWMeDwDRxur9wXPsl0rnzmbD9IPTJ
O3kyAPtTb28FCdMoUonAFuBcy9hwzVQnGrV3APUOanjRQxGwIFhJzZCX7bowGAyH
9RS/aSx5lmyGxGsQyW0zMtF3i++zXHoToDPv1Bw5RJ9tZK2fSunKRonzdR12Jz+P
fRXAWca3TcmUDIEya/+uoSJiczSzgUC3Au/qLd3KIgXJNcYthJAMtfor4QdqzmoX
`protect end_protected