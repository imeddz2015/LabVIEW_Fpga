`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 13008 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/9huKRhRMtvnNqb3Z+UU7TahEoHV+T8U3P3ufru7l1O
3DlgtZzb9QxCbOjthp9+wDkjygH0eUfDrEl1ovhZG61E/ULyjJR2qqSbnFkazFzZ
96dgd171ppCCeY2OCHgDW132rNxVjRGLGSBmuTLAFHIUac9Xnhn2Dj8pjDzzx7fd
7tNGZdQJv78MY4T6GkoT0ltqfj9YKStJw0DhgMPMfwfbHuciRXVV8dkMN1t4e7Bf
b9AreISYw+T0kbu+8U0pMHhVdcpyqFwbcvoMUKVRF6/srzofu6tqVAkls656m9PB
XZG8M4vOMRbhe8zIDbtyHa2ymVwIs6lTC5Y76lzfHxXor0lqXY7XZt8A41OQvFb3
midMKX8DBRwPOFaRhM+0tzhez/HGUe8LGvRaCU23ePOhErmtu7wiWa/8g8257FPF
YcLceHKcoME43c7o+woMnSAYvxEfM7dgNjsCP8mRT5KFUZ1DJ9kdPxs4cd3cCr10
c9W9I2QR63ke661KFUt35OeQXHd0giLAgZSGZQBOW4A8g6hylLS6GWOzZ5w40hXU
w8shC5zhaeDzwPyhOEYtNZW40Lz+ujMCpC6wzyDHEWj8kOB/pOvBOtlFaspyGFJ5
NeReIswSElGQV3h/nxvEg7+7cR1q5/2M2LACB0H0ZGXeD52ft/N7pcXFzUSFx8ax
8D4hr8Gc5pNw4Ef1xPS6n+KzCHuB1LOyGardpxDtCT3EOQRuzQfFIcmKup54C8XG
MWcJi3ZqKZ5e4xJbzyS1teyJvFlVwxcu1LIc4IToZYTVg4DD6CmG/iqM87NnEg82
D+tmUCkDDD0Qa7q6kWOzb+VeXLOqZfIEmvG5cKRyih8jj+6g0z1IsUW/aZIstdsL
ODqQ6B93HACcAF7lOED67lrHKALrnetGSC+VUDPLxruFMeF4oQ/Ga7NSyDtE5vwU
c1jxyKCc2UGRHyzeMkumF0Lb9Wp/lIVNgP9f2Xyq5SJn74iCLfA+Vzh/qvY8LwlA
bQnUio6afFFSprS2lE6gRtqyGuBFz+NnCJ6g6Gnw07SWsObb2hudxlGf68RH68J1
mHteK9fiwyC+msHPmYSNDNf06/hY87JSB3HlK789FtsRZXgZImoYJsnR+427naPQ
oZiIsYpU5qK5oCzp+eLwiFaSgA/j6x5HS/UpGU0+fZsErgCxCv5BSLuRXIFYm8Dm
Z79odId/sCtN7kmSLsZypJKMXs8u6/oVU+KKig1w5bePo921NlgFJyLBbQcBMhOg
T1v4wXPu1XlkusFRHphisFsV4ko/WETcKYgh8QZBUZd0ywgkN5aXpz14lHurq07m
yZeJ3eDaBQKAdPyo2gDciLhbWQXcQbP7TZL6/00KFTbFGT/tTM9cHM78QZYx4kwO
m6X8pyGQju2mmsBWosPkfuEaw7mpea0I2swfHe01CoItpJDesu8cdKfYvnCKFu2x
DJD7+2d+FIcrC6ktu5vPux7FBmLZVcMj4oh6W3RwNucVXDtF0c1Je8bYSCiHo8TK
uQCpTDh10o/tyORrsYaOzR2R7SAK8b7ILkYb0rc6x1ErKiqiZMN1W8WAECFuWkLw
9RWizWq0OGfQELdYGf4koK0bhnCnrZRqlor9djvylCM6hgn8XDD/5XigR7S9y47D
IsabTZEUIVvdE1vjPh/lkFwoJmKp4i60QFiur+n5YDzSSHMv22Zx+0K1CHqvcU5H
BfEMcXFLI1m5OEhLN0ke3ksfLtC8bNs7hmJulHGAi6axRAwuU2Xa7Q/AvJpQ9lBb
JCJHIvhqoPBXkx7GOsj/XPmtkQEG+PhtUOj2gM0NbLCyQhe8/dF0TiSqe7soBtM4
o7LQogwUcN5KH+FCOSM6HQRdmBTI/Vlou7AqFlVogZiNh+3BruPUKWlXck3lgaLZ
z/nRPb7JNdV5V3a4szHBnTZ4MbQ+CTx45bpBlsXTcuvwp8UfXSxAgYiaJI9mrowf
S012r+OAGZuO3C/WTJBWNM+2sh8cU99lxlf4iXvPSWl1xi7UQklRLb39fGubkTdM
BwdJCsFc2uILlyOZ7TuWGs5QwFg2Zj+WZTCMqLN4IYad0q+wNTfr6sRmDRD//DEF
2cnO12yWUGfBvQ9DgRGOnR1cMiaUxfLrdfGb0Am9NSHRoEtWrq4s5TQ7mmvH9kXL
pxmmjbYTkRrg8RxehSstcyZ/lEVzHm+NyzZR3dvwV2KyneIXYEulffN11GIHwfg1
0L5L0z0gZ/alrfoEBo6/xZY1JLr38S0Yw3HaCzpxGEim6qZmqwHqJME/zF3P46/a
j4SMcSPkbTfkcz42NbifcuJTW2CfNVbPsMBi44G6Ei1Ojs1OmN0Huv6skWGSYpeA
ze9Z9whNKnjNO3o+zJXFJs1MOz82/Ld96DNwDhEAWUbHT5Gc8opltvXvY07ShR5e
wrVaaits+LlCuOiAngAnrfqhnkDUXXgUpGmX2YAmKGci+/Qpe2qh44aSUXsDQQNv
DKxMbl3pcLBd8g/0U0YAj6krQwtk48um0fx6N2mL0hMb0Y0zGuhryV0if5IO9Cnu
DDD49+kxHTwauUXdHNboyLPPE7eemSxVNDzCiTFzui8p5ubgjelmYnJrYSihAdQX
Suez+mrvl7pDhEpHRQ1XlfcbHcXE0pNe2HNe0JAW/xEL9j3+7/GWdR51yjgu5kvD
v/wIt0LXd6LqJP5MEHY2vVqcXRmPrrJ6Ra/7eCaMITNDT5IfWVM0fBYZ+0FsKDak
DqMVxuqoqvoyggDVSzE4sKKnVUwi3NHBV2AXaXFrux+q1JwqADKRBhSwPmgEZl8P
eKZnRBHIjzsjqR1/oks51hpTuWHcp7kPSKTj9Yq4phzdv8dPprRbd06ojU6S+483
AjTIH1ln0i+/WVfT5wPjGQy9tCOYXMyKq3KpDvbsabbra2KKtZXdNqIi02jFi9cu
FpMkdoispPPuUMbR4gxnP8RIyH923/wlHAYa529GMaX9xVOGdVALnrAsS9F5/tAV
oMgzWhocjaoW1dg7Jfk1HCr1OSofmcXNyhJQvLG6ZDwL08HbuPanEP2rMhu0HlF1
PARPccsaxq5IxqQsjcMZrqrV7XVb5Jnuz46pnoe4CE26Vc4KbhtbqpEYDhISIKvC
YwnOOML9uBgqbG4A5pzLYbSp1eIVKzGPU5twDPhi9UsQEcXgZqfaGSW4vOI8VcJa
FZ5LrkCZw/9xC6zdLPkk0gC+K/Fj/lnIHyl3O08NC3r8lFpjkDJPzex8sr7Hqxhu
8G/9JBACLWSQOqOah7fxnTbv9Hy2PB2aRwN4hBLTuwTygflQOIMfLxtMDVWtOQl8
L5HddWKpeGCDswawwmbFeMvXhAgK1Lt8K7RoddiyqqCTGgHy7CaRjp/RYW+tLHSx
2vsX5cIE/Fr0eG7QxNSkjPFfrn8KiTWrQyNRu+GrFKfkCn3UgnESN9StGDt/S40S
SdrGe8B/1xTJL+ShncsGECZgWohmafScuGlCsfQDNf6PzNeo7RLbrWUZbZSPINPm
w1Z6z51pnfXepFVpAdz+H1pRD8DKxlZGfgcSrTmPMIV+cBqH1EMvPApE+y3RB685
uSlMHOHGdMoRotzdLki2Qa6SQT6Vtolv26XdMhpKVyHNUUjjh24t2oSy5XIU34ni
/YlRjhItQnU2jYOkZgTcyCVBvP+z7qCAcWNGLzPuYf7DjLFTY864sRxcUMw9TFtH
KNTFZ7ZsIQ/6NhU4a4yrtnsW+ylBrfsDKwRVTgI4y5IbJ/cF/GFJZWh2wbee0CGb
P5sDOtXoE1ew3PD76V1WQhLTOKffE6j5Qd/QhzJ+kSwX0tVcriec81I9FtAjQUhi
OzhScYKFgS9eeqGuermEuqo4Oo2oDOuA+TkAbukau5v4PGD+H4MTZijvTuBnYU0I
eHkXdoms9XJhi7U07f5J2ga1r/iZOi3WvuRzvYyfeIoFpGtgmlqVMeFcgtdoW1BL
2SxRLywnwbzOaikuT5I86GEzZjCofIFd+VNe9ZaghAzBp4gm38IQj4n3zjpikfjH
6cA/eHbwnGvvFfwntBh1tnOGRhvKf9bLdk51t+ozbKlYf/lAPhJHoQ19lteCNNid
yxYAQBLh5ao4aoCvHorSF5BK6wsTudwsdtjRu5u6laXBlsqy0yUg2PXi/byoiUUN
KK1AYCGTfTGixrjbx6C/yOSn+F2vGsiR2DvktmhElFyPmPsPkDQTvzNpHeepPTWi
rQrn9GJ9ZGWe0c1a+UNk7++jlmZSsOlMmHNh/aoMtiRY/8+1aL0eysJ9+1usB+zK
WC0AGw6EAcgizxfRGWF0bj2a9ynrC13AtKbS7GOF27M9vEgs/Sk1aY2DnTCMmuKW
D8Ou/Jy5hBfe0DtGZIm9p6hFOXzQbgr2ECmy1w+1hv2YCY9YZETOOYcB59PYAbye
03eTbN0eC8xvyE112trSl4WphveBB8smb07smQk3aNdhsLl+mZvjM8H0pLOq59/j
WMbt1okjixhMTpxFZfUaP0O5lCGDiw4HxnuCJgbLBOniirl5XKH8TO5tOyOc5H9J
ah2acNIUPtPdXJXSd47yblYoQwbrQLp7hoTLTihtVMGh2nQboiWpOYXHpYB7+jap
ZUGcD3fXJ4IyOsCuUa6FI0zVHN4cytGdiWE+of3ZsN7MV7j2IGnz4dq8bEf/8j30
79yySCkihIz9Wf6RLYDRl0UnLm0QgTLwbikvrtb0B/NLvWGYDCGLXphAUYNQGNOT
TVglR42yxj++cEbQF3Ii1pePTbyEbmoxv9ErI6NnNOuKEc80GfHckC2YvTCAPRkP
EG4jveUGHOg3wcA/ahUzBtC8zQUlWoXSdncwoQyT4z3FpPasowrj8h+gi8yLpuHR
C2nnr7woBmlTHZLoMtDSFC1zOIp/zoafEIv6+gPlzBwUWmjWRu4GtKCEt5ujGpjf
sEvFxm46yQXOIzraIUk62v6n+Lb7hJnVvmK5LAJQsYkO9M7tz++fbS6PH7/Dsbfo
PtIm28EL6fH6B9TYopLF6FRaMacbjUV3obJZpXRIA/WW4O2n2QeJpTy2wvPBJX6X
vsgfC6mD8BYhXP1xln7YuGylsegILfJP+OIqf4csekr1Ksnzi2PObbY9dJIHxbRg
nfSzq+la9Dw3YLRKHV4NJCYi31Rrm1GZP8SxIu2tyJyU6ex+6UAdbccjdPF9hivn
gtUxCikHu14geNPV5hirEQXPCfL+MPsn0mABeyG4dloQCx8/VAxMuBGQpauJMeZD
8Ar/euyso0xEtAoigamLOx3WEFPeIHetg076FDfF0z3bKru5Foak8pdLX3GTBUNd
iom4PeBNsQDXcRuzjBpw1I88OARhkBabU+EUGd6crTzOSZPNBTdTyYbGIN4f81w1
UTBb7x0IxJKsgOvgE0jz9mhPdfxOM04GvrhwmjfDZ/daT1NcUUAvdXm7M1yG1id1
ZuzGUOT3cXqMj7jS0JPoKvG0mavieYBzEe0yMsM17YlXTSjxiW462/PAtfs/RHRW
WUQThvZqKZjD0BBFnoHQ/eXgR6oGNA3YnnxJWWzopUXjoA41yj+1t+g3WeCGa9c4
blKzAntQkFsMfD4e7qdIV5+esuNL0n8ZRWnQh/EF2yTUfnlPjJzebvWyeDwxMctS
2ZIPQkFmQfKmgpfLz87tNCnNB0+tnvyvuLRS8gT6OVAjUJJS6VZ7WbNDmDse65lY
9kLVd7qJNgxdjNAP82BvFzte8y8wQV10TEdQvJOAasBXj7VfmbnK5Cvc/KMJvsEU
2IGGtcN8aQQUt06AS3EiNPiLsFP8OIJxU6AoPAiimBEYzwMZxmwLTyd50KEEsJ0n
GUG61nsRxGuUxds9qSKBW/ZLvhnBulp9KHi2lutz2Ton/0i3UQziOHk2H0MmgFT4
yjV7AzgaIi02omoSHKZmfdpP9+ufvJfgmWmJwduXDrgd5dwiogiwIJXPyXe7qBk3
/MoTOQCYQDMTqBqVguGZ/BLwJK9jaZgBFGBCGFaVHgxdaEWChrS4HsDifkCdvdQM
pIPLHSjnjLDKEx+cjZt1t2wNxBptpoRX8lnuSbujuF2pm3bfSDZyAwOq2vEgqzao
3SWybZFw1iQj5zn/ndVmD/cOGUd4IWe0MWt1v31jXM1LYkYvEUmKNkZYslBVror0
f/pAPOcQZ3O6REchB6ByTolkEEcbsxPpnrbOz8XeNwZhirO4dv+MRZgK8y6Rm72D
6bvGV44hwoB57iFX94lKQpa7N5ZR+7DelZmaYtwoaYep+PFAlC/k0Seis9DIsG79
KPm4hjAMD6BH62SkDJzOA57H4IeRr78duMDBc9ekfGrW9ovWlFvcCjGjR4AdLoly
97BotZ6BmXVC4c9ZkayVx6Va7AZ003iyhARYO//6Bc133QS+OCYK3674/gqtIPPw
0Hl8LJzntmKDoJjNCUzrarkbD/p/TLSI3XiYxL/Gt4htJaxO5uuILkGzBuTUgzZQ
maTsKoslm6cnJyqI/Kgf9p8FUMzHsv/maNj0uY0DxBbyBxREuQIVngFsbct+XNIQ
CMu+TlXNfNxfpoMBvzjw3CpCaIWV+1VI1KGRbkJf2lYNQhQEz+pNK7D9NMKnVfB4
p1abJ3NsFdXUu+GdQruT5RwWpv9sb3s9pvMILFCbq14kj7r89zLPFvAArcFHnjPs
2OsrSAU+xLhYg/bytArtHY4fSdifwQnZXrch9ay3wfAPlbOrSO6IzxkOvMMt6hE+
AqDauBgufEezASTSl3vOTKNJ+NE5MHfJSc/rBVlbUJPn21YF47gbp3ImX+zK0EUz
SvZHVLO4sK58GyFAowjaNtOTPZ6OeM8H9iLS0rrlfU2z5KxLZI//oEADPeeg3N1q
3TpOFIg/dZMy/tV1P+sizqIgv9wi8YYgf4XMF8oaeiOD9KlfmILjihnycc7GMXvM
99dAfqZ8MGnOHXZC67hfw1wggytNlXbbdU3n6/oRYUKvJvRxErHpuvBZ2MrRE3Ge
WqgLYQTEH59uvHvc/Cqy/lKl8YCETv2od516HbP91MeGdwHl+trMqh9xU/KTHA+G
Y3hmMzBUxfo28TyCmXZJSdahvTAchQnkmAu7+4B3tSMX2DueTxeePOirGQ0ePkOe
j5jvoPqGytNyq4hB7e2AtOvsm0cSp+n/cRMjxuGh06sy908OYvSdZlETV8w85l8s
XIjJG5+jYyvjB1uD5IGCPSsh7xDbHjowN5NkR/LGO+9yrRJ+vXgvRUTEtx9vXo0y
SerJkrCbEHIZXD55c4cChZHy1GO26kIw6BxQXB8f0NGU4+pYvtdASubUMUJHhv5F
QxqhPoqtvt+ioJcoaYiJK52A1XiXyOixZNyN2vOsC5X6E1ZGfLFjDTAxRhBMgzzV
lcl/kvQECaCoguf1ntIO84bXBPsJFBCRgPrQb/anAmJE7L84TNjzEcaLJHnqxrMm
Mmd7idpkh6ggCSlKOBopljT4UlVYA+NzlCYFhy7rt5YNBSy3XtFuSBGM8Wme508q
IqMO1v8yr6HG75M+dQaoFx3OLeOnvNELUTWrqRWfgBZfiIh2zUeO0AfApyiCKTxm
JJK2zDif2IvXTYCHCCwq7rYt8ZKtJ3/6pkvhhEFaJNhegRm7HH0KWganIeeVDg1i
jwnv+OQEPlWqk9TsYR0ojEThw2N0rh2ahCYKrFCZYie0oAr5t2z4g6uyCBJfiA1F
gfO1O+/fAIpUvC631Mb88dJVpbDc+PirgFGhNaAJkjhynbDuZ5D9DZ6OTMrcEZWy
Cqfa7MDrzFSzpkCy7QFFCwBIl1HoyCYMnXYpkrtxReY1AjE0+XYc6GAGUcjitUdE
HKGijVQPLVKXPqAoHSQyr95PcAcnSG7vB8P1tGvutSUzHDX4DfLKmfZiJTexHhzh
TUTyYcT/ZormyJh0e10joBFVwGJr2FrkFdl3IIy5MQ52b1aWJoQkHvu7cASs/o0b
07MNyMm2/qLKfa6ToU6g3x8UcP4nO0WPMe2YKtyf1AH2EiCeFjFuGijWTRQLomkK
4jzaUdNdeNCzWbQuXpcQ6IFk23QAbCzI/UtfJFatJZsM8/ByUzwxwPvqH2xN2RFx
nXxmhabGFqPLmT4llAP9wgHIys2TOqx+K92Fq+k8I3BilUUQXaRMDOza96PkqI4/
d53RDuwUNT5t4D8Ez5WC7Ud0oVqgSMEI7jfvrASSCy0YW4CgwTR2bnFoTs8Pxq91
zNGCl7F68moxUfax9CKfHMwPSBNxT9kNHC4kfT7yJUod3/GPl7sgoz25NAWOxkGq
cLais+K5g//7dqjklXvuRrprKu8JFRGAyQvjDjUElkiUVLDgC8zJ+tjuo259DcnN
gTTkRCCkiitqPY9LzhashkOELWnYAFwC+wqEw4hA77FwjCr4P1I2XvoJoG5S/81p
vIzjDCx0zoKgNy48US1y19e5vAqP92G99LD35uDIW/GC4lwLKVTbdiCM2hG5WVXt
64d32IUr03hg2uJ5YBRczY4jcCPenpm0aBycyiJ1hz84umaYnWa+5xTGOQdFq9y7
TqRGh+GtQ9qPdFQlUQWucH5oB21JTSkaWjq/lrDndFbE8KK5sd95wGrUdlHppMxT
3+eB+yg5XXNQ7OH0noiw1wpTLkM7xSJ49+ZBpV4VvzLtr7NdTHtC4QGooh6QF+kK
Z0iZOcDoBgkWrOJxbfn+kYH0WGiAamr4/ObhHLB4spy5HlWEF68AHJ6NPk77yoPU
q5Zbb5kAf6scjx97qr90I/LRLVnpmkUSr2BjwEw/84UU70+M3kvh5eVaUmtr5GXX
cz3KlF3ERXwIk3pQW7ON/czd38EdXQViSmasVeO/Qq1tHVaQm6607lsADUBvOiEo
/NABpMHuTxQWxqOfpOK73i2+H0v73CIQwRcx2vh/7fiVUhKwavzyFnykdBmpvZ9S
Fgf2IiMXaresmWNDtv3NtAyQ+qQB18/ZEoAqxoJh9MKFaUc9fqGHWNse1kwKtXCN
afKqrFUu6uE3Bv2tvmW6GZj22SX0yBdL5wvKuvcSgNg2JHssuHxIDyupLcEmj9YD
9ZtZ2KpPNA/Jhekl/OvLOv2K2E2KA7xI84p2PG0dz0/v7t0BQWeKJgh1hDcDcmyn
XFFlvbaBcmJwW5sLyI5IlVn203holmdE107dWzS0t69B85QGY6stzIz2/G00b5hb
ASet0mXxb5vGxHAW/wY+YQutvyWUlC9p9EVD0GUps+R71KfGMEk7W7/c+zMiBzwr
CIwgtqBUAtQPQQ+5cfG7kjNTNIBD0xucOQEaZ3hjC862/YxXgdrhgd5RhwSlpmOS
7Y9mkTPkuWGN01h+BA8DwICtOYq2Fgkrw5Xq2SpuNDObUnz55DBs2YBx+qP38Pa/
iZHBZX0/JtHyBvVpIURpLtBw7O+6bXoiGZJc647knhyeDx04y2jeF9a4yegrx8l/
8sryc3JoKbMvnGhFLVsuPuNygFwOgVjzVIA9fx90s2cvjbc5GaW4Cik9HQS5JHB2
McPyum2/tWnWULx0YYyCZvnb27kyOFzLlJlcvD+Pd7tPP2nLueKWOOhLZw/ckWTY
RiECVxq4EkYg5AApa/F9Zyd4Lk9k/sbD+SdngCSzwtEMZzDTQAbkSq5mpQ+H54Dz
075QZ3Lz8sdCXOrIKgiNbDDkCkwdL1kIdu1R5Nc7SymdXAs5bgtle/FUTAS4QzSe
Yjy04vJLoA1sTYlngwCxZkOc60mYTQiouD0Cki309APZc/AJPWwuoOZ3nwxqC5AB
5+1aFOtFiGe9HPNnGGlBif7DgvBWX5F2v0L64qHrW9hzbjEuAQ+kwlVoLuXR467/
kmEY1uDqGKeZtWsYM9O7fhAv34mw+T+O9LTL8koadHYOVduAN9RSrqOyAegZ1ANb
d7ilsuTFaaj68rHYhtBJlQVBmgd+W46gJKwFN6b7EU1/ltkMLamUWcre1s7KQsqz
HtwHgXnID8I5wPvViRS7ldVeH6QDdx0etiKKQFx8/r5yqeZd1jzZnFakpOUfMFDm
f7deAhIzXX2Sg/YL+XcHMPEMU/Kpk28gyiGnQkoJMjQ3Df9VoFTCtBHEFjApZwQO
TzbEHsk2SokLNw9NPSvKuFSCb8rEbSa0KazeRlEwK+zACVa0wD6GN8AYU/gr4fMM
VjfS6/GkCumFp0gSPn2wHXQPJ0ePnOIQR8mcrskdSbiT4WB3sW7tZ9DDsng/bMnd
ZozK5ajVhVMr/GeDDqiX1cY1hNcx7yChI3k3bPVktIzoKdkaHJ7hja+yf3SuiW5p
63EL2R1AdBXmCPZIqFPyQqRJOTkZsPvE6wUstU3m1v2Vq5UbRwc1EdLJ4YhooPwZ
uWOy12HtEq+exsM3iNzr55ePJFGIQVSGqtUYRtg8cYhe5XfmUUxsxFdEDNIfXn7j
pl9y5zcC9mWVUVIWz5+LkxXneEfSZN4gn4qhgKdNjAKzV0sOU+A7VCIdsxv//Xiy
bEDr9v4RZ2ulNKLnimwQSJVSUK1Rb0jGFOUw9UzKPeZVOW1zBTW2MqvdW0nuatXK
JyC0Dvg08jC9vaeo7YOZ9Drc5lH7GlKukjQO4Ktd1MO8D0USpVb6tQdsmTTAztFM
oGsKOdAVcxx/X5hbUfII650iQXH3nd6f5o8ZdhsSTF45vO+3hOzUGxsaVqmtXUPQ
nknGWVS4LEVqVVhZQeWyDb7iVKe5aXnZngDUaly1wgd5hsH6LUJKqnYPGqZLZyYd
hDp4Zgh16ileY7a6saZXUzANuHKdTNCtRXcMe3BI0l8M55zsIEZ53ofwUeQ9dIti
5BsCeVywdXcmoE19urwqk+kpp5HwKOy7uD33VWWkn+6BEH1qcG9K+NBphRSrCDzE
uZu3NKOHMgpIv/7ZApIRf2nDc0icJ9/ymqNjaI/obTt02TaXxADyppLlIzQ9hAjB
6N+JnSN7C4NQ4dNJG0GFmTlg2hE3SdGF7oKf2scsFLVJu9hK/IyGf80yqyJBcVmD
VEZT7Q+FwIHJy42CIZJvAndb7sayljdKofciMX4aBf3VxNHacTTQzr/yD65+B8ye
juiP21y0TYIKU8+/iKNH++W8m0oShva+k04a33e6Nstmf4Ks5wl74e7F7XSiWtPz
DxMASjYpPzw0Ofzn5daMuc5fQ2Vb68lLqbYHTTZnffpm1cthBo6kfybFB5wVHvhY
RkSHO81Th7e2NpC/JILaUvFB5pYVkihgsvHAB3CwKrNlptyBlUxB+dGFfLAAm3vt
OipFVk0pqs9c78zkhKS7HPwv5bq+mKoRPThEsWDcchnZ25R8FbGl+ypie3fMXs5P
ifhGKR+knQ3FvVeLxbLRVJBDtXjCJ3bRMebjR42aXN6dtv1274nOm+/1WOoffzqx
Cep2qSV1S4MkIU463n7gOK5+kf0yVgXkAUxKFqjdOXLo5ngyYTvg+cuMMLkHFu9f
Qgi6gVlvlYK5QYdlOlLfF/n26EA6ibzjjM7Tr9K/VevpjOBj1lrQNL6rx0qMbaKc
tc5AKV9kiFW1jcCIl1+lLNI5uYo2LD3Lqej6JPi/4VKcQRGOFy0cCNcljRM+m3Cn
vTa+VedJWS12Ai6hEMyEywEZwKDcWSlSnV+UmO6ou1cg+PyTA+XkEB79mEXFD+7M
DstQ7WsXT7NA2tCYV0xgijb2lGyZ72XnqXKOEfAzAGcFVSf4AEq+5Gfl4Fr9dqZU
cvnk+mnuCK+ulKE+6DMTgTHAzY8V/3mIvtBqORvgGyW3uhFpnx915JtjaDGUMIAu
HMUzcsf5Qv6WE5T1FZInbIt4SrLt1O6Yi5JDCf66PHyT2Bd39e31+qkwfMRVzbVH
SlCeAxvHQTK5qQE9moCyp3Cwi4/pblKFVjL1P01xShIjisgG6B/bRaOprUXrl2ge
XvVCSRXa27M4WRMPSlzUXwcZVU6FJMFkgzplZudYyTJumGJUt0ENfehnvVNx6ISG
mXdb7q4hdY5rlelZKz2jpi+TK5jG0M5+vaDbIZXB5ybcUAlc/zijyhjMbxz9Bwj/
PFPfFC+IDCmZhi4oNuBbrihG6e1spIdI6AZFJxgspzLVy42362EuYCuA4cr5FdFP
LUoX2MYIHE3wcY0B7Wd/qlH9sgnkkzwe03A6pZ1hdjcUdQWRrAO0GFmeyjLE0zAC
MWU/YT+DlsmvOHkGL2b/H3hX83b2Tf1mVzxbDiwsA6gwlSpcAs0JEa7PuvnrZxwJ
DBSHvFDi0gjezV610vQsl97bpjI3aNIyf2zd7LDa0tzTpG3sjtTLftyGxbN4Rjy/
LK3aYmmbA65JZQgDZA8jDp8fmpRyBtbuEdIMK/FddggWwqopBb5TAmw35+fVEt/y
CZUkDE4oay1ShmtcLYM4KlG2nS3i1J/qOrlMdeXHnaNcVGz/YR0/KPa6lLmuwAMM
bmuhFf9Iz9DtCfuzxAuQ9w3Q/9tb9dRHEv+NNCkIQ8lJQ7cKRJWLtPAANgqXBN7y
xUJYRDP23S4plv38IvXHonvRKUnEeirDZ5TPdJkmEsz23RHQadqlU5cNxbTmERxS
Hh+WwtMu7CYcMJW1o7ICp0LNjq/shfZTue21A0ojOwdIYUJ4Ezn39tGDuIKfhMJd
fBnKqL51Fk0AChwU1VA/vd9C/UyQ+HyZrZNGO6inAhbxTHpmCpE3PFcywOXLgjet
VE6zp6eEUfjlUJhVg4fshHWcXMRaFwfUIZOqCF+ZgJDgRANH+gmOjHxGAHHNXMzv
0smRebH5+GzTafaAfsUrgC5DYsfnzsP+c75EQpJhs0PDe8QLI3iRY7MtNWWlWIhl
A5jBV8Y9WYth38Y3cggFJPav7v4nHdpRBSUSqHvdXfVaw+f0SeAWsCLTwKzlDo5A
Ekyq9hFPQR6uEaFF7L8r9OL9H7DyPM3r+sjZmiSog84V+g0kZInXXRRVoa0/bvE8
VljOFEy3rgBwdUr2bno6+9XQXfW2bzxry7AB0TELfsSe9stUVdk0KB5g1oqm+cnK
AAtPjpdo+ro2oNFmAlmxoEAOXam8UC4TxyuuacO5RX3N2C+H8e9m9bDHUg0ffBY+
rMYQo80EbFRDZ39pI/DzuB5Wj3Xo7cTQtX8YHwQPuICUS3zxshiMnA3VjCQr1sai
Te4GvKZp0CtJlDYpeIKdkKBNGC6l3IbX7BjrKSD4bzAELMx2VUvw7IAhQj8iWysn
nud5k1ynXb2fBr8UQEiC8wmvJQ4S8rM5FbP19JdWTOOFjKhEmFPAt0+J850z8x6o
+j7796zaVMSYsZnHvkGaiCUsQSVcx3hb4Ehc90TcDa08sH5V8DSKKxbVmcegPkgc
Kj8ei35TkkKAFwQSH+jggVX5Yt9kVJ6AIGS33cO7+JcZJsmlXON7IImlgpu1hdPk
1ReOZ3Gfgsbx0zT5aNJ9oiLtjvN55h2oHfixEivzUx9qXvga4Y9idGYrrXVZ7Aa4
kFvXylaiL/dBnpP9mXQP3a+NN/5AjAuppUL9Yd2PmlGdkoVA1vlN70rEo3QBnxZ+
2n9dOtZ13UAzOgUGhS2JUYc4xSUIw5RSxFSs+nGSUIilrpeC80wly3RfmsJMcLS+
UDi2yyhh2gPBZis9KOGac/E7kZZ2ShukzsTILIOpdxAJBIEyFHQelayiMtoAUMzv
UgavmvZLEZiZtSZSVC/B3emu67HRFXyblRNNgYPGto3yqQQQilKOW5VW4+n2pNjb
a0up8z1P+hUVoQNUEknCqz12AKxe1BpcyEIXaTi3ICeTfvI6cslBDqzy1NetQ091
TV8lQm13cMhF4iVDs9PGaEdCyhoAEtP0pin9+0aosCp4ZlLDxEIsEE9jvuCFAVv1
WX5f3VkibbAjUEJWhkJhB2B9oBQ9laaAtCnYhZMgNDvvZbMnb2Hgl++Z3iq1o68b
6IVHIWkol1YHokRtKny//lu+1pxMutaioIgQnBsQMxD4k+MxdQK98aYAiUwC0sbK
mFnv5anYNh26c2oA1lGZUixQf2UHJHEdmQ7rI+B/4D3MMg3gZgJOzwe63ZNiGBMO
49Bmpwc6CChHYitVfSSlcKGTDt3+CcavLZVvRVjmmr101ls8MVuA7j0XLebm8iyt
JVrs6RhVGSUgAQUQ55Z12rx+qlxfWoHDGI6xcFDWU6/A8rOWVGXghD0O4y0RQJxJ
yljTkJYOlGH9k6JdVeqfHXvAOXb5btMAK8UPBrmTNNgPMiXVjbsppRe5eQhCWyRB
rQReKhVhYAAJp03YcEqs1j+hIHE/5fmOV2LtL4wjy/VwnUkbQsF4igSdQjugeXeZ
Qqo4weIInaWCKqifYNtzX/imRVliZD/NigXFoUiGphxgClD5lERUjxAspKrlvu+U
06jY5DKneo2qtfOZYXl++lePAW6xm5vAlR/ec0ldABY+iVDmXq4MNedipELJBn37
gF+TpeS/NJiCtqBaTfNIC0dr4tBYwIBDyYA6hqa3H3Oqvb07meh2G2CqtlSNf8Xq
OayFySLSFGZEQpbEu+2RwmwHrELp1EFvhZ8bIgcQBdc/ankOVlFkyfIdUqHNzOus
eVwgo3CwEcG33+s8JXIOBLjyTUVSS9RWPvPxoou16XOiUKj/betz9SC3ofObsq83
5sRJ7SYoMRnNqPGaN6DWR6I3z+pqaN8h5HgrtW+DZhdmvJKuFdrJTUdRXDhIlEMt
qQd0HqQskp8Af95ihz9udH9wa5q/oUSTbQ9wu+eUkhV9jhgtygiVCtvKPXKTSuye
zOzNdqOqdVAxyBqmSxFQD80kv+bGIHha4mW5gQwxtn67HfuyTYQ/9dhGlkboPoau
Ib5gHU4jhgDnvHwGiA3IITiTtNVi54bbZ4ssb5jGfZbfNSdhyFUoeGIICOme/MEd
s+ijDTS2Oe81DYOBFbTfTZi8VnCRLmUVvzgT8QPfz/XEvYM8xR8Kr35pTGLxpo9X
z9bxe1coomQqk9ypR+Wxtyh3cim8tTY1wbRGHMV2EXFxKZmIFGjAZskBcPW+GPel
qRoeMUHaz51RzpC0BjDNsdUCOZS+Tfz5olGEih301yluEBqISj7DU6vvayjKDxrW
yBIih7WMS8xanPdV7a1wWjCiScGuusxPusJelXSIvzlZ5dnzJjzv9zpHFjgZDk5Q
SV4zLaMN13nN7QPwyJbq1Z32iJdy2wUwjPSWoPc/7i+KOCobRBdQVVnEkHGzedcF
xWgChJ9tl74mUPuafosZ+jT6PEjDssJlflRyrITUSr1HoST1mMO7OGRYFAfrdkwq
7+/22+IF786lCcE0u7XL4gn+wjL1ij/3KQjJoxVVIAALT3oKs6YmUbuVnk1d5tJW
E//r6osdd+76c+HSEFf/oi6ok51odYmE8tFiwQOtRhjnOQUomblvaope+HJEjpNo
Z5A2NFNgd5pm8qcVHLtmUlMulQOB7ehVMxegmoDgg9t9aal0ZkIFmErbfhn8pUjI
jKrmnLSQW1uM12flS3hqt96Q9aXwAiV2AW1WDRMYghD446RQsTHnktYlFAPP25NV
4N34jXmpXQWs938OtTshUWa13Uh+TxrX5RJvxRoFu5UMU+kzVYFldrpKVBcCSdgb
7RqZhKFAfPP8GTtL1qS+Lnyz/1HvkeMOq/Ac86ICozWGDTN2Jc4RVEc3fY1XGjRi
XGQmPsS453K4heAee2g8SleJ1Qys+baDLQcAGxsojX2QLmQilwoW2iC9BBHAD/ce
VujlhK2rknggkD+JyQTNY4+diib74+dWoEdvvON/NY8mr3BIt82XQOwHf0xaRDfl
Rbz/w7VmOByamBiEHOqyB9R/Xg19XT0VIkpFvGQ/ODjvffzE0/FjccUVzNQ49D1n
62YKjSBofyhzArjWQEHmKkMj56cHGj/4E4TiW2ge+lGgLFK5T0/2qsajL5rBMr8Y
0NyUft3DXOpKVm9STGKW753226PAj5i3uKQJduxxrpFH+9FpgAjdQqgXRa0tVhP/
EVUSFr8Q+bIvDRNSRBs9jpYMCQL5uRUKsgkUMnLaBCyssY+ZyWvaO8Am064Jvw6h
2JHiv+tVguCCt8HxdIHsPi9E5jrV4h8OR5RjhMdFpOGgCm/gCH3okRVV6ZPI1RaJ
NAqMrG503YjvwauMgkQ8Wj0tqwctl7hCUO0Sx2HXB/oKt0K5E8/qRxjjD1xh/ONF
8eGqrlo/dbouLRf6E28lJKOK014xexqokRKb9c5hqVwnEniFBjc+fy0hgOcC+Fbx
e0TY3zXxuAnrhc9+ihq7RHAOsFNXQHFYc12JCJ0S6a/yZQYoeFzms6X+Oa8oxZwG
lEXH1jGRQK7c2Uj7xSwUQCphMlfp+O2NHH6sYurJ4q/X964XsQf7iwY9tVacqSCO
+atK76wspN3pEoYItbiwoxYCsaBArl8nVKQq2VrPpRK7Zw8XJY/fWKTsLdFZQFGK
gKYaJc4HosM8v3oXzgD5tw1fIAMZhiRlpKDuODfDjVL1OSF6sDVfRquCnr8eLaKp
M8bBc/6ltwxWvWh+JROX9jlwGTpbHUWHccQC9tyFZP9v06il67zqlnE6pjGWujpi
ldZP+kcfrOsYMjM19hMB4BHy7b+u1YxpwrPe1wa988nc0psS8xj4HjEhdL9LkBe6
bEsJk3M2JBxuEjmU9Q0DmAPAcipT322048D0FeSzZm+DbPPwmXeEpiYh8A0T1t0c
LbUgCVOWbF9Q0qQPGCeU+4T5+ECA1IBYeQ/bjCh4woWFxFQfWRbyRr0UV1xqfStN
EQeUD6NG8IoOx3lFVfBAXma0fII8H5Br2cWBATsfYXIBW9MCuo0kZa9tnnAain+5
SmwGp94fQcQQjnBXr9lSPT2/ybKBBy59SDZ10ZeiUpBEEqSgQaKCVT7iyeH3yErT
GOvQcGleNrgQVEvxA2Mne21SYWtrQkI8KoAf4u2cQMiGuc+buoAiOVufb/2x+uzl
GWahZ+CYVjQ7aZHaTsd6Vh10qfifBTc//28J/N+KcVEG9eI1CWVWNOyFAlOkj+mi
MDGxosvF96NEYnfLfJRXiRrHQOKlZd6eUF5adHVen9peGccMSr/Ob6NmR67H+EdH
XNkQVd/ozlZrvXpw4thyYGACqi+SrqTLv9VyNZ/G33xLVIp401HNCYpE71ZsEVrv
wYBu0XnJKe7FZd+80GJWN0Sgb2zAof0+GNtsyM4vWf3O0kX7Sd43pWB/u1868XWi
qSgxu+K8p5raPbYVBpM2VBOPkkabYP/je5FnpvWHybn8XPp0YULJGnx+r8Xdf409
7EUezlYUotqyVj/wMONMIQs1C2QpxypowQ6rzoUXLmK5SKmcDa77vfaMWJLWy76g
q/IDtD3EAubZeFKftOuwfrad0sPXtr1mg7HGNyK1bkqpEiuvKDgpZWJR7hIFfB27
XJahWkQdup176aF89xQCctI0x5Q0Tnn84WZZgrnQ2wr+zmEScwen7zxP3LJYtA2V
`protect end_protected