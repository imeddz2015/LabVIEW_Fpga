`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 1584 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/9huKRhRMtvnNqb3Z+UU7TahEoHV+T8U3P3ufru7l1O
3DlgtZzb9QxCbOjthp9+wDkjygH0eUfDrEl1ovhZG61f4MdRqxq8c9eydzUn1Pqm
jAGdQzZHVEpK9grDG+55ezqbKqPouKm4/Mhg5s/MwmtLAQZCqdFvx2MN0xe6pPIv
8VNJ70YNkIDPrBFxQczFZUYWX1AScjNY+KY0vPhN9BcTYTub+Pt7ZvYfDzYtD1QF
CcBwJ8UTFXNtdmaawDTyolTAhZnPDW6KqF5IduhjkfARShickplbf9Uvk532mhlC
gFuFBlX6IR6TPk6dWuZNA9yqrijn0BYw1JtJiGlrVDezuzfNC61swe1e2oMJKKlJ
FcSlaQ7QDoXbJKneCjx0hntNQMdC1HZLYbIQ048hTCqm60SoUmgVQt0U8+JIk1VE
VbtGWGBuOEwRCukPhJB5vqE5OIk0vflOWpD3RjIdeGBOXpNchLLvMwrq4Uf0NXGT
2Pb5HLxO8Fzac0SwTfjuKEL+3zDbDWRpYWIQ9+Yttl61M/quM8MhgRMIFlStxQsy
XuURtTrm9KtDUNfB6nX+0qOsWedShMbKPS9+NTEJmRdSQFhja9MhO64hhNi9vcH6
TJ07ekb6MVoD3AcLsSGWqbRKNgGWTBCw/n76jhlT1+gDyCpLwY/KEw29/CpSobaG
EcujrH/gOcZyRQZJvuSNe0PVlPLGAk9EZ48OTENzf8tVI7DtmOChIptYaOUnMTbJ
Gk0omOpQ/9KfuM9eFNVkjQIKJnQ+K8ZJGuzXoldj8V1MXR7J1Zqn313V0dbjemov
+AlFKgELJTggaZifEQTCGNiNXL5aCuzZoWNKXpDoHSmb1hA2iyW0DdN9scngTujF
3divf+th4KGmReKdtaf5Lxz0JCyEH1AjfRrKjZhJSPUXroBohsQ6hXX/u71HrvDs
uje4WBK3spwdHbZhl1/IV/fiKoFBF2oqLiQ9YnZBOv0YTXVDvuwvmnyIE1kbH8ba
XrRWb4tOal5qkiypLCEBzZR+lPIA9lYMTGoGDlqql0rKnbEDUnG35u3vTwI7MOuO
9NqOL8Tg/5II3go8D40qt23hlIHkJ01zD7yvZ7y/Ht+xs9jZUygzJJgfFcXmSyJ9
FztZsAmA6gq54/9YMpLFjl3gFzRTQMI/47WKHe6LaOlBiDooAPJYZE6PLvSce2Px
xa03ObH2EBWKlfOfQN51Km2rxunUNfbkrqxZ2kr7mUhECyF+ajZfxyPbWoOc3GVr
sSHMZe/IlS9RvAFKBMXHSk17H0z97AwkZm2SwqgPJgvATMA+o1Inds4yjf2i0LjY
jO8I5nM8wEThlH2mNsrm/2Du+kOoJzoN+fg/nEt0yrfsnnffOizrv/vLRjoVMSD7
CcNFDgpAHKXCEHN1Er/PpF8UmGh4YfYL1kuxVL7it6gheFd6qzPC34jTDG9e8hKV
BDi/PMaP6/k3lU/rsjyp9t56c0wfRR8aV1b0OyujLra9Q6MTcJaDKDDzMBEFFw4H
SMSCFUpGDMgXS3GUod2/i8UTcC2m5aqUgI7XlvMigIF9SWzXLmL9YjkMELWXl87E
QFuCOZ3rxpm2ZRZC3Lz5WWLO0PxH8OWQs3KDYkSYGnDF7kUb94wCaApGiyeWpS7f
HHJoPWdakEaoCELw2FJnT2QxZq8q/AyGa7CW3H1A++f68zU7YfMLORiYLRXRO4br
MPnZkLmLgFq1F24KxrNmdt3QkPqQ7h68MokldqTVT/xa+zm1H+dM1mQylXtDBrbQ
Kuz3AhfgFqZyb00oeFFm+CNH5xxJRF6RjrBBK/A5pFKfeSWJkNdQCDhoP+Hhw1od
N0xYBglO5ksz0QomPfyIy8R2GFJa9NlhVD97elRZ1/J5XB1Vd6dn1KFFY4Ba5MjC
uyZTKdjZjCm+7zasWme0bN8yiXs4wsGQSogUkuGqebFUQpcmAAMk4qf+G2Ho/mg0
OZIIp9poY9WEBeqkNEfvGT3T7OyE5R4O0uPVNd5kJPmLgH9QU4gsU9kY3h5EuyQY
EScI2q9hrTwxepFJNNeM6Hokbhaxl+OA4DlTIiCgybKBlwL3QZ1dK61NbMUaQ332
`protect end_protected