`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 6240 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/9huKRhRMtvnNqb3Z+UU7TahEoHV+T8U3P3ufru7l1O
3DlgtZzb9QxCbOjthp9+wDkjygH0eUfDrEl1ovhZG61jZx2Zr1k4zgeERGQLOl8T
mkefhqeg+ov3zHJVBN+YWYUKDYnZCF9QVjvD1b0SUCNwnwgY15RZkWqhLqeflRgf
4lPmwseJ7YqtUE5KMYZVJ5/zioFR70XNguKLf+NMxGZh2Ik1A3RKyi7js+8FdDAW
l6LZst/A2LD86R/txE55AzEqVQQL6loqw+lmEjFl/KdXPe76X2s/uq8SPWBmU5tT
Y2jNZOf1FkK79nUjwcvfuX7CEc4XkRU+TBppbB1GtL/+BK/G/ZEwUISPf51W2qZx
ChFSU9Vu0DF+QQV6hkQVSpnc+u/ACOut9CueO7I66XPJlfD9Nr3bwH/o75aFpbds
ldFtvmkImNT+32GXYiOD2Ua0L/0Un4wEPp6aekWW2aUby5Kg1FEjkWAszi3C1OAd
BwwHb+BmRcpM8CmBK5iB7YB9MZkB1kKSpqGLimYCkvpaw75bjDtTz4OBI8pfhPj/
zS/ZrBBcPeLKOnCZRGNzEPaC8Ft61kDkcy5n8PVddD9loRk42q8Twu1wH0CiMiWS
n2NlOeFP1+wppx0n8eFDh4UcJmUeENvmGFAKTc1xjGJexhUZr61rRVIOMug/2A3z
6ksMg14tslJmulfx+tu8c4GfLhYwM62BXCRsWQzyu9KYzT73s3c7ZjbXb/+OAUMx
NW4UvsZdwEDReBfDVkfWPfN5wqh4597eb2rT4/G7G8V87J/svkuOMZx7KgmlwbdZ
XocFg17vcJYxkTZ8X4pa9RRoca3N5FeokVo47UTc5q30aGahFShdn6AT6jW9HVho
AKEwtIjH1w0GdCLn92tbcA+pzJ16SiaqdYIHS2qzI9pBMik+EheDZtvi8oYyZz4k
drnhWUdGjZ2L37vqiVUoVqMwZsptlznZ05rZ8uBkVTsCuE9rwwU5gPTL482bY7wS
IHJy4ziFMS00+IfgPBzv5I1mummyuV+N3lDfn5M+JI6X1+jaAlgM1XR+SE8Pj6EX
XlmMfNOExL/SuIQaocfS4dvsO+yyOMgSAstdVQPyFVWVm7CSrOaB3816dUHAN8xo
9x9VWNwAHz6znTLJ90Yu70VqgykmhTIWoLNCYRUpvjwZZX41QAtVGY8SbIct8wvD
XqmzSTCBvVvFDmLExj4OSlSu4bl9aHElNjlrBCmMjOt+wwXXkXs3IvtRmMefmte7
FLGZ6ifd0OkDaYOT0iGW4fNtzguvyJw5yidwcPMyFrrQD4FMYx/R5c940RtkNRFU
GiHBAS8BKXKTG5msHXX1sk5qfJT3nrYbQ4XjwoejYELtg9HQMThOWSGVG8qz5xdp
H50Qa5cxjMVpGWXlKlSKgjlLxv8+ie6VSIqts4kgU9r1VZc07esRAqsUjux41Q5C
/sstajMHXCBWpcFyZr6lIoQtSoXn6h4GcCgMZrwwu+VHAxuSK+YszThqE7B5zt5O
0T+DpueypRkobO5UNpiYpcuISqSK8IJPjLrR7b+/cT8txC5zaxwZAE/befbreI7+
c8rph2WuotiZJNrO+RTG+yNoGvUlDXhBSCOcDObmtywXn/jL4BKOPIZ5a+pI87Pa
BcxFG1RPk2E8na5Nz16HZuTXp/gM14qYElP9lNDrsJHdYgXMTCswdu9/9Gg/rSE4
tybj9NAqK0dvhSORRr2sgFqAbHCtdOgFpRUXPCBxLFIS/1w4U6mR8ek9LNVl9biu
8qssHuJUyzqwU4BELO1arN9kp6GD/GLAluMVa//ZB9Hlehj7gOqeCTltWoCKkDM8
j9CycZKnGnYGD/KS5QfJoZbqBAIm6zGqLqADbMZzDpwIB4UxzJQKhwAIBuKgQovm
W1ClgdYxwK52kTvf3cXDjufViFTzIWKrnl1GncTX38AwID2zGJrIGl1nuT+Ldttt
MuZQWGLVSnCJIwOrvqxiJ8pfMccb0qd/r7PPeeMlG5mWoqcsNOh1fmTkRbqrs0RF
REeWYHkAW4ZLMSEYkUpz7QV2yKCSFxh2dq89kcCZoWVsLSeAn5I/iNm8Ol56P0/T
457gU75jOx3XziwWMCT22wa1JqzuXhJCLFdGhSk2IHXX75V9tI1TM+hsfQIuNh74
UwynPg3B4e6tJ65Xae60vngKAuJIb8Hg5qbhbn9zmET/5DbXplruEsqyvoAR04oa
piKFhrkRjnAkWB8rlfwDTp7Zn9MDmGcGheaJE+QLR758X4czmt9e7nDuf89XNRbs
rQYBAcxlmnewAFwFg1goyuLzgPCUqwU31e+VSTK5aeG4qvU84o34jjEompj+VUhz
m88mppoL+f6t9OtbE4b5dcwGLYnxdrfmV/8/PY5WWqbZdQDazOMUq8WnM9CsP8N4
acxtfu0qx/5c3X9S8xuaZDKzqOb8NpWGdI5SjYJgn1LU/jNjRy09Zmp1vwOOgt0v
J5apquWjic512PmagrW9w9Q7UFkqIR8iyC9Kx8YimDBzf5Hm/MrVKkFr9iNPY0/z
Bej9uKGH8vOtQ0wSvdiT28wxsDw9JV/FsENZ8ZEWnk79WE8LU5P2KtzGg86Hp4bF
SOX7XEWmDft2T978lhblMGPKBEY55EPcS1FTNf++DKQrhTiPrRwqorzZLvG8fsuG
Y5g3DCPBJtJSy4Sk5mIfqZWfUfyD6NML2OvtT929BoXR+b99dH3ugEpaInGgaF6K
NFpQs+gXB/xrFToexDQBsXRF2OLStDTRCbQi1q9MEugYUeE4R4vGdNNbI18LR3UY
+J2MS4ZGsVlaE/cuC4X8r9OZbQmLMaTSjGo/RD2PnLYYUmyB57p0BPQK9EwU/eD0
VwOJhXFMPSR7ufJt/Gf2hEK4J0rHwCM2GCehxRx4KWFJ1NjJYk5VU0jbIcXT4U+g
P8zeknoQ2ByDG01mDTUK9I1B30bT3aRiChWsdb5NhZQblxS/0nRNFXVgQwoOQNBY
Ox3EGSaq1kv9DcJMbsjqIw/uuP1VRssXbwkbGno7kWKkJquqjvqXERtW+hGPu+Xt
sUy+FnrekoS6mKjWncSpRpfWjsTM0lAIlyngYPUClNzHe3spB3afxMrsrDObjM5C
UvyrqOK/ubjxkjpZXskHsMHXwuXtMe1cqjccX03VLoyR88BoTSqLALSgxDQ6Te0V
k/DaFrsuWR0MnsKL72km0W14NFutsAF/v1+C/rNH/vp8TS3zqyLZrCDj6sYf4myf
UMc4hxehb5P2UQQLaeNDrQScQgAyzMEOT4y16/CbQUoZyiWvc3e0RFEHnxhnFNle
lslDK1XmUPC3d51hzU6/PDCx9UGmfpNVL8ld3Wum88OFuoORRWlWLLpktKhF/nJN
tJExDLuIShVPozj0In9z1WkPMFwn/nJWCJTxJDtmRpeJm/ITjaa4U1F0nWC6dbrk
i6rWQQpdILIYcWnSTiXhI11LMeXsAOJROFg1xQRUoIwxl8WjpXRXqXJ4MrN+18qp
TzgE77+QLLPAN6UtxcILv4J7F3gciewe7lZFo3pYFTqLgg2DsrSa07tMwQpwxG+f
Ap4p/fUlNxTrET6ysWyXZuqle5y9N/Old8CaPc+XezmgAgv5BsP94ZLZyOQQSnh9
UjuVnW09533j5fzUCvtVKDNcHQAHp9qJy5Mw400bNTnvzff0dzq52iO82X/ojRbS
PsMq2T92GcJHuZI/k7OoxscSNW244W+bzgTOukAnGb9TFNeYJwswemKyRPE8LmNu
B7qlVwBtTESDoTCvdouW1g4x8s8zrAmNM5swSLkQlhZPe6VqlPxAufVfm3hQiWWA
7wOA6DKOG83IzN1CczSg06OxSlLkuyz9bCXdZhfyENApbnJWQhXrRYtEWLMo1CQB
RQMZCwM8Ph93D3rDbfNJk9tgrLUDCexzJvoinssJv5SlZ8tS8jWeBS5PEvI7S+Of
KIwGXpMpu/omjTV9uhkvDXyR/jhQBRV4KRxNK0Xy6zbBOZIZI3rd5N12j+L8uesz
EL94rtsnD21hdyI+KWZ7vyIo5lzvUospKyFQfWcLd3AKcPa10s3aB1ufbdWuVWq2
QLtar0G5N1VCJRNx9XS4hWyj3W2WZGGWzEzlLHytGO9aL7BYoDX48Oei7u81T6iF
8XA0dgvnp9IYIp/LJLEAUDb/5tLndYnO//kkagIPPLbG3X9qSSWbhC5NFSNh1myS
n74ikJUofk+A7xTQlV8feQz6LbGe5YCHj9v3NsvQn9C0tFIYDtdxOqVCRKDu92RL
P6vdK+jPJ0ameTQzHTymQlkjG13oOCYyCR1FdcZVdaW11G0U0xDnEFIXLbGBnvL4
43r76DTlhwNspCOzMB7wgHPyYiilbzH71KF5nFhw45iL7K98GyfKtWQWT9yCHQU+
RHukM6btnOG64lOguhhHYXwuFqJIiL8dhsXbWrvpctiwEN/+7QK9/+Duugw85Uej
OOoONbf6WPup1PIHSdnh5QZlAcJO03didAzjnk/hlh683OvAFJl9RmVP2nXrm+4+
s6v0kcN8PCYNYRDHcEqxQ/zz/BI0EuyDZLcN5EsbAHhhUo+kbDdsFEgqI416WJ+k
B0u0nGn6Krz8kDJ8tT+XDHsYa5u6BNEx6oW6y6Mz41IhNHemaZfqiYUmVUALJBs/
BKlNwrjSr1JoxmJRi6eahNqxE6lZnTBtwo9dfR1PoP1uaMSVFiOsaLFYvO1QhmJF
+UENO8mf0WAtljnKS1p/1nG9BVQpmauO7ruyJgsMiZXiVpSG4CWPDocmQM0oKFtX
Jfd1XCvNTwQTaC4j04dH4q3x7x4lfcCzF6MDyFVTswSDSvUfXDgJXJQXtabWJSx9
limR1G4CU9YmxJhATgEanZOlhVhhXj6wveJAII3xtS0b0261NeyvJImY4VkTRHCi
qD1TiC4d44SD3EPOxC1L37perA4wkaPl9JfcMYwMKTEXTOH/BGrVMc0DgaCn6zEl
vgvHAr72RLbHFouWvvqPjbSbllgmoOdHqvlSR24sd3+SitK37Wt71oWVEbJBvFjh
Pe177Jwh3TB4feemP8x3Hh3iOhFfl7p9kbPu0rA0rnXwxssUCT52PkhiO113NUBc
9zuwPSiiqeXgLX7YIXXtcYPYKr8FU4K1Qgj2eEmIXvjAY4shWbDHAeUIQLH/KXcW
K3sv4bXX058rswq23vF/BmnDRvEZ0GtRZJFsE3KaLQI0aAwGjRMEZ6mH2MJAsra9
LkE5XOjzdxJDIwiLqdCd6YKpC63mM8aNMWnASvSd8x1C1vj5HiAiyL1bXiPoUbgj
/WiLUtSBuKBFXJgFXBdWCVvhXvWsu0Uy1XYzEOUe3RZ786aTzlqGcstbmFxa2iae
IH9stRtte1F4r70F4o0g13fbGuVK7mngx68TwaBflCj7Zulxpa7TkRydAEkRHhR+
n7Df+oyXekE9YWvvE9l67FzCefI4thBqUbBJtVZlBzu2Du9x9okd/ahpcu7jMZ/S
d/o+qRKVDZiVL1936pPhO4L4pySl+Ls0DGJ/ued5iK1JM/2oOPp0op+BPCAhBb4m
vMnt/Ukj+sbrkCu8W/L1k2UpFUf3cmgI8uUWbBvjVYcp5QQLPn6PsicPKTBoSTrH
ViAxiy4FBrWzQoMMxZm57Gdncbc/VbG5xr/vu3vYUjErj1YV4oiOdJquuLxQU/lr
f1IpmrMz86SOM+al+IMd9CoxvapOiHWCDZpkyzsp2lAmeiftX+mLepxdN8AakmsH
jkCyO9VhEBu9VAnwyDqSTHciOyFbJw6Wz9PGbS9twds0UDcVHy2NxXuwkgu74TNH
4f/BMy2vY6zgmj6d4GLg15XBeadBDYKgG8+2J+0LX9YqvvSFTSU/HnlgW4TaISzI
mYip1Ov/BZEAKfLF887OB9eFFR98XbtTqZneaOgsKqLqzwkLyqJ95/u4M8VTxjQE
G79eMM8rQoLcNMt9X8UL3T9HXzvhuomVEm66AkU0lNOTaZkeUHFmzZ40WwOry5d7
R7Pjs3Jho/ElqSGdGSdY+Qc3v5YoUt9NYEN7fS0H5a6fn8Fu8JkDQFfJO70txFIv
jpsYYtl9TNukj5LzD73QTbsQlngVFALtiURSP+p6DpQ8+3fec1aEicI7qPaUDo4m
UIykhtKgzYX76MZQ66HgdCGBcKQD4zetCRARKioN1bam7RfdeoGR1dr6+lqDacuD
pv+j5l08CKY7mb33JnoWb8Mq9q+NQj/eV+XNOkOvCBVrdUIx5V6OE3pZ6SXmZWaN
DV7qgdRJwhZ+sRjQG6rH++8xd1npsg38DgcuhOqpPldvNd9KKXBGK9Xnuw4rLyw5
2vSUdNQmUj/4R10KaucVkHODmdmekna/5e6xxcW4uZ4mp+mMyWxVv6Vd/2l1YOgJ
gp+mgQwMn3+2kCE+9WjCC75Oo0IMXpaYlVAaud0cDpt077MEoeOUweic5QoU+Q6y
CG/MgbLD/Ecls2dfC/RU0WjkSD3vnchpoITflkWDn3nepsnh2nRqGppVaHI1IGl3
H6SvmasJKxvBFx35Dg1teDBoYnG55sQmTGYvGYwhtcM3f9YvNv+X0rznQwmUFUb1
MDvsJ0gC0r7+0P55hgjIoMdDTuP6wHNneLo5S+3G616QyL2mW7xjKwtEgelFt44j
4lPUGkkKqyFNRVVGpCX5qdWlO1Rbs0wvxqjG/d3Ilz/ar19GUI1s/f4+HFUAOonp
8ezAAac71toaUFoHmoACAfPS7RVxgbMiCxtl106G+oMEHYaQwh9UoGJ6UEKi22na
RLw2VEMXsbgv71c7IyNqRWbfuCuDoXJ0GfnOX1muQmpJyhALzmxl2zma086N0eCc
Dnlq9MIJ2tKy5YP21Hqz7U1NJ67pMeKAEXgRJ3BXIu0Xvf84vwgM4eQPYTYcpyXs
+QckWssfLPsvkIbi1tjOTBEA26yyMPrvRHYRXPdvMGFRvHMXQC3W2zXAAJhTgode
nFccDGK1mOYdYB+W3wakQpYSauBPynHl6wLF6l8oKjMfFUh3xInyttEIkHWPzEKJ
ZYaTW46sUfQM1BVj3UAv5YKAgu8YNpoM/Od4zD6q8hUjjsUT2AvS5TG2+ie6axXq
cG+T5d9GS8diMMm9pIWxKhkxljtivo8ZwHzyI9C0LPVVATf0Ng0TP42/6+t9PqHU
2HuIgZpTgAGx+Bn6EW+QexJ/0E2zy6agwGJrFKOMSdWUkUqoyjqhfXIKnBc5HXYq
RubkJuMI1Vf5YpTDuJmLG7NIhUuA5OG2BY4e+xrV+lTPrCvZ+6WrYCak208ymWAp
SaBbQUosiVcV+ZSMeibu0DZMv4GyFfHvJiW225tqS3j8v4MVLL5ThjlIZVMvfXoH
KpdAYar2J5x2CFVxdwWsT7L3BgisVuw2CpQzQky3bZ/+OOe4DqNIsjddvQkjKKf5
FJHPyNkWQ4Flj6/rSSjRFIMAyxGbNumgfloi9p4wFa0pnWJGypv3lKlb/+OfZ9K0
Uk9nR1FjdqCbLErRsUYsx1+ZHD8fRdJW1XOzY2CedVASQqfHObbPaGww5KO6x8NX
QZSsagOvRl7MmHlMI2PLPSbSPVrZ7vhEn4y6e4X2jgd6luIZXqOSgdfTzUazBECM
Nn9ZgRC7ctpEleat0A4UaghM7MVkdckr89Yo5oGEtKYXK3crBK9c0TTfMZT4dX4t
n5T0NZxB986cjpZuQp4xQCNMJmn2W53frcK7VM4upj3hyiHBEk8VT8gMXXFOuW1p
c7voVmx9cXRHokgDeuzz89AMwMzLmw76TQrS9hKKSq18/+YlxnLd67sc/Gqj3TRa
BrpgFwYgzH5RkFs75IrLTEQ2W+kGUtE0FpkGHQ2+xKbJyI3/oBObFJD3scUQH0Wt
Y7bVS6NKS72N1YoPwpyvpYRCk92jEQyL1HAanv2OaMMsuPin1Hu3CEmE+KrdIJU8
s8YG3g43LS83mqW5IlaI02g3+NqtVoyGhleSZ2wKoW0vg/rKmneydqtvcIo3ubUU
CFsLLbhJVFYPJYXy2NzxwEDZBM3ln22yX2NGXwT331BDTsObiEx/tXQuZYIqU8JQ
9fDqUJj7zowCOV+2EBU4joxg+QdTQ0IZ8ms1we8KzaxsM0sCy+wOVb9BRLzSomWj
ECzXJHa+P6MRIKRnCoU2Uf1a+1U378W7BMD2xKm+cSf6xn2OEoTMHBTcXNWLmYjM
9x0nemjUiAiLsRJnpUMHMZae0tPSiVCizM7caTAqx2bGIWgvG73JhEj/0yhZPVAu
J+PDC27a5NZ7LkSRMAQO0qLqn+FQXMMpNWRMOebVsMoYrmqMsCL2BMyIpuJjhEXs
`protect end_protected