`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 1904 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/9huKRhRMtvnNqb3Z+UU7TahEoHV+T8U3P3ufru7l1O
3DlgtZzb9QxCbOjthp9+wDkjygH0eUfDrEl1ovhZG62XW3ylm2JcFKIzD+72jwLP
JPuOOUgCYNfPZ1CtLBG9dg0q522nROPuWo4lj5Jprq4hUChShqwP92CTKHHC6LCV
W29WcvzhbVVH/AIXilIdd+eRfP7jRIGbZIPloojqFQg6HNTfUK+MoUQZrskro8Qh
MLpFPFrrHq7hRaYQz1Yom95/wCEFEUpZBYoEfLZ7ElblkrByzijKM81Pmw581dW3
mOUtBbBe3hvCvLb2ehS4+JaCEkkgLsahCbcT9B2TH4HmWhW94zkRZpyV5oUCNVpS
550tkTQim0HFc9MN0VVgrt+p4MGZAHTEUXL9fn8J4Pa7D1xWyxujdS0FXiBCXt8J
xK3hLgiofGvM1D2YOlEy+r0SV1fE7+QmGu2HzOKC2WbxTSfIUWED3ch3GqdfjO7l
E5CyoU+FffxbgpMMm8ag1vitPuGucspjaUS3uQJZHs5D2vT68rbJF3ea7fR/wfWB
yu9dXBasCfiyZWApMpiE4IsM+LwYXmO0wDRY2zXty6Yid19vqae5L7eYR7JC/74H
ZpFGnEkpUW6zJdemYhdl81j5jM3bUg6zTdXXHKQDb8TnVzw/g+azp2MvsC8vMmLw
F0YEeEaXeDrQp215jDk8PYco9GfA+JGljfqqBBLLuUW22MljBLQN42/IiUf14dwP
4MUBOPfHNB9Ple2v32WJD/YN7nyvCzhP06rMBSCi4eca246PzjGNLivRd6YdLPxu
fh0G7U7RMIOrjoiM/lJ4EZUs0LkMipHZWqTmj9iIaUelwSfow6iSJ1m2ziXWVqfT
mJDXRkH7OHq/J5wA3IDRMwXfo33iqM6Idyc9TLNf012iMEmttR592rbvXpYJMCC7
e7Bf0azNRxqg9qj5PlvZsym6ET5mK4ZEvvOMIPgvyTA6lIHlcaMwVuyZ4B2a9TOK
E7JsDAnJymNzFH+8ff5YMcYOlefBSG+NupoLjeRISFcSWEUPDBu81D0q0iZ1y08B
8OKY2XeEmc+1Ay4Osd9m58sVfeC76Y8fd/86TaciwD2RMyzIcQgw1bCrJ2v3MPDp
qMMblaFk1u3EFHYWVX3e/AeJXmHVpxxevCSCTfK4CwqWxw1RWDX2wX8fAUKX9ul/
eiRfvM3rm8f1kJKkTwhKmyPzfEeFm7zxJPIJvH0e09FBcYnIlhGZi+rBuznYJ85F
uVf0DEr/ZOinXZUBmc6VmdrNiLR1xK566HmTcpnMPD9mTSmlKe0VURXSmLND5n/Q
v8Wj3tJYGdqZeXP5kYvjNcYqV0hDpAaLP/vOiwKnl6l7PBXeie8BcF2bHSn0OpHD
+qlh2aOVF0iH97PYNRb9ah4wc/ufUv1Ocow+sMh+MqxDcuxqFBesHKb+PC68tCFS
bRD+xUgTvzIyVww/KtpD7Ci4/khVudfVF4OLWbLP7NJjwJMYya4br2D/S/aT/SfY
/3B6vTPpJ/33kSsefNa+NMvaC/fNtj0KMBnaGNRC9UJ43Ds4kvR8P5Yyna2qUMFK
DAY6UWi1sZC47guPPkfs5vxzx5WQSRGMZFd2GMxITZk79J4GX13POGmmurEB3KnY
h7fwr6wpY+2NtkgEj4RmZoQ30wEkvOXTtvpch2optW0CeYg4vIp5gXsYiPVUZEZL
LMV8OuIdjysoDbhQ6m4FnBFT/oa3iQRWiJnTXv3myFERTQnJTuJbw333aWVtnxel
E3qvSawAUjHe7BZi+f9U2BUysNVyXSwK+TlnuJ7BhzsxPIIgMoFghaUT5zjP1T8s
lRalDo5ivMJu9Rvo0mb5tz7lVObpqrE337TBJmXYVblsZEXPdacsYgrF7stOUdxL
SsITMeY5wSy6IcyrrCGSuBetddIPiVJnrHWglnVm19Oz+0n7O3WJ/NvsqsOYlQ5n
87BWJcCmEA3oXdu6zdrlwVbb0UEd82QP2qBS4Dwrzq8h56zVpENPSK7qBKpy4Rra
myqN3mhkJ8XS20L/ri/Qb0iqmazui3PJmQ/Z+TBhy/DZtlmfx27KFmslTOvZmVyX
9Rx+NJkt4wbpszciVJQ/XO3oeCgWEF/bmmdPeHf22T/lKtgCxIveD5gnNYvFnqou
VYDaV9PYQiHG0AV4i9K71sKyGiBaVTuFwZqs5AZF788zxPbCdmlkH9+vJ42Y5UUN
23JQBPFvCrHRngTKOo/XMRpf95KNRYY7V4j3ZM4CiSxuVSqzQjfsGWwcf1WbjbDq
b0Ypw0Qon1UzcHRF7c0asek3Vvs43o/6mtNp9oEZnqkm/gOuNxCxi0BXDlHajamS
ITE7GtlODbw10pLRQIf7/7bQ8a7qNcHpdW+3/74bMHscrq/4xTB5agwZ2sDFsCfm
zCPP82XB+zBGQIGGJFFAxYsfL1BJfuDnxswmYP8BRcrEQn66Dbsz9vNk905g7u0e
NHT6cbwoH+kTopt0ayvxk0tCxjyOX38rtxoeUUJTaQk=
`protect end_protected