`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 5424 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/9huKRhRMtvnNqb3Z+UU7TahEoHV+T8U3P3ufru7l1O
3DlgtZzb9QxCbOjthp9+wDkjygH0eUfDrEl1ovhZG63n8osOUkmmfEmUlQmtIZxm
8eyJ4ZEH8xAds1oWLJgQjs/5TKT72hd83WAS0OhsUSZQmQGwvIKyUfsNEuhiGx9D
UnZJCsEzNK6ja3IidTHF2CG+CJ+z+qOPwt9WxOApDnTEG0ZS44dFyvsdwSi/Zt9X
lfdTG76mcDANyo2y135PoEU0HOVCVyIi9GCZbj8cW5/8Jbg83VZQoRX6htVQwLFP
rLR9CwnTm6tuoCM9+OYobj9gtYE0h1jK9K69UizwPhIo9piNR5ehC83qKn3xVZ0z
HmYOfSh+xTdJmaYC1SJWIRmnpHzjKmGjoFxcjR5Geot8Nxkbp3QEvQd76g1KSW1/
GAEHVbcyqNTcpVs3478lfks4P0BhqgWE+aXsN+LcZxxIpBVNHzeEtSBNGOR1RfRS
wyNCGCy4875vW4IpA4pOWnZgo0qGh/ejOA32HbdGcGthWGgdeMymjlb5qf79SHS9
TCWjIv67piP1wr1eMym2N+Lr8p1LZ3jDHKG0AMe9QH35dwbjSDkHPfTIx5STv3Bm
Pcwn+LOnqM5i1Kj7YKyr4lYQVu8wy1hZaiA1kHCmL/DBM2x6q7nBJ8jGXJW6ba/j
gtDLIa8/36a7z6OtR81WSBGOSzwrlA6425Ct1b/RBGSf/C0+l5h0jgu6cLW+Y4gw
OxWSMiRJJZLxFAlDYnWo5wPvehI65EyTJByl8Z4jR9P9R51+MSYMupHB62FchkJQ
mnPmosKDy3napx+c694GidVm/YkyEcfp0+HrzOhulmy9Jdac2EKmkvsTFHn5LHBc
xrcWEF0RK8nGiRg2J5uwaba9cddNf6Jnz496ROfU5Dld8WeXLMMzKp9zsLyOznrW
FoSetgNjkqG6WeYqlpajfs5HjtaSK1cvgssxjZx3XEPpyPy0wH4zTZr2zrG61Qu0
nacSlh3zFNhir9ntY9CC8VAHhyhvYU1cDQ1SoCCEwyBO5aOhoGRgtcqSIUYQrTIu
Hq9UDo7atDh+D4OUFDrWkXig+PyEh3iOmlxtBWKzLfwgmWvYrbQY+afNcF63TiFk
+xliyC4vUOe4ff6bs2rTX4PVmhEBRFYgwkYUJwuwCY4gUHWJkYdLiPdvWWJQZHvr
LzVC09xTzuYEvfESsJpHIjSDlrJZXKlY551cYu39RPX6io9Hf5pQqwJOGyrBpR52
kbxWo1W2z70Wmir4GpmxEuu2CnFNHPjK+B4mNsVNLLF1Ct2+iu49kJUpZ9gMyEfA
v5VHXQpEnmRQHXOQUHEmTVPiIL8gcYpu6VSzEfCOM8UfZETi8eE01A9pJ0HHulSf
/wpFZH64U4GCw7PNbUDhfAabcxhddyTVy2M4JTrGyn6lN360RquCAgFClXChRZDE
ZMKMLjsdmnlFQavbap7DjYwArrufRKyxQGXMo3QaFFQK0qc+2ttpW1OB08Uj59di
W2dBsjDVh2fAmTl4chHtr2JBpCtQ8yyTE/6aG+r3u4vkzxrzkoAuDZ0HrGHHG4Xb
8bjTsjGMtJUMayA/3V3g2sP9XCRawlukQdHDl8fqjvXj9nc1QnNwfSRCn+KrFDkP
x9l/LC+GjbgWr5+6ZD7r5g7u6B22NxtpxCXy1r6b4zPrpp2owiWtYsG074dgzvvs
4OvyuM+Oa7b37K4mQa57S/43Yrd8v3a4ptQeLZVmsiCEHnAqA4eOb0Jsfrldml7a
MrlQya9QSsgIX2FySsUdmkV5C5o2v2y0fm6V4pBYfgCxgI2e/nXyrK4mVIhmrmph
Fl8+2VkaQCzT8weI1UxhZVPanBCdq71voDuEhbzjmgBLDGTdE9TAZW3Xw8jRCDs+
BrGx2bVXTS+qt/4t+S0w1dmfGjC5KRbyJpDbNdmpNFtsIDbyMhU0WZ86gjoAkbJH
PbZfeYpqoXc9EceFr5f5VMNRmIPinomhZoFVaAVqjzvP04xIOHRuBEqngRZOuUS9
4qyHefGgX+HizHB6mj7DirDJeNyjMmf2dueChpWLG6DI3XzgkVwuMeEYBp2kBAmS
s15oEv7zGzQVAegGqD/2aMCqdDQ1U4kpWZzYUwq3PpwkqLcnxYXatsM+WhT6Yh6+
FQOroYc/VWLVXXzag82VQM7lehmrCqM/8fzEZaYOxCImdScqYVjaV3WkQtMpgDWm
yVEQdwZmsF4toXnWTAP1YRt6Svdce5Ippxq/qNEGazU0rEMTzPnDMCQ4yWhvjV2m
E83JK3ObNEuGYdyble6G5z9Xzxr/S6qzGXNqiQTbluKU6uL9ILV2Ttg/dkbmmkpL
ba2WOO77E25MQfW5o+FiRCbYsTK3rdxoGTRYlIxGzCVvxzjwCILyqQa3C2xXwk1N
DqwEoLEEmB7XJt3YA9WYbYPVdPjr4hK+4Isyco/Qh6vuJS8CVt47y3pyS10xzby0
x/a/UzYDZnRDEXvZ7cYYXQe1cjXo/I9awKnZKBeTUlNmH4/68SZbDOvANoFwFLyk
WJVtjfmmdPWdy0U1bNmsjC6pNfw4C2x+ZtQMcwqGanA1qJu+jy3x0cTg6smBGF/V
WseGBZtOz5GY1Z1Io4WW9j96+o5OAntei8inKrsWpb2QXlBWE44Zndngy1w5ULo+
LUZyT+tVQGe/ZtqaT6PY7iuFtzg7UJJRVcnSUOEB8GqOAalbvw/BW2S8kzG/IPSs
veI103n442HChwobU7BCCOvC4FzMxlKiDOoUeSbh8oDR7t4rk6SSH1Kf5SAGGw/a
14X0i5YMb8KPw87ksPrV38RnRGWMuAm8sBCo9HhZEmEmztWEPdR5ncT+JZuwEic4
fXGADz0WV49B2KhZgyfmsPLWfv6U28hH5o2vQHKIvLICgcHaPnPIEjLAc0hE343I
6TibGhqx7K9CD68Z7s8x0eX2/X1kOht+Yyd9CEKOgapM57TIDhqZyrna/g73stDE
mUCtZOIPV2/PbOI+u+KU4zfv062Ln7hfNBUJ4+IQzKKC87igRNDiMW29QpWeAyAj
l2/VSNBD2qOLRnm4FXL/zOGYrC/z+ETwIB1JVNWDqPeqDjHHPl3zpdTE+QQh1WDC
fIEZiymBBnSoegDMf+bZRBM4UUreVfAhNkskx+29CcUy7E8JVfvEvZrFcQKNjGR7
mJr3rCOypBDv0PU/7fU783u9IPd5OzXBkX1YkeRZZhttLg1uFDaBOlbm+ZvhO4/d
0h/o3BGV/88QW41lJjl0VeN0T7vlMcoDnFgoRXEX9V9eLgdzM6VlpHUtjGb3dXhy
eejHXN+EdmBB7IVt2dsHgaEtQVPFVRpfJBRwdduMFW2iC7ImAuayny1oeMyZDcvF
IdbE3ljshNMCioyNVqShsti3F7AJckfoAhcun8SgQZN95ktLkCzE+fC5yDJ/9y54
jlD+cofCo0RaRTZgKjmdCFp+lJmtRGAldjJMIC1Z7Byvi9SAo+msNFbdIgZlqDpK
pUSRFtWbPhw4qYnqqgj6c32zqEvD+YXTHFNxCYxQzEGoZjLxd/W8sG3F1t+0meD5
jAwr1xBq7O+L7u2igGWsqIERtoGk+sZOmUu4Xkude3I9CrPE56J97IWRtupYfl+j
PEHBJ6/IR11VWR6doNhEZaZX1jD3d59VoE4ajknRlfOHGodPS1mhczNh5pFCRzU7
hXTyJ0T5Xyk2aqBYAvoqKujqQqC0CsTJ8yoXpIY2jKjrgZ2KTCh9uFxHRbnidNxR
dbsyuFW0920lWLd3TjIyHgWtrQ9MzJLlqBheJsKpScCFVVwCa243Ctv2ZY7ZdVev
Q/F74iIlfFfM1SiXjvLA2IBDyJdZR18WJxVMZ8sg7Sc0TanxQ9zswm6XmYkhYaBa
9Mxc+SQ4r1s4LQclmRycGteHBf7atUgyGuyFUBdiSVSrKf+1ngnaiuWdtYlsanK7
TzYuwY9p0ijNZOF1RBgCQ3PjvOMQZbVvN8H894qZHxUKjur/tB2g+PxwR7XyNGu9
P2/t1KYiekUofqUmKtYLISoYwzguJomkfH3v3rcg1fJmB4yVyOhqce/qgGs5pjMG
cB/on7KJ4pm6ETmsIDaRxBdRVel1ZjZbWAzKRa2vHkowPWIz2uyD/RQ1QsLgYP2a
iyFJQs8Y+IxxOGGSSYLz+ZP9WcqeURlvvIRBHbi8KBq2WijVOOmEhTCBaB1RkT37
/YqSAfBknQD3uO8BkKOm7ZeWfX5Mf1h5/wLnHfsa81pw/QQQca+CyL2i/Oh8YJy8
WhyJqdQAEPQEoqGYBkhWzRM5wqGEU8jaxyRJFfXkNg9vWStEYd3g+mqoK8TGe0IA
W2ObeijqV7CFbk9u68GIPyWmSfMm1rQCK5xDtmggI5/Y1dDX69VhZOmGbl6x3jZz
SpVDkGbZBwV7xAdvy4CZYz6oMM6N59DKNS/95A1uFZiBpTq2vO/vGkXO8XOKhaxR
KHe/7dwOKnKts6ssxPaf6NXtRGhEEh1tdaslezTCKw5yLqhANMX74YYdyxSlc7IM
E5UBoQSRf1+famNoWgkPAZRYXnnDqzqcw9ZMtiooQFXdjDEiNg1YLeMqMghIWdU1
x2oYIwUyEVM2vC5r03tMLJl1QoOcCpIie7yfZloKmQ1WifNlJrD4Swql5NdGODJa
vVPJEGXDsI4jBW4D6O0GkIzFWlUO51Lmn0hmBXnVANflrvaZBX8+Fn8WAPZU6ioP
vOvyqsJiWothFfGmmfFOKrwMcqwrPZIvSoMSGqHAWVaKs+tCDKtDod0PoQ3g3GKZ
+F4+9TWTHTr26jKqMTwoeLyWC6YZ2xaQzIXOrBjdcJZOFn6/cW4PKyPqhyXvTwQy
s2NH+ybCmn8eiYS4uoVWlh2+8iP/2L/aSd4+c3xemvbW80opWkeAqKiyHYaEr7tf
KxBI8o1vfcC6V1wsxyWFQc98YM5Cxpg+3SmTK0OH7wXUNkrVnKmMWmVK+WyzSXJs
zSySFWnvkFmQPPVH6N/Vt/IvLw1K68eSQgtqgD8h6zmNnm8vVEHwjOxMNI6CBrAQ
fh6SUxL5Uunn5B67zK7LzsJ1ipDwduxl+wbAV4JOyHegu5JzAZUyzn58qgaqgBZY
h6bLu0dyPpPDe5UjgNvZ/F/XRWKDOYHid2DQRMxu0C0Q1EQJ6SGfczgG77BhN25U
mhaQoqzFm7mtlZEi2EW+kW7L2TW1fqv5qbWzmxGAQ/wlcsd11WZOMbR744Hb/8Vc
AB+u5liJBZGMTcVuEiXGXMePsaEy/lCV+Kiw6n0jJ33Uk/FJ4H0GMnGFJnhVve6I
a9emDcfPSjgpJPGgGFRHTcfZfn3XreVxLAR1Lc/tqoEFAtshG8gKNd67DoVGuQCi
LVG5Ij/c2/cNqXgFzZ5Nbk44lxzqiZhxWdOgtQshePDUkWvXdF6L6tPh8591jv2g
34N2+w62D+ot2N5Ggq8jTLjl7/lw6wLW79zr5YpEvlcAaYKNOwjZtcnSF4627q0S
91R267b2Q5swCCrsw4puGyYgSp8OxmxKzOI0sUqYKifRLIOhDSUoRIVIilVPMZjO
c8wbVTt+JnUK+U/hwurpA2rvu81BsJ9r8ldaw6Gmvh0+RLfd4yti2YJWhfxI28Fl
CaLjO9e9HhmLHIBGGpf4alRRRERqOswNpxOMXSKmvt2u0FyrD8CmyfB54xpC26AU
DLwSRtlWuG/rnefOs1LJaW9TxnLGCm2uM/5O9iX/kYQFm8rkVcqAnnIGeAWOsK63
UUM/Pt7GXZiplDFhsS6sGUDqCYdoOsWqRPYMX6i6GPUrB6GADYYaKo/T0cImjW6b
m0fjIhxYxf/swOY5BhoSeF5JjPiKkUxCvQIRYYlQA7kx9H5hMLebYg2MgbOG8dB8
sKvkGuI54+mwODDUG0Ufja2mdotV8vkxESUFU07zzPp69Zhwdr2HL+RIXeRUkVGm
0GoghMbO9ihocGrwXcIM0zH30OZMASt/XHdgywIG8WPQ7L7p8GNNVftrflJJUV9p
MVWzKP9orUOFa7QD05erGg4+dSzwqC2zFXxD9yOfke7JvmRxjjlsES3IFCs/d0uH
gCNqNVmdBW/mXRoQUg2zSbZ9aH4ItVRiKN4n3wgivGoHG106kAjdHRa+Lxcm+N/b
GL8lwY1xl/XhOu5SKV4Ipw90zEp3MPlJ6ziHmBq6de9pJmPHfpHZw3ZpNXqzjBXL
vz+gOAgDg5c0pXtuKBWEZwx0PVthslxCSlkTdPBeQK/tp7S/3JuZl7a9+iHe+hFU
3MPV5dfom8QOuBcVvZR2sRCd19jtj6moQFr1YFv8nNafS6Q7kb6J3Vi7Km4Ctaao
y4iczEfMJS02QaJbEN1kO/+QlB4nZ8ru5XqayHivaUFxDbMFgMRzH8Mqq4he3901
jkrZjik2unvzf3lW+Tc9OESQwWjeo+Erye5m3NArkonDQ6tM/Ep0VdNliZPRPGJT
snk4umVV63KkwT8WonF+uD9dxFHF2ZdMs5scDkA1hxEVK4j5JOjkwUBXXbXAbp5K
CChcnahq5Gd+IDxRHF0YtcYchvNehiaPzf5uTnGTHVE5gMxysy6gBOi+TVpMn/az
z1OquEyX3Awbz8NB8sjXEKMZImcortp3Yt3JZaG3KvzE3xCWBG81pmf2UWTcxFKC
+hL5LjmHt+ji9MsI023NiPSXxYTpXfm7JHk7oA1gLiYxHgSbLzl09gkjUjbVbOd9
tWjgVwyZwKmQtaX2RrHB0IZJ2zZIX6wSq70clGq9g50XIXiA5jH9wT0eXEQCrU4L
cthpKJKvHv/ALzJEuBbGNWXlUuxDHDRAhB88gbZY4x1aGnFMHqCeTbY6ituh3DU5
+z9JZzLs7U6badUZzO7mkHui96t7Oh+oroDGnLchmQzpzC5YhkmNJWeJJNBSIlXR
onmr91q0g4OAWTWckg2Vdod4GIMj/AyF2lY42tr+ZnmT439WVyiMYS3AzCmd0Q+Z
eBHta77SWRiSGBA5UvHVJ+bwPx/aw79qhlHn3gDEGWlMX+BTpzN58kRm0YdY1iRS
yKkStVuGiUvu3SUslSifNQ8W3+GrvAUZqpFGIbngn4gHcXJtVjvDx/iJo+WuQ4su
J7caC3z/ELBselwTqBxbjy5quvZLaNRqctM+P93eiq9x1PznGiBfd2t0QVkmhE42
BbPINWBVCBqN0Za/StTY4m/1eqMPXDN5qYdXnhr1j9fHyDYWDiFwTZrPkJzMWy+l
`protect end_protected