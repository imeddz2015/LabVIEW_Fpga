`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 14432 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/9huKRhRMtvnNqb3Z+UU7TahEoHV+T8U3P3ufru7l1O
3DlgtZzb9QxCbOjthp9+wDkjygH0eUfDrEl1ovhZG629iGXw3AqQPNMKZvQKCsdd
yUeBN0BvtpBmuFwjYFelezKVCAQOebHoYoPEMalffuuIUqlIEv5naMKTpfaNJjv2
APoUNM8SAkfic5Uk/qlDQ/8FTQ1jfz2cK6DmD+Y3p+uuWNfs5vlkTYKU7YRZ+Ye7
0z8lPr8czVABFaJYkDy3AIbCU8LoMKFMIC4lGzByQg8pLg6M1bvUns3TYn5XfZ/s
x+LWjYmuxCshzI+jeHDIqafw2NezfsdcyEPOPgV4GGebGQiLeBuk1KumlI9hsFh6
nrv9FaYbYmP/1TXP6ZotbLBYyXeksDl9bQNdVZNnK8XZVM6m9TOJAnzPRYds3Wme
ZZLYXL8lEYS85Etcwh2Ds9sy2bS/W0ee/ujzAKiwVTQl/114VyWMYVHYBykppdev
/zubYz6d4j43NzI8xxjZER0s0p2PLNDyDXDuoZoXWG+eD8gC1D4v6UJhlTBOgIsv
6jjn3xuBDFWpycDQqG3qgazu4YgtYJDNAOMOgZB+cyXhQdIh1oRlKVh8LlcuaGeI
WHsCDAWJTHqkwszo3OWlzYwOtzJEKBgjA/eotVNSq6vSzEkwgeENYHTTXuhAs9wp
pU81rcgIbRnA4KJswppX7igK+dwIEJUIqiO6/6feZOOKk68av/sji7xiNYron3i+
R+fof/6a5bR5SiNzVcGqgGtuCMbcNJRfIYsyVvQDS2sm31VNihBmoUjjjUnAQw6O
lR5ovdAFoTdtGZs5Pc4iKs+FSuqtNMzaeZcqhIzFrGuxkT/StN2EaSZRGTlxIk4z
s479eiXPVqW5DlI5mhpJT51pyVj0QKsCl4dydE4DFdEUwPFjNiMl+dLXPFkJHe+m
XO1IB9nBqW5UVl7hHDZWQaHn8MExk+j++G58a2hJJBFJW7Enk7y3zmByom61746K
d3+OrfsXu2HQWomgFRemewU0tOqHDSxhulv+LNXCL7T4JSiDyYHJ3n1hsn1b72k0
axd3iqZAOvjKCEp4pWAAIFW/CDmFua00nn+CaMZGXxrda4BTNPznm3rxAQ6YrBvd
xMUiz+PtVU46lsAmCuc3LiL2Vr/od6QbzJIdEwaxCv5RlzYYTz/DHZekx3/Dc7Fw
s36JAGRzjcJKrVHpubmdxyH5q9dlmjjXY3MkgePQC4dHZ9wLYkk/m9xhybBxD1w+
JoG/9yugPPgp00IFtmmbbuijHbIrPBIcYgmTZO3CknaYkC/IofAAafBHameJb47v
VW2O71WFvOeIz0cCkVLE8KH8nSp5qP1o1azKDGYMeANQr+TZ6GSS1WAItluSe2Jw
fY5OaswQPzDp04gveIp8HzzvJU/Y1SCG7Nr6+1jK3Oe/MX/4Ljve6UhfGgPOk8k+
p5cty2NS8t+Q5VaC8ZV+6LK60e/oPlGU3RUTaH8XyixWICqZbEHyCbKhjw/lU9CF
5JF44z4EP2p92rMMFmBH8aVcCdWbpsNWI9E2WT5slGSPw8jy7LQ7MeOTQd0D+wcI
X0/JmkG/zYf85E0mItEiecJNUiVWzwht/WeYnEgqMd5ks0e3cZ5loY7Ng4dTcI4Z
5zBXTE84IaCBi8xYU3hrcEH5bOZkMshhKLwEFYm4DmIfxNwZRnL09w61g/JIlSRB
vVXuDYskhtdmDGo2M3C1d7UubY92I872hclC1dSnPT7RvH1l0/W480mzw97lrgAz
i5bxRx6upPbYI6lS0erwjZF/pgZMEd9+I8hjNKpB1ZNeqRmDGIJ5pxSTwca7xiwn
wK1qNx0CgaCfVHFTixu+Ll9QLp30l/2u/K8aQqbDe5t1mjMjqO2GUNue+o3X9bxc
Qy5l0pQzwD8mhz+JyfkoaSgX6YwJ4mX4TZR4UIxuAU8LshjvZr2JkdfYuL24AmQC
5joATms6SFo9jg+PQu4JtymcZ+VAjEHoS8xM0UjU+bcDoSuAV5AkkbMqrGKAUHLh
H+UnYymJDU754wfEhakOKHTRFa3g/cwbamsj7R0aDYsaesKZ6+ma4aATYDYd2zlG
S5sZXqsyIFQQMuDCJ/EZLxiWyCD1UMBIACNMabMH8dFSsh8523N260QCIuufBRX5
LGy9nUlU381sKwUftoIDZiW/83Em1XaV2n8aPp6CWezYvU1FbehODVuMw7hyZBc+
6J7kUD+FmPP7R4EuMdKcjGeCv97qfvyTLs/JQgMD0uZn99vrcgNxXJ2aX3QFnxQk
Io3OgFBjIb12WtT5H/uiTgB3vyj8M73SI/BVkTLFsF9Eu65JEfKLQfrcLDeWrNVf
lgkOWyjPTeyBL6sK8+eIFViIaabbDRXWSl4XKjQTawC1IsOEtmhOX8MpmNZuIyts
/ISx/RVC7w2ekgqZrJvD9hFdY26sb7rHs9BovNR5WOFWMp4UpJhqvF9/CmFp1JRK
h4Iot4VS1cO5WCNkyeNIxpCjWF6XsCpJsC+SKSHH6uZ0W709KD2ke3bv0z020EWh
aDrsZ49Es9uOfqUcQF25s6NQ9GGGhFM6ayzMv7QnEip2jwMT2WBwdNASFJQYoGRB
+PmMuB+ZycScZKA3o6JWd3AleyLrZJBHz6omNfjdNJZ8ECMsTzs63kC6i5aTRmP8
Mj/bAc7mwEuNCXseCv6seG841smHi1e6LZRA8SQeB/uc1M1sq1eSnv2mTYsoxK+F
ju62iU+u3RAgtmqBmwtbShjEky0SAb1+WYhoHlizsb1iF8hmYbEOjgiBvNyCoNH0
RTziz9S04mUtvIXkNg56jLcciBwNG9vQJ2KiMNdp8u2LOiBhq9NUWwdF27EzsgeW
uslhhDiSOULarbLp4ze1/SUmjrhf8ZRP0wws575WJy/gVItl86BWJnayQRgDT1F6
T0UoGAZGYcqWUCNj5N2SprVUxpEz1eV4/Z6fOHLp7U1TnQeVHTT87UGsAQBVvqMc
HMWRls3YJ23d9wRnbdrYJD/9NTZKj2YImFI2rM1sUxBT2UChRl52qTAZlifuqWQx
8AsAlhE9H6U+KmHD7QRaAhRpibR+2s4qL0Lto3pqI5dpELAIdUFcdd1JGQ6Iec6f
zq8qw0px6FxIm/dE1PFBb9T5kwylBa3Baq50Iih1xL8vklFClzXaFNMqB1bPudBn
1bueNl90stPInerO4QwEliSoWs/IPiDEyfrLzYGQCzSDVGGJQOypjDIG9tLgQ4oM
WbdZ/IDRmjMgLZZktTS+EtXHVeKCwR+Dt8g3uF944B230WzXQdxRRBU2RUIOiTbF
F8x/ETu6uVyjKvfc6vKCK7e5gudoGEIUoc1Nbu/oZkxf657T6FuEkyPL6W+C0xTI
1G9pl/4hdvRLay5Vjew5q0ZXmBqKHA51w63P0Q7Gf5jgjoAWg22akMADC7+VxHXn
9ClpeiRf/sZCRgURbymoEZ2FycBWJBJntAW9V/R+CqRX52cdCzwXSzps7nThBF/b
1QFaPf1Cj+KJPWki1O1XFJbgZpy+74B0kwGRxfxalNJk1LwQIAd8iTHEUeonaE5c
rQjYhpUwWAwf/j669waIrUz0dLzqL4wckTCiNSb3pPRScV2NLtbnb+v1mNgoQc9s
7uqedlrkELZBlF14OV6rgu7Hh6Vb8HSU4FRL2QMnsyiDRw0JWc9OVVgcldQ4jaPJ
0JEP/Go6I674K9DdZwM7V/nL0IfeEAqhwhJfhLweQi17CnNkciaUx58HGkz1bOJG
zzQFCzpu2u7IJM9HsY8hMXlOsk64i8VXyZM5CWJOPakjR7NAEBTfovO2h1ty42HP
s3vnX8A6aKZUX8m8kyftYA6CrBnMtJIrMDfrHm0tANoSbNQAubY9P3gW47XFVp8g
U0mBizs6hisQRfWb0pOvX5qO0aqwCMkaWZv0EqJj58OC7T4g9DN45/4vJl5uIXVd
W74W5VAq3N04Q680azgHPAZeej48b8zf5v/86Kq4uf9Q23Yy+Cw1LN7TDQ3OFTFS
mLZm/sQ6JEdeFHrjy4n6IGqjFn+Py2riRQbAqC+71n1zQtAeAzeTjdPJu1zp97J/
Kp/MDKSW5EOaxx4Cz0uOHpu48lrsPlWDmcc6ZwVuxp89jjeyQP7fDEz1P5lL9EKU
9EyL2PsvrjXl9qowzKk/97RL3v/QhxApgtCr1wJ62GUfm3KrzblqU5i8JkYjf+tT
xah/vGWvK9w5x+gxVfLp70WmhdWz3gtl5RUTPfLyDyurEf44W7QmV+JMGo4sHStx
milzPbJHPYP6lRWoviCTJRAI/Py80mshd/xlKCoPqN4p8ga/UuzxB7pvMvfpstQ7
H6h+eWLk9jSw8SiASlY7xsXcvgbA7EHLTPH8sImldxP6lQPBphRfTpFMET9B7rd2
ycGXJuJGjSRKCOrUbGZAcUwlDoj7f0KAZ4bGX+lYxEbRTJY3vqLtmD1aQlNJwUVR
nFkRxG+PlupKEsiV31aHM7u23tyUTM6WPZEj7vbX/2m6FKc/u0ulCiUVArIOVJjU
Ye61yvXt06GtVuVMXEWKn1YfX/I9m4v+MvzeHaU9+RzvqmrVBX007G3zFcjZE/yE
yi3EwtC6TVYh0JFqaYz2vh9VCNGQtNNPOLTslgt5fEYQRND6cFd/ePrOeQFeRtsi
VBLSJu/OLLxz14tQxCriZSFWx9cIHSImW2kPLP+TFeMacyEwNbZBg6ZNXD3rINSZ
aymq2HaGRP4I3bxGcPXFhudGAm0EEduC3Ylpayij27HXXEBVteYEFg7tanB/z/q0
BnaUAZpFaTOvNHuBqFVEY5sGme1DC58xgXQKq0F4CQ0WuiXU/tKaAFpL3TGOa7d+
aO2nZypiDR3QBdge0ddsyC6Yz2N4IeecUmGY/hyIygpsRvsUoonUU38CxRFT6KVg
mqG5dMqWhU2B/eW4Yd6WUDXe5WN67Ti/GatIuuZ9OF4bkO0JXjooRGTC2c/XUZUZ
zfcDLwEU6JAGhgiiHSgVhLRx3G0/Hcpgeikidxnq0Fo2AGuA+JGgqskHUk6x4qD6
wF2zV17wG26eSbquZlTsW2fYsiMMfMcV03DP6qoI8JJ+VJ2Ute8dKe43luTdNstP
6rglwcq3lHool8GA+D3L8+7+7j+FS6V8CuH01MFHHR6077g/JPRZ8DWbyssHBn/J
86Wgw6u8oN7dSirQQ1s70EP5RNfydYHIHgPZPlzRgBwYn4t8HxPkQFaKwPCdrne/
vpMkCSThS/SAHQZ/C6D1RXmvirNJIL0QJMGU86tc8unZgFCx1pH2vVtNWTQA6FQn
r754K/y0dzgaJN1AKD08yVfXPO8Fp3gW0MjbcrQ3OPqVWMmK+ndWFfwmAQ6J4M33
k1OvJj4QPtTSoszylazQEvjVyPAoSKoKO69JoCZgqH8aZQ4T9hgbNRGI3tKZz31x
bASRvQQ7IWgJ68E2031KTimWTzzdIwPmWAr7Z/boNGQQWByxSQQGRDv6sp8iFnTa
plYH7KdokpyoHzHLjzk3C4A1mAgEd0w3WpoY3gCB56pVuvJkQbCn/d8EWFtJUIZL
PcKJuYnFJ0kdrTMusHt9HarlcP0qixw4AhK0Rki4+62SfCadaON8yV+/jPI6o53H
7miV9hPTNbd+n2MGuYTKODuAB0xIBrZtC10XpNPnpT5D55YGYDhCeWz2z9y/wm7B
unsI36rqYQPpTtJ6ooLdYYmfN+qCa0AZSlsgfeJzpH77fyV//LyV6soYcaRTDg/U
Z9sp8RfuCKr+svCnjlZFIYScbNTtGmBFwwlGw8eAx0xeMoXBjAAEtRjTEUNzDFH3
XeZv3+RGoppCCt06/a8x5/gV6Qcgrnav4TqX2DrQ32E85oH1C3cytNdAXDoVgm+h
lF9wkPC3BHvkG/fZHilSpsR1eeAEO/fOB2g6+M9kF6+9uGrFjCpn8j+BGpvMFsuv
RtzvYfvYrSGMQNDN+n+FfriDZwjd3BQE5GQnYSXMEZJo58Cci2+ezLZxC4W/DIfP
0rsGGvp5mHN9SHgZBTmWXqwoKCAxM1083xYv67/JSxouccDoT2Rtn6tEJXDSMT0d
9A6eDgr0uSUUE1kLw/qnBqZQFan3FV4OFD0YEJvlRWsF0+Atlfa6yBayRGY/IpCu
DPmQPkj0uwBkbJG4vGQqnMXpsbhmsKNqn5kXmlG5bEBOsNGowALMS0CQ5DZGWwno
NTL5d5nXoIrV8wCu9Fv8Fk1jjJC8XZo033C0mrty9f4uxyHokYzjtpHdYJJrNk/l
0yQMBFZpWwPDCzX3WTQ7Cq3IW+YhZ3kxrcOwY1KCaqkQlZu4TTN4sdk14bviwLJ6
nDZvXcxImajcS5MzDDZOOn3PfAVX+5/YZXjp8jN+JpdAzAt1o0keDWcN/sZgE/Nr
OzTs/peWi5j+h73czwWE3qcJbQvT/9hv8u2CVPlTN7TfTf9DrqJlk44svhT04J7W
MTBktdiyk2uNZm8FePQW31WNdQCSLtY1BwlslOl70LWMuAdx1EdKgnTbC94zlK+V
xKNKjVz5y6PVfgSsWEipyuwl8RlNoNto3ExQ3mlq7LMd5eVsYsgXptNvOY5cXa78
q/2THtCKG3YEbm/vMpGjSngENL4RI4HDsIkfDfVzLboxejgKhfRuuBAxiYGpKfvl
gzspry8SlOexb0GiSyU3DmCFhjat1B2Ez0otASzwvkAAcpGWLqwL+RoN7VP5IC42
F8b2YywsZq6EkH9gFVQ9P0rlW7MFN2lPOfeg9J+NHK9987vSwkAABACRJclT7mcB
dviajpIRE8mC16YtB2nwL+x4IWIl+c6aawLoAsW4rYZ+FLyocmoXnHlSY/uyTgFw
NixoeTm2sNDUMoefbRdXAeADOpHw3dO0G6PidXf4YxvxOWVNJpbXGV5SHm7ncxRi
GyiKyANMzk/KWuLz7rptF2kpmX+i7exWzsd6QEatWhgAjNWBO7bjeRUorB2zML7i
1G1cI3WPPs9iAB/Fbn+dJ6/JA2po9cdaONXKSzCv0Xijx+2RYvXW+2lR+Lgwxh3r
JdvSbpME/mVoY6BQ8mmBJkng6quBip3td4ho3U4R34Z2sDWVYR3hkNbGWlzWZw05
lKmO9v3Z/ZWFzPgam9jrTaxprSnfBv/w2bnda6GqxywXiKmBGJv/JRyuX4a+NBoN
02hdgYPrtJ1EuatINsJ2X+qCyKzHIkixL4k9u14davTOEeY0ALJt1ROSQHGoa5bH
qVhPJnGun92GFtitF587qPYF0xMtO/fFEScboalHsAJQOX/geszaqyAWWI3MwQyP
EEm8zqdA/nG0VKySXtUey0DVNS2qhv6SLoq08sy8JA+u2ZZD9RHZUMpGcYDU2N3P
NO2zt8+s5fyRSL8UpqaaSjyFAa5lpQ8Qd0FkQ6rWBW6/daSQn2jHmkrhYq9wOwkL
xEAPTOvaWcOTx8Z/3KiZ1//WSZe/C/LYDECJXY2t5fAIyInNy9LgTGH+25GJTvxQ
YMpoj2PPQ7mrCpANNF2KE1DCiht7k1rOeUTtSTcb6lctq6tWFWz612+dHCnwNVCl
cOhiHCD/9Gk2bTf9lAkPClxcw6da0SQoHy7GTrGrY35Zkkz6pl2lb8zyN9/50vU1
7sP83ojJyJHIjxlaSv644o4AspSFKD2ER8AGbBMyWYi1Bs9XWSqGW7LkIlsCk9Zf
KM5w89fN9qGdxy6jIuT1+b8/wxD6J/6HxFtPkI2zzrtloxPwkdZM9ElVj/fwdTSi
kYgjaTZAJKkCS5Pa+IJLCkEv6cnn8L2TTKsLPfXFMB1lxZ35vmGJm21ZXInLREZX
6e5zr4O6hhjpFL0p6L+A+Qcx4Nl/WUNvZ54LeHDo+5nDy9Wdw9d5gbC/yaT7X6+d
Oa4JxMarABMFS8EnvC/Gi0LOKf0Xwg5GqRbstu+dPl9MDmKH2P7z6q0lT++/WHHn
8i5m8Ku2txY/GIiY0z5QqkGfkZtIuQ61N84Q4mwoGo8ToBSiI1Fty65cq3pquIvl
G//hua4YmTYIyTvS7ajfez1VNVq8tLA8S9b1Z6GTxTIRWg9C1mZz8BgaYy5AggPk
rhqoTg7M0KK8A1bVr5HdLY+CsUJrLCisPkM0BI5F2kSTjjRpy0DP+Zmd2ALrZHII
kxOOqQ2HZPqZJg6bZ9v1SiZWQTJTCiaNBQy2XU6bQkHYIi4nykA9pkP26gDGdYI2
Db07ta94T6uE+R71oe8s0TzPEQgsn7CVguBWAXjDD4G+l0uheEJwsHNVn48ya8EP
niPOYlu99ivs4xqaJXQzxJdbvsQ9hPV9TV/oCdeHL6sj1VOpM0N/VyN3fEyeTKfX
YRCh8v3yy4Qy0LeEeP35zJiT/mSjyISL4j7bmdWWVIUNlpoRh4UTa0bZm0SnYgJN
jP7U2g8PpXtFxPN0f6BlMU/xK1GmQiswRk4IM6YG1CzNfIXYd4p63saevQGh7dGN
Ezdif08QNFoyX+U7l1dOJrL+RVlXUhuaj4sbIZeUu54VljiXW/aINbWBPhBtgrB/
kasmF6Av5gDuyBZZnOMHq5B9X0S5NkpvHvQFFeSjXEwspfNoJEwbGMkQUAY9DI0d
iEYxH+E2Fbrc6UAc/OJiSvr3a+Uctmhake6o/tvDBGdqxDRNYv9eV5EsskeprXKD
hxbmTnptsCI0sIfsk9hN19Ehfz+vID3z1me0kGaSBNI3gyyxEKIqFwswOMbfnNU0
WxEomymqNloutCavFZHrFkf4+FD1oFkHEB1kVOja8+G0AUGO/gr0weYRRl8GMQAE
wXo2BP68mOw/FNVS2GCPKlmO+fYsDvFS402EtiXBOPCAQbIzCDqICWv6OiA62Nhg
xX/LWBvRZNJoHTD8PoDM3us963qqNLqJ9Dsc4bybuQqOVGyqa4eK2njm3KNZIW2d
2cvuFtFhvEX/Yj4aPk3ZCu2KwLAd/rCPfK+uyOl/S6MecqaRIkbb+PoVRymdtx2d
yOxlvmq4OxdURTxEklbBcIH9EAa0qiyLs3uPtc7u4xIsnLR3R5d0n9txYG1zUc5O
uqzV2l9HiQv6/oDDmDmFgzPWHtRen8ug1W+pL6oHP76aYmW5lgY4AcfG7j8ccvC5
Y5+EsmCViWgMZ5Gh2AeYWwu+Hv2EiwX+Me652OLxZqRTVFqUcizenxtIl4Wfwqhe
C6XTe3Hk25CFVZSeKb+QEY8IkIVPLw2OHGZGEXk6nZBVMkzbcQLQV67+Xyes2YO+
VWakfaMEzd4BLu7SmT6PRQU0RqTKH0c1agDXGoCRdDfaQgR7kn2ibK8nnBM1nn5w
aEhlNqCwz3ID1bUkRtRejXpC5JJ6RwcKrnZhvFLng8mORPfk2GphosfeXD/RCzqA
qN8d7t2s/HLoqCJRymVgEiwUIJEL/acEAae5xoHCemu4jCBaFT1bXQ+LtYkOqas6
GbCY7SUd+5iXwsOHgu/Ioo/CL+wu7KlCU2u6EUPGqvlCi0Nubh/ACSLn9MatVkrE
dDf7Y3cMVOLeqvzN1ttMK5J+15l4gHuOLiFHBi23GToR2teW9tSdQxTkU7jEWOF5
ig14d0IyUie6euBfXeT42fCsnyQEIF1sqaMcjzE2oLOND461s1cL5PlA7WjdxCBK
TtD090fTNdOlChZKsiEcV+er2XbZGKvtNOvBro4Tj6UMJLft18asF6x7aK1LLTxL
LnWbmRiB9tTQN599zk3UFmCnAA7sdMLJbLY6ad6g9OpG4NW8NcLYjFew072oyfPF
EbvxMsoA5mmyVvzMtEpdseOX/+HZgA22EIWrrxZFAcih9ru8opPcP/5iKB/xXf32
KZH4ykvN7ZDVf9q1jZCgc4OBNjeomesXLtls4sjF2Tr7FB+PEaRR6VxWf55Qt3Nt
DynHBVuAdr5d38a2rdQZx5aVKIKr9LpqPH8YmfN1gyxuLwLUQHXvvTxP+Ss6IBm5
digZK/jcE9qe3d9/w0WU2tTdUdgkFxhzRjb2b64ZwDDV35IYYjHcpXt8HRQiyiSs
qkuaOl9j8Zayz/3rGmziH/PMXzpmxha5CqahqEPYyHzshug9daC5TKRkUiqzfJEo
F6lEaH+ClcCUn7Z9SzwEwvpoU0x3dwLUL5gN/dxmaGJQJpqaEo6iGDq2gjt6vePs
UAIjIE2aaY33ArQETna0V+4DwtyMixfeA1ZLpGD7pFtssycRhfp55UvkiJNe9Erf
pNp6TlnWuhtG4B3Xr5tKJJHgrsjCnky83L66YVPuYo2Gbr/bXxys0+QzMFGVqjCC
XRiM7R2QGNrZdtYWeOU1Es/8zsUHUeqPCp0KmMZN8p0Cvgt97M+XRFxc7Vx54lYr
6i9t61ewSP/836Ua7KQMZMvGmhBlDZdBHzT2F5dymlHlEgfq/kfUdNs50/7EUQLi
Ncpb/GatF0QFTwV+vFYMEKd9Liw3RqvbubpEw/Xc5zdLdWX0ooyFw7cjdbz/bv3E
4d4InvYr2UCsyq6/ZzHCNn1sfAkdo8kSgVwJi0SRlwlYORKF23oHeDnIvNzqKO41
psfAmC/gAkrqYUOVb+XVHwdp+45UEhr+lTObwgFYaKIqVMEztaAhThrDE3UJm8c7
6GmM/QHlqUi4VYDR+VlsO6YtxdBJGmiMyZwJ78Mg39ICwsdvlDNZq//oeeJELE42
YzmCb6JxwDJP+k02W0eddBO6N2X83bSNIGBWYBg1qqju9pQmcLEhEvGWYqG8KXTX
qAAonMFzhdpZEWSkH9RiqA63Yfpw28YYVreL+LnvWtb9xjZ61EZ4Fo9+lAmcyAho
m/llwX+8DueP2dX29CuAsbguuQ7FOQ2iTJnY/lTkRDI8DnXCdvH8RnlDEYM4T7oB
wHb5Z1Z/6zP+3su4a5aqVrWgu2KhpfnPq+1RwnEyQ1Oj1HR/ZOMLD94lBsCotaOP
6PIoDu9F4zokabRw4oJOkp4gysU9XDpdmjQQ7SBo6FVlZ4Zg8btzrs0gVddtbCZj
nes2HPHHMfJ1ImTdicm/Sh5G79euEg/32lYUXC6ijne/8ymb2lHxjK7m3Bj58lPc
FAm2xdrf3+dI3tb44rjBrxREGQu4vgspQzQf3pdAFs4FNDsvrahk+Gf2p2+8VvcY
IudmX1jFgSN4L6qAvjL/qZ0vMtAZMfJWeh54SSuGpuU0uYB5a0yo8dFaVpSxybrq
9mAiQ5R40YZH3RA9k9cXlV2nveh0eaq5XaJXKLwbV+SmUHDl3UpUmNXqOZC/84w7
k29DjiSxWWoevXEncBwCqa4afTt4ZuvTOePySpY6GKP6yuy9Sct1g22B2hZfbdKz
C7qbIhdqOP5bmsLE8iSpWE5V0hEpTIYOD4lkomrb3n4/eanT1gPWCxG0WCXuq/19
Uay1NslRsBAFeb5wUcX6RUKNFSJSTPAJShDCVMgIq1Z+k5uhY6iRda2Dsmyoaez0
0Zi8iNpQLNcgughPs9xh7YGtXcpPJzs0grhaoIb695FGWSq2x8q73M7+jzm3tGqd
WTEPQzTNxaZ2ERmF//SS9R3keSQJQ5Dcegkf/TYO0HK1Q2POHQLcUHwswEezLd28
5E83A1vR1cohYdcUTSRuebtasfkIktPLBjFXHJm0stmcjwPxnQx2vr5gmm2c2L3h
6Hx0veEiV/2lYyjyhPe8m1eVO7hpc25SHSqxb6Ph2rtV4PSvFlb9IhsN5kLw9TDw
Wx5d0lZhNNNJa895ocjE3iN5rQ7cz959Uv7jq2AFEj4HPD2BF3b80Ww8r7oW6Qpl
H790FTR7T+aGnCLjJXmSqdiF3u6+v9TMd2z8/+UZpFRIl+9JsE5YFNhWfu3Bh7jd
5K0t7g0+unJCdPGP082i0OwByqU1WS6uSWUF3y5j6wk/cWdhwZ8a7csQ8KxFrIXC
gxLhDky2j7x0ybCp4eMLGcP4PErlG+SzJ/sWElDLbK1VsKwQKNjxAhXtk9GKnaUM
tML9b4xoJY5UPeeaTg4q+kv9ME+ySuuEIYlcdPX9wr0B4X+xIV8uARBOBL1C7rsd
5ZSlJs+arq6uyhp9GTYp5PLAKavUXASa/frskOS8WKaqaSullv77pStO/YjSflDD
ZxbOIAg9aG8DGvO/oorAaHenFosZeW0dOlOJES5GHsMgTaYskjVETi6q0KLIpq7R
yrY1W4nAV8ZVRrbRbs1DWXJ+sbG1Cu4FvSz2wPPmZ3MJjTtmy8F3+1AgO6J4huzw
MYCZVZHkEbsP/PJLAFCTgi8nvWmY4Agv5S5+Mh2Lum2Q72r3QUFQ7eJ3qJmG2A+9
Gnz1lUe1wZgfQ8Vye5zGIRK2uD+r5VTir5M8sSGEM2Bt0zlhLpBJrZPdvMCZg31y
eECK/TkdNhdifUKVvGyR3S6Mga16gj6qWWVQD0Qo8AKoXW7XF2pcjCXkdn7X6V02
RwZ8bHKGGflxIDmBtVOR4BuKORvClaZOZcAwVIYLM3qmZTx5QOkRlrapSHMIB3fH
rY6g1H33Hht93qxdmSSdwsHDTpthPYYcbpUo+kqs4IrpdwUpXurJN7J/xm2qvhMo
a+v8nsodtSIy+ooTHWqRDpTfpenVRYwSjUGPlzl4zjtoiS4JhLo7rOb5sQfmPtzt
41ovqh142/DiC5+0E5Yesl7PHsYWPgWU9s1pJsG3VRQUJidkoJfl15n2ELblfGtu
x4b2kVAdgFcLhHTW8H/SnxRluqBO4ZWZkoDm/ua6tFRjMFr71CY6rRnwX+r7ly/c
Htn4mOqJZhF2u1rUFq9ptKKmMb04dDOsfa2KwG8NlQBdGcTIIvxDIdTyCB1Ls+i5
h7Hod5W1eUwp1FxoQH33ucLfbMPJDeUMS50+zOxY/4es3exhqcr38jiWaXYE2lEw
1NNkmaoxdOynininSV0lLeP6JYJpwt2xyDPmOh1TRc9h9EsA3rstoCdxwvsMpBS9
RBIAxyYi6gGs3yAH+MSY9v7HQeP6qPDYMRFpbmXu2gr4PqZ2kGwjG1uRTct2kL0c
Yr4tK5wuSumve/pY1U1MAYgJhiZ+tqHykypyoF7wImeg9pXnFnQf3J3yCXiESZge
naFGNZz61qzp1IcLmly13h0fny8QDtj0eutOk9GKgRis/zg0nG3/XkQld2f113VB
JcwoOXLNH9o/aK4ZW9UQZrhvBMFy0PVQW4hMaZ6Qp9Q/5gVM+O2NAlVdcMbkkQuO
BoRyhSXGZhefsqBk+nzAyL97Y4meDVufFPpE7O9QPnvMaVca8YC6ZWmxfe/xi7ON
v+yxnJFo1FacmEJen9bPxA+hS1Gy0fz+g915DLapYGkNMznxOpWm2FV5NTPSg3Sw
+X5WZcLmq5yizIKKS7vn+7HiC7W+OVzl3+37HqyXCjDgLY8YEBBKiX06ZVdc967M
Ed/nSYjQx7VH4piD4MDvlJPrH08wMdU8vabnBehtny301ylqSE/PrhuEysD403aW
zzHY2VCICKrU1VdFSJMRY8edyShS7d3VHCgBK3G0lPIDciCgINUhhpn0Z578QkLc
0k3zXghUmp1tDrtCWQeXFo2kJ+Zrs2EESeS3oH161NnjwBNjHzMG6/BwgWir+x+n
HcZueF/gP4dMkAE1Lo14QvsAn66UcrxdaJpLMQMQX0z7sw18pxM8bZE/DgcrjYBr
t4IRJ3QlrmTdbJw1TaZu3iLdadu3ZF2oIZPil3YIK/Kv7AyzgQWzinSBGKdUykkO
XlIMHejOLFcG8iXHCWiJsOnYsMSNT86gElLFP3SIyGx2uiUSKA3E6ep5Ah40wpNZ
eqkBM7GxaRLVpITOBVCxLGDGvyY7lHlg5Fk8oGK0YS96g91x0l4LumaeJ1p7oyuo
NwsNW/1TIb65rVQIe/7gkoK5dznO/HBTK7BlUnPscdRjqyxLj6FjWU84nh1AO4Ef
Pww4hqVi167KNt6WTsNnLdBIuQKBunyLIy9/8b1Q/nKJ1qCOP9E9yYFAi6O7CIzf
zB8SycUsZWq+BL3O75sQcWdqeuybJgBKBaR3V+l62S3GQA831EABc9Jif9KGYRcA
4sGXmcwq09ocR8tAIKZ77PlPXfm2QQ2HkpmHGhCQKZwjh6tRhbqQy4+LqcKEmtgA
jOWcog6ksUMiUNgitYBELL6rP7E9AjPqabhMvGJTce92jwvBfuKJZXMkh7nqpZ8c
Tkp6AGeFLdIrSeqTXdZLeoOeOIEZwePZoyCwLd+4NGrCYMLhXrRDylo9nT89PGXQ
R3koshL63tEsDoPoEBA4ICIbxYgZXC2ofDhsrS8cTwnCsip+G8ZBNa8BQgRV/JXl
PUmdBbnsgZOUjWdk+xTk4T3DEfF3XmuwK1WSxkMFRqZ/UbSccls2/KuPROzYh4w5
xrvuSzPK7KHKoM5EifSyTkgXhS1YvXsGG/k4jVqq6bsJFLyTv2IGt2P3CbC3hR+c
CAsnWbWtYFCa4rXaqGElWtZ4oHCqLHLOE5Pj6VzMtCTFUYvOEUPERK6XMqlRqum/
27r2TF2U4oG+6h3LDV1UNV5xPfzvDlnRPbq70aUF6jRa0+T7z/87/PlVSvMnxQLl
ByT58oHP7WIQvBkjtgP4MOjOfTbsUSikTKf6NsmBqHAyvhwC+67LrSXkwmrBj3y7
Vy8lWzgSaft0fCDRM132d56solxtf2RzdNJuYHrIu41Yhm1z4m1ZzXUP25rwAfPD
ZRRmKvMKJtOKUncbB33y+gCdlVnUenyGqtPDgho/+x9oiyaS0QLmP/YjIBlye1CF
tIfdtHIh5tWFrZ68/M38OgOt4NE7jEWaneNHn9qsdVfj9YOOHXufw50Nuua5DK2b
YRc0C93HbYpU8lLx805Evd6HWG18XY5tRi2RJp3cpYDNSwj4w4F4ew8hr1cSn3kH
Mxhqc0zSbiY+jzA/rS9pJF1jK9M2zMf+I/HSonDdmWzKI5Dc2eOIaqI9pJv5Uec9
UYoskzs8i7WuBWnp7md8H+A/iXZlyDM4QxfPNPTb4gyJTZpiM2EHoAi53MWPj6w8
vFvnjXi8EO2Ljjz7jnx9ouKtHW85egegsOSamOOgBb8VaLIXGnSe7GeKRPnE0L1c
GiZUQV6P665dkBZh8nhagR85KH0CCUpFR8T/AN55NVjDYxRKhrJPHOLt8yjzM05U
Qv7Q8eGsbTB+VjQZpYuuutQB0J2m8bqidXbhNK8Ll9u3U4BDvlYNlPvz7MPN1XTg
0aGtyL824UjTCtPzydX2L5PuqLbXUBcI0SwoPM+ZkKdIJsgZfb/dM5badc+2Hwmu
7Ln9RvSZR6x5LpI1HnpuKOj3F6kW7pqgKdYK3JG8iBODs4rWzv+Ut7E7E5sAaj5u
f4E7by2Dr6clGzyFsvQr7e0R6tZUqSXqVnMAW1x2OtDHKdx9QLACCQOcG18pJqMH
Nz8v0e3hq3v6TMWwyWa5fj7fWzNjOE03a9bMDbxYEt7UuCKWwi5+xByshi/B1XAh
QB/+HUzo1Gr6kunBDA8KqXgx3w6FPZnEvckMQOz3fa/V2IehuRAXTgkSLbW29AjH
Cw5Ajl0IgwSvPSJgIU56NooDi9UGHy/w2zGSpS0cTBG52cyJsSCky6RYjPNlYPom
HR0eqRK0cqGU9x3mDLWrCmWptlKTZK6yTOtxedEj115Yr3IHv6SQKhZN6UlRVrhw
8Sf5Yxc8cbUUlu3BHspLJuC6X8jBfhB9hMbzoQlpMf63jUK/UEggZgzKJStK9zJP
dOR382J9PjhKaPg7Qne+fS5Gf75R1QcHnw2ARaBh59A2qebSGkSIAERdT4F6/2J7
S8HSny/R4ojAi/kZa5dd4FhIwfBtbcpfeBSSTW9Y6tzdIFl6cKbW6RCj+HVzNEEm
NHkNhzGOsl5SatW/XEr2TEyCEnMrYhxoTfR//BBosam+cb4bRGqEc70W5rE9KLXN
xTnk6VpQTPeinNEOmvOxEYCbQblBMZ4S/M0GKqk8Uy5fkZm8d9YnfTKmcInkFRxt
LJydRv6kLC3ELSlVy/msaFNkNkagzRHe0S4Kx5Emp/C6Lv2o9lgBubv1G/16dpj9
GuUnmTph909pA1NheiuBFQHjQYXurlHECG/wC9/fQZ14U2ENREUJ4NoURpOeGrk7
QOYB2KWLliSZUfcTbh1AMBUjbwkokdLjwdu3f5asjXD2QIAI/bl81NkKEb5f9DYS
7n5pUNEzftD4yoOZAeFkzIINctuNLq0+AMbXTyP9OmoJWDaET5x98lkXSNQU2FCx
xHH2VNXkw6SglNktEQhtHJg7BozIHDAgogBJBo+TyV1Nqh+nrcOp+Fk/tSRgAdcv
8Opi2NbCXw5ujq/nXdpbUUzAuNVxrL6PD2LbDm3tCHP+p3QvtMSSpbti4l2yfdhk
36UXK3CMNFWzCaiG50BDWGi+IHGI1KQ+pylmc/DopfMW0TE8U1ZPBE+3v86EuRzi
XTk2vLYe6+ZlT7TqDS9mISKRyrSzyjJVY0zcpDW5wRYVAYce/1tgEv2zwlXR6UVZ
5ECXUl6lXbHOZbyVejlqMeuzVH3zBw6Q2eeHKkVtA9d08P1AGTH4tqiRbSOUSmmK
4fZXO3jqE83I6BNx85OB/cLu+Vqe5aWpGYSt17YFzv/klTMP9Z8GnDFez1TKDK3A
s/VcXZvL/m7VXt49z9LS119mCjjH7Qu4FngB33CzQZs39TuozNAb/ltIfCZ9aLNM
MDRnY5438I6OI/rUvqn5ReHR3XaUuuRGQJx8afZ4OLS/Fbm0ta/tOYL5Xd/PtFpe
JUYrNUYxLUVV3gULKwChqB+5N1SDJZrFL5ZDSlmdHIIg1TA7s8QlrEH0xODyPVLb
GMpWiwYudQrFwZxOVAph7nk9+VUSNCZGY3CP+OVqppnoURobBI6xRTUii74i7eJl
vzZZKwQGND5EY+HVqFqhutMRnNXrjfQTqefNqLPI4rK52YQPfb2967ydPcr8vpD6
hHS/sdWmAL3Wjs/DLg3Ocz8oQD57+RtiRKZdQ+K8/BqOeVQ72a84iwzluCIc2ROa
vSYxiYFURbaRYxolZmBuLl9jKi0MyXqwBljA8uGXJ5jQuEkXJD+OJGI2b3f2xva0
BzopYAsy5MeqnuAsHaRbxkJqqZqfhI9lkiAyUw35qlCwEyAw/721fbMdLvUytOvp
AMHGxDNIgaiabQ7Ti1vw3VaDW+givxS+I6Jg+0FUBatZC7c5RzJpJXBRzxIXaoFL
Pc0bFXoz0W3ctwA9gmhwoSbqO6etlNebkgXHpDsayha7wSZjK1kF7f0TijKWsmnb
QNvxsGT8Mkgk9VeHxV+jqOgPMgdeqXP1vycBa3F78Afj7Vs+Hz86YGYFKgpMHQNG
XoKNAEskoSpqzQon8VU8jaedJhCuLngtZQ04+jNCXxt1d+XygqGEE5lXop5KtGHq
LmSzG89o1IMt5p9HKR8r03aJJpHgHzpJWEvwSNeh4BFDI15vKtINC3nuzrlVCAmP
G7SerE2xiEs1lCF44scQpmMCLBvAnc+ESudczTPdGndsUU+gTz8pM/J7iUWvXOQz
PDnYwXAa3830fuy9AplX7tJUA774NsQ8NxPETvOfFdmFEIfLmVbdqHGOOhCRWbOt
ue/FpN2/ytYNlQ6CLyNx8eqQjq67StCURTTJtm4Bu768TrdfAFWHtai9cbsI8UCA
mdGXBopdRfUSyX//DRGQn9m5aEEo0AEMj5W++ikuISrldFNypYpnqI60Eufx5qrw
O128yuftL5Z7y1MpAjInkQXfhpa9J45Oa78JnLrxEVyUKPX16zvYARuo6XmSTJf0
tGVKB37mlAaOo0gKl4pHgKZnWqh1Zcrrel9IOlR+bgpYnRqOVrqxz4UJZxSXzipj
oiQ9s+45t7J1pHQNtMsodqFgYB42M1GN1dv8A9TeFxEAdQ9bbQPE1LuuurzQ4qDR
ShKTdqeBiGlsuuHKBTjXHwu6V7ddLRsbkjaqydxxDky0zTLZUq68eJseOOqpftP9
WIDZicqOywBD0yBPIj8aQuNfWkBG/Mz7/CG8W97t1sMZ9tkFeRA+REY1b/pJQca8
9Z3vvA2iUcBLF6j0MhWONroU3j3z9bBcS+J3F9wgmj9FQvleusOTn7oE9S6ipHR6
ZCf5/L/gLPdHW49G3w0pJ88GXicSVdgUisREaG5cnK6h3KILEMw649Zm7M4oDvQQ
JKjA5sBUD266wc+lTb/oKk7udoLiVcCZEzXofjN84dEsPx+n3YeeuVrU9BzCRg3O
pw5URo2m7QCc9BP9BzUCt+dh+ZsvlxtIqaVWlrpS6N+ea+g1WT9cVPKB2RHk/PQF
vMXOzibnlN4uSdNsS76BkAaciprKUPAtZrbtD7eHl13HnJCo4PubxgN3zN72WJXt
K4RDOphrpsVV0U9Vb0ujcFP/q+5styIozNOvQa+f+s6nYih6xk3jMiE9U3RuEp6d
rnbRVp4ksze7ENwgjsz40TusMRWSl03B+ycI+CY1bqmmQrAaP7U8Z7fYHb7neC9Q
hNrW9J2n8uQVW0WOxRiG48JRoEmOsG9Qwp1Hcu4ANy8ObWV5OlXejEn5Oy3CMWX0
SM/P8h2JQvIpWoyzfkFfUXlSiCX38MaOM/8kuQsv/skwb5avRqGZk5l2MSebXZtY
VdaUwbi5qXM6eXw5xbygjWd+qGberbCZWMpALHOtHvvirNoMJnltyBh4ETRw39Bi
NXoKEf8FL744XKzTAM5k3Zh6yUSIcd8qSV2KO0P5BqKVoNfWVy7tBQLc9NE7sjPd
VGxDIayvC2hjFmu6RtpR3YW+nRgTxgMcBFrX11/PIc2eYpB3gs24QgncA6pUTLpl
6dMi4UkhlAj41lN7k6ZC+4q1lyCg6+m/nWaargcgfADeEyek+zi7AXnOiuB5Epto
jBy9+wxOg8WvTaOlTly6pCTxm6Zh6CodFI5iQe+n+skGE1FFartqa488QEkgC48d
1/7ObdlhfWfqDTRnTY6Tz4wVlRXUJWT5OdK518eNlCvCtbxv21J0iTfVrw0+/tYV
Qf1DepbM3RYlZ7axJXLZLr47o7X/nwV9YdEgPDaUWSjUVn8Fed/tmdX2V7RSTrJz
jy3ceyMpECxNadVHQ5kW6tZFdIeboZUjxWV8CVsyVqxsEpm6z+wxvuzbDZg6GT6q
O70J/+zrBgtZwrN7fNDRQiC/f89WwMBKYrPP9MwlvoZROmcXOX7PAwTA4lj68RPl
rGHxmmnud5cu1MuTCooYMwpbs5cAF6wQGqozumB4Jdd9MvOI9fMJ6GubsUqWrfhZ
M+7GM8iiGxg5rN02SZn0cZPz3Z2DSclndBdSoBzLw4gaWP6C7gnTLHPR6rCL0sqk
1JA9qJLGDxZVkryzh2fURTe93fSK459x19H9diDdQUw=
`protect end_protected