`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 3312 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/9huKRhRMtvnNqb3Z+UU7TahEoHV+T8U3P3ufru7l1O
3DlgtZzb9QxCbOjthp9+wDkjygH0eUfDrEl1ovhZG62GJ7z0J5RzOJ5eFhJKp7u+
4U74vF2M6HNyofjztNM9X/M2E0togArb4UtgitmdK95eS0LZaAP1htsnDJ4zQOmG
UZNXUAqNEdWwwUQ4pOEUfxXXlF8cVpPGOXYoHDGuSXiQ4yiJlS1t09lOW24Z1win
L33rs2KlOQY/5q7iq0CD9qLYiFyg4BN1RdmNyNwsSmsWtMx4Qw21blnCqUCW8+v0
ZQFymqr9NF3g5KConYbJLJc3BmPBAMZxj/NfPRWuSXS6elGGQAx+NbNkRHAEttjj
j30i6ldjlCKt8PB5GG1n75lzRu1PdayORQTMfmNLGuCs5MA0kE7reXCvS4xlMk8T
VuJkhaPmTpL+6MM86bG7lLbheix9BphtXvm5wXLtnaxasgzojDyw0X+4zHA0G09K
eWMBiZNptlavsXCD0mIMPeqtnfBIbVRBbEE9FcSBP/6mzN9ul+bbeRFViv+cbeZC
Tn5D6l82ZiTJ2/6B/q+ds02s5WIGWiuwY2OdE28SysxXXX0rtxZTYhp09s9yVqzg
2jAxiyeThYbiaB/Zueaxc63gBgJLCggpopjWr9+PV8ly/iKTQjjO1w5m0649Ct6Z
CrHq5BhZNCKOzp0lhWsSVNpPy26QU+bc/XkM772+c8rp85MDjc6eSHelt3WsFylY
PlIXYpWIa768Zic+cUZcWtBBGhtbb/chz4YtoPGcq/srqvhpv/3LAaD+VGSSjSN+
PDFMsXs3X/WxriC0GnpMEBHPI8SX+sO6zY1QMg8T3y37Kwp1IdgT0cb4Bx2GBcZB
FX0oUa1ERUFdzhYBTGiULz1xU0fEqnWjlX5xucETjHiquB9ZPzQXFZ9uyfOz0/bE
lG15NaMTGJEAkKXH/l1vMpdDmqSIht1tXjbjYReyzij4YI5uzxaXm+DpLAwnHgGM
lQQM9TnFWN2blOBLTEfZa39fN/saIske5R5cOZrXEe80WHO12X2KDvm4jiD5FsfZ
QHcyaB+GKa4+P7UFGoAfuOx2qX3qT/o38U47RxjAuZPzrol7R7wW4Xc1Zb5nQM/b
ehVBn0Da8wlxM4BfUqLYaZX36fjx2w+HDhl7S9hFwGruHE/93xgYVjulj0CIJvHw
BDfWzXZCBeWwJT7tQCFZRiOyOemEo1JuvWBp+gb2f9vx1azL9dnIxlAoV8KdgXkt
wpEafGG7GbmtEWBe8kcoSxrsgtc8t4vaS/FcXCdF7YP6bWv8+ayDgPxpuvEP5taq
xGKBFscFg/KLUbIzQkLaQqaI8GNXnxwSNzn5+78/wPjUT0AcwN0s9CgPJdZ/zmW2
Q54DjSj/kvH8YlxtH/H8lZHZadoBtlorkBy+0Q74xmi/gxf36nZKWQV2Mlo4Jo7b
SmzcdFvPT0bM9DFG7iFanJzEDfygyXLwEvwx5a6N26xnkPeR2MnAm7trAQuaO/yu
/aCdGD5BDNCCTx/Ll7lNAtV2Bb7v7AA8BPZNFVj9fttyVEmUzCX/7XoShlwt7ov0
HyBK62gPHVAK49j7w/bGZRU1Xz8ANspE5q39+MGdCrlgfQlfhq3os7hSEbz3MoM0
xzuxvsCunedpoUMSMkbUe1RfiJIqkXK5pYcvMMCM2qzcvb7PT1f3D26/NJfakssP
k5QqngJqudRsZghjSoG+1u7u18/WOpFcfFocTUYsRtHeWeOxZr0HhMairaaR1OcT
KfbXFYQXS4VsMsi1EI3QWOzh/djJYW0NNlhd5PvgqpsZEGipFx6XJnFHlD0O0pju
0wqDRHPcW63Qmgiw8bOJn28VAV8KsQkcXBLH0THXqAhGmElZEbXELoE4AIOph47A
4SOC1p9875NeTw4KnN3H1xJrMrX6TKuD4jYMaithmJDJZfHCYuthOcwZMIrG8y3D
QCn4yzKKi61s7LOvW6BwzhH7lK3CtTBJ8bJtyWZxjkoM5HCpastBjMkSrc/OhwFo
uRtRy+05bzrZxYXjmbvnhz878mbNCUMp4UJAgSf0SA+FOMv9livx2FQ7Zcb7s7H0
8IXx/LXrcX5QGZGhVtHfOOTXLuo1VL3BJX0TOvCyuhGbQ0JFtB/TeZx10nrfDF8o
r1ROCjL0rew+37PmcvqssnPH42uaserpPTB1NOS5gIlGGiLHiqzD+rDDMf01i/ZQ
Y/9fVGe5JlHE8UZjpSNlffQnoWtucLoMyTFoUx4Pl7fOJi4eHj6E6y5MyQDiSfM9
seRQkzT9DNIRMWriVJy8YYs+eIuSPJ/PlcWkua5qmKq659f+WNCH/2SQRSaUZnhk
whO++xAmdzkFCQ9E9+lFNqkDva5QXsJ6aXUVjoROCgqLy/zsmNOOQPiMM8uOuXJ1
JriTas2OBWWhOuPFhCBBUQhE4BlJRce6QQNs+7O8czjjfYVBT8RjrhzUf63IMRbK
GoDKezW5qjeKlKw0kGkZGzasfnC8AB3Vluu8vF70udqEljvgBbHrcbfTH8DkR95u
t1j02hL/R1+Hsa6DOA40aJn/nlAOwRIu1cTBIHmGpyihT0/YugJRaZne8acjl7tX
dX5uhnj+BpO7ZW/dumgag6p3mXsrJmQT8G9/wd2bL+9XljCjDcxJZAYCsDNSr5V3
7SUncdBOUP/MCS9vq/6M/0yLqn/j9C3tQHf25/+HalqH9G2XygfOXCMgyaL0EcGb
nacXvlX15KyjC2a5KdP3SzTBwrNTBP5BvSu38oG+iREb/k+XVkUTwfy1gaBiNJzb
CgkGTo1CURTKyVOPJ4qWv7GbFRiSIrW7vfTg09l4uavuGngJ9sjJ6ieBryGrDX14
jD61HtCwqnboY7WnsPr8Sb7t/Dn5SWXDuWdYGH7ZVh2u3vuSsn/xWdkmt4ui23vr
csUd4RxSips9A2UhII75nJpEoXtw6FHjA+xIEHunbsleE+FAC/vtsT/wM56eQ1pk
M32wYQW6VVsUMIZzOnpbfaRV4yaEbQPCKHmmavLsEcG+o4yIYK/6//lQvaW27bOw
OvIDXJGTgEzrXjfPNnIJ+SRq0tiWiqPcMthV5PfS6bNehJdWb2lMYXIZMMrTlkC+
/8XpPdhMHj8TQnYBkcPEo8kUnEB35Z6y3YBPFVZ+QoEtRN7+ufJi7+TnQeRKv2mw
Fs1jCGCfQcoEMcke0WdRaTYIFzKfJs2gQ1rLOHL+AfwmQmEyFQ97Gw9QjUeJWUut
Br18IAHMjJT8GpPbS5/0z1jnt42oVLgm3ZQMQGhHn2mBNCdlm4RwUsLQ+JfIJmh7
5oCdJiyjivgD3dlIDeJyy2Q8Moe7gtWCEkwzhD3gR2IjZeHc2YIeKgj/EPRt+WIZ
M8CqkWXE1gqAfH2f5Kra2f/2XqoJEZyH1MbyEmunDRT/++aPLycvlI5t+GYukdp3
oxKvMEcV3n2jPgHAV4TeZKrKvKGJxlpICWUy7wGKYQcStAc0d/hb4SrqloBqgYE5
v8STG1MeE3Nn5lN1dGT+tqYzZjXiXskgPMKCRin3tMpAP/dgMnekLwAxqAwLi/iF
U3oF5jj1w+NteCevj/osS9s34e16aEpwHfttXo1T3wkSRZPMBqce4cve8INjevb0
WAbiaLQnWOcvl2uGJ+PEfYpki7kzCUA+i7D99Y6kEbPyyOiJXT0t98FCgUSpiw0z
LGl4llTKcL+OGuZcXQqU3E/oirZU4/MwTPcSuiM6tUtB7qzCSHWV1hcE4cJbWQd2
t5eES3cH8Teoxlfv07LSf/Zh9FvTUygvmJTa6mNfRudSynaswx9IZVTbOtjq7En3
7z/QybutMjYe16iahvvcuFf5HztGEzQWGQWB/oqsS5E6kFtge8qFSEoNyrFBK3Yl
9BkTTtidLfZe0M6YenAPlAEc4MC0TV4GWuf+JyuPvjTEl/mEJij2jNI4LWcaxJHe
Or9fik6NODOjk9ucl+0iJNreniMe2oj2bEy4lcUNdLqLTr9AMJQOAe6ZWgdlDJTl
d9kpBqHoG2hc1nWk6sVCkdqZkWFMJg9o1TDb0LEX+9I98/y+slE7wPdf4Nk8intw
h7jdE9LBCcv+94G+zUA/Go6KYI8WOdlu2HUoNCBm8FvzZPlts3E9pOCbwKiXjShm
96IYErWnsjZjZ8GmnCekNx7buv7egk/p5VyuE4n0gNfGzLnXvlDML+kyVpLKMrsC
HwZ5rajj9AHQpcEKWs3GsXzCJoKrUaE7EJ2kEhbtFTU06jqmUWD3/DF40ICixmh0
0EfwGarDa/g7AW/FkGlIhLfZ5e/TEMVEy07DYHua2zW4Q95QtvYBdnsn9VY63+1L
ZP9H9mX6BT2kDM/E2WHegRgPkB4VBi0K2kdtUDGHNsqL57FjuhmRQUhU5PuD7mvo
`protect end_protected