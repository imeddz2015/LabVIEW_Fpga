`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 6032 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/59UwEX+aE7FohaWu0/8IpTj7mav863zUNIsgIH2BWb
Abd9opeuBjbGF/waQMI2vMJTwD1ie1YueHc3nSNpEh4OXp8P5ybZFY89uyGz3ztU
W1EsuUnchJoQgbHZ/sLbgtGRgsrAFn+ZoIeGN1d6RAF2wAESJmYP8zw+p00RvjZ5
1fQ25/jflXJ8bWLKnubPwmgtk9GxoUEcmLhAVg21Uoez+hWi87ZtOEFJ5zI9BCh7
mP5i9hBoiSVIPtmwWYpJRfp/zpDwFYYmpBOlwy38jpRMz6l/4WmsKtf/QrfvFX3c
Iy7irQVUm97ShCd+u/+9wxUhIr316EW9VlGmaBO+STluOWNR8ZMma+2m7PcoB1Kv
24K3M+uweYFuLFnHHDj6kis4K0phMpKg2G6dvw5aNEDcrcBabNtcMYp9jcOVH8Xm
LZPtq2JY4z01LXLw7rzFyf14WgQfqlkWyMYn5sDwXEbngm3+n71aTbnDk2oz6vyW
NzZGqJdtkzJBLiaGm1SNgamDHu+Fj3EQiIyEE9s5SbQwLk6roxB8thPAUyi1w8G1
lUky9AEhXyksNIpKjqw7qsa4FoQTkybQ4mw4TI1nMbC7U51iUzWcViagXmlJeaEk
2QLu5OVfFHZ3+msuYjibzwi7AzEU/6thRRSLrHKdR4tTv6Zei5yGwttPxrfKPFyY
3TgiN8RtrvATSsJcoPngxeqKj6TZDzg222ENJysWJ6Zm6XjZubGiyfkrAn0Ap4CD
TSawdbqVWPtugL+njCuQWuwif2yIpmsp79mVnA6PmN37O3acEglCZCi3tvyzYS7U
2zXac+bhyI6faLZd78U+eFAmvk6NrUCYXcrwsAoVmaMy4tXZ0svrqOiRC9eOb+vv
pJbtX53/+SiMVWLQQPMYoHQ5Vy+CZpU89kERSVP+8WJHwJJv7rvTTYe6DwudDgUP
BjS0DEta+dFk5VFnvciMI0oqfkGyJMAMqgWIDvLD/VvZVIoHfH/0KojDJ/U0u7pQ
ECrw/2HcE78sJsSIpMj3H/sC2Wj+3oDtyIFpi5WKYp9LQ025Xo49MJH5W6txhyfs
hYdMyUPUwJHid2vNHqt+2Ns/F61OoV6rS9N7K+d11q28b6rqKdqeqtdmgonX9rtc
7cJA+kuY5Zi5gIZw6gb8GzQfuhW4tNunPgK7oAIFrqV4xCqfd0FGxtUZOYwS151J
Fym+TgmVhvX9TKBO+iOtWrR/3/4hkPJvA0rbiGltRCbsNWADLD1labjK8DfF91DZ
0oqG+oQR7WbrJVNaAP4kQpn1u4mGPH8FTf5k36aQW9M0++Si8XMIRHbhqJ4lDPrd
G+nCJqZ0Ey/smkSFIQSJNQliENUPwBycE5d8H74p6CrBMa4afivQHK8X/BT/57BT
+g7orvsYvqpJpQ+2uDSymoJBQ4iKdJ2UFyDMsIqVkiLcW0NokUFsWE28Ih11jVO5
Xo+VjEb6SY0ZXy/JFZ4bPDPJIYoxcO5pg56wxNOPcmt/lk7MeS7oNcoV7Tzwz0Uh
HUdUCGilg43QZq/OUa7PNJnbU7Ab0HT2amZvcwxqjaFPA3zaPtckUSFXgHFE+t3o
6PKGxMdm9DoFUmPlwjh5ZIlZ7dS3GWC4aPULrjNWNtmhChnD8TVaXDNBRajyoxlK
p8qkZsL9NWvwwU2w3vIyhF+VX640PM4Ol+Br7GduvE6g0FoJ386u62Z95Z27ps9P
D1IFoAwDbrWR89+j91hoC4I/qEh0ukn1n3GMNs8lkAuUdwGYEOyqrfwlhqJliFUM
btVnUrpgOZ+ZLaKIuTSNgq6RH6Vtjk2CR3Hvg1GaMPWB1AzR1elmRsY/RDuI7LWZ
vR5lU5nCCUaEtDH7+tKvUvaUr9Pl0TgpeM0Vw6Qbs3kpTUB/h1VlH8W71A4EZDKT
5D3tPttQvZP4SV674dDn0zltoHV6o5IeXY3YGMINzgKfQaxnyYqGhFMOgoT1q7QM
b+0qQOFGIHKXWuNSZ2CmGq7p6ofs5xEhnSMkFMFApTqWdnBju+u9q2IyL1zMNetb
uMl2e7ADcWe8pUPHF8yIFHEPcuAr1AWD/X8XARZwdq8nmZ+Cdf+Qc7Ag8CQs5MXo
RQp6pE1oacMUNm2WKX6Glsn9Eurf3vHFQfdW1I+bh2PxpwEffR/DHi8MGoVXyNbE
agL/fAfZtbMa9wV61cA2L8cpI2qyfCm0feTTYq75gmnAhWj9tS/KHkHpq4zIam3l
uhbwpcqiDWXhdxxYG0RKDSDjuFgE78Kajb1/VsIqzEnZcyKJyok7mVdEB7pdebjO
S9vWJrKK+7SrjwINiOKswcRKms+MSt0n9hJ6eyoUD8u5VKjRr8zOtz+JSMIqxxNN
9rE9pmF5Rrwmx47gmk5iNjFMC6stSlV7HZaycY3WKH1xhxVoOLhi7O5rQffbpB9D
59raX++3CsZA5CpPn7rkZe96eqzEe/0/QzGPXH1t+gb6jOjjsYCx/AW5noMALTGj
SZJt1OPvUVjddWP/WyXurYju42PMmBHvEo234c8SHbc26TruJybjf/VNWPWKbqoB
JBVNBz/IRPzOEFRYPbKOXI7K5KkxbhHSByG4PcQhcdECX7MYP+FYiR8UHuNYqV8m
d6XNMINQT/odlyv5DCDCXmBEn1/0F7wArFX2pWT301dceS+2P+dR8p7lNE5zmWGG
4OdA7ATaAFmjUvJ8oribBjXw33mm0yhTZZGDK5bR9/Z/Pb9cHDwvvtvGnnSTtzQv
lZ71pkYMiGmvd4uk/0bOqfvteGZlXZplAedw602FIGH7eoKFRrHxa2UmRx3w2mst
fNtdq3xJXkYpYv3eDJIGMhLx6vekZycsIDWHazj6W70nCHkc3YAaMNSSVsON+Exo
CROD8PvV8v1aqrXhXr2YMUwqQ3Yr0qvPRy4fjFysCCYZi67of8e/BirxKe8aW0t4
7gvna2fl1dwGOyTMBhXJJUqzHDhIZdoGZ5KUEvtkAjkc1XX9qyhLojeg3wGsxbZx
gCgKAo/kF5kRkn1vIF0jHiKZkybm7JZQu15MaqXrGQh90VwzyDNMtPvm4pk4MPDZ
EtZgIxdJiosOuK5LXUD/QojirjAk7EqC7DyRRgDXR4p4Fvo9QFeNPvHkz7O1VCQf
c7SS4ktA8LK7nlfE1jhSgrVg8r7TgnW3xhVbBH+l/YhZHR6ffkIbeGq/SkPPE3dj
RODhihgKqDAhlpKLTteBZHpETRH+pWCebFV1PjQ5gcg/zZq2yvPNUKVBAgdYYkYI
VTvsMK8SpZhG2c6c1XwPHLnOCoyRP9oKXSP1i1kjiv8vttu7Fjw+/G84EBgaS0Z3
uQi+p0oM8aj4leq+wqP5pYPzltqmwsoc1z9oMcvXpQfFuM9+xFIyraUKww2CWcFB
sx4fwcpe9dP6se2JfrM3IrndYQyzA4FCd1D9V1KRLavFqBeuWKsaP4Ew8hgS7dL3
QQJlyIRHyUb3FagO3v40cllTYwVZ45BQs5Xi1nP+OHyZfjzswzu3k1KlXDYYKhdK
QzpojIt3QTbu0879H92awvUJO8Ln4gvo2gAn1TNQK4WP0ewAemu1PL0HeKJhB/8z
yvoqRw7DERy+2tRFpcRLdRrsoWola+L3HqEsH6w8jv75NKEChn4rt9R3yGX5rkjL
5bVyEqlo+Oo1X+HNkHSnmrmOeHYp73yzgHboQ+mhz7olD4voWiUgSDq/HN5qY1yp
tVcjjt8jyJQA1QBAbbWV4CkaAmeVT9lLy7rnlWC9I6Xb0qZfslDTYlSfVjYZd+ru
aKHI7TV7HITBVVf4Z4F4tgLshqJWcxgLOKOuM5T/xBgwx+vzOXtvq6UwlhGLjgOC
1YmYTwD6EbegltE7U/m76PbnkxHRtB5k5JhYRCV3zTCl1OkxZ84ELjkHUv9T56c9
LHqXpCJXW2cDMavgM2XGrQJIpk5s9i5tV9qFbf0PltY56gEVUB69Ti4VWi4CIe+F
URwxvgoXqS6CvTM6MvNa+f6w5q9+TR3wdJPWrgXmBFgQGu32fZX39ydrAY5lYW0h
5wTcPaOj1LPCbw2pL73erW+uHHUUVV8jYvW08vbhnozFOVWbWHlGHUI5XNRmM+Px
VnjYnljmGlDJNYAS8Th7/twZrb3g5jZwINyPz01+hm9LW3tG1ydxkRUawR50fuvf
E20Fxm/uduVyXtukuLcFA2Hio5s/hNz+Dp6PFI3F2YWNWhU0+OxB1nw1g3fnWpi5
Wm773wzjubh7zWCUGegUBU4IhNSmgYPhfYZqVAP/RKtkq8r3MJg3x3iqmws7W/00
cm/CMct2rQKJnYd3l8E1hjNNKy0j+nPpP3d03/nBA+ZJzeqgpLl+Pc+VJ+ZVwN1J
FrwPllT7R+hVYbJm8E9/M2cqXrFKWAkpsLniKIM5qKpAbT0pIWV8DLXQw8PApbXp
QyaSX8Cr+u9PB6oJNlnanVXZ68/xTNgpqFgLIemd7K+CWsytfSzxvla4FKWWC6tK
ll+WXdUAjibNYvlTLeGjnrFEheK52GTWsE9jniSFPrMd3MknoFu85aZ8G2AVlbbj
9zPQyiuqvJVBnfbrhqTIK7/PmBEAcfrAiuBA7rGxavScxilgCc1i3Cm/a/5Fuev2
NX6tg04GZrwUti4yx8cHKLcnu/nCYe8TTczZCjPTDRHs+uHZmEzsQ+UwB835NEeC
wLeRlj4rOail/tlG+bz2HgLnFmppVNPTwhKZplK8cqw/nWJz4cpY0VXN9MialquX
oZYz6rvnTJ3gCNt0AJhMIwUzUNPxWw6QYYAFt/zE7GdgmNA1eYU0DIk9Ujhbp7cn
VilM7ZyYGuyjmZppeiKU7rAzknarh0bj785c0o8c1379w6uJBh/8a7QAnpC20LWI
dB/AaHzbsA2cst11+DlpwQHa0OYP128RJXB1t6qdvGdQS3ffE3sMMalMkT8JIKp/
v2wgmXUJP6CAuteubKxS+yCu7GrWJtVMYjXg7IZTMenHZgEAz9thHzpp/YnbA4wy
YjXYQh6kI/1dl1Y5ixY6FtuDL2cah3io6pzBQswl0bAOk1A7UVM1dbPpGzV1k9Dx
AONyIhW5+9gvhsifb4hgBbRA/0Jh2q59ymPm1msNi+H+W0hcyRbXWy3CuYp+91nF
xo0YPA/8U+I2wAXyvbRaCncTCEiLU2BiFPBKNFcpKGitJk4O0G1FLFN1J38H48vw
dmRqyoTcikLC6TcYwHj/8z2qumCCjrCwNpKbluG7Dmi5rjsSCzLHTydRub2d4la3
a9OStaNggr+/nsdu+cood4wwhd0xy986HG9toa3JsUHgNRq4sE28lF9Lm6vrSe6z
dmwO8fcQYewKa87tg4plW3wVqndKHpPfuvX0HbQhiozjHVMNWLBP+rduRZ0OdbCO
QzqdmUujuJ0M13CBEUxk7XILtgYE5KBcWUC81tbTWQBPlITh5iaPtVnS/su+eMon
ByIU7T/yuIbmH53Y2vXt4WZ1NPFArvhSxpwvCSnqQTcdOpAD27dFz0wXat7vVlYp
A3KlyKqf6BCdUojljlJN+H1AwQTJiEUKL6CA34vN4FXFI8ACniCBmo0HMpbAJX+K
UMEC8IpDxgCql+SCdAwE28rqKzWMgQXcD50LzqvTkR2ISCniWwZdO5yL0q5WpRhk
A9YvdNDxX4gLQv/rFKLOjG7mCTZmhAxcVYTfWBjAENhXtLJ52PIGL1hUa2O9OX3o
kO+yabAtHgcKvf0TPpJKGOycA8ZgtbAJ/otzDoUMXvTIPkUJQFDqZdszRwTYUDxN
GvVRB8/AWaVe2XBoOgqUCFwMJwMkHUmxtzMv61g819vi1uKGgbzssc/tFDeq1bU2
r0OPTQEFa0K6nFm9WqrEEDpEzkEjcpdXM9xnxC3jV3dDsj70Ab+deHUUteLSaDFx
VyWw5bbUBuGzMVdSwKM0vWBe0pkXqoQYWBzJeGucN6Awv2k/50UWDEagmnvLKSKD
UnpL/Wj1QGNMJDBIcxv5Hyb6wS6XVfc3KuLbUL45iapZpwa54zd+OhfJr2LNsyBG
rpx7FMa3KYraXE5DhRssd7zjCeCQj7BIm8b/TVdGdidqn3MipGr5D3CKTp8EeGy1
U3EYiFzXacWI5ZKGV5p5i6K6uP2nGXs2tkr7Ly/8/ECsIuyi6kPY6OtHJ89d45xH
TJd4iqAdJo0ieokxvQLYbSOLLW9fjb5PH3q7sagur7Yfgip3wDjxUQIyieGMB3XO
pe9zwri3KUhacmlXL7twQuY+RsYeX4FLAR5ddSYIqmMPpCFQ6/pupv46Dpp5rfoc
He069k/eyCZZYyZ1EbSt+JQxS4B5i962ur3+1ORulU9PrPuakEOSKgYNnw4lMs+P
fd8oYzJXigJQS88+zK5n2T7fJwGNHeEmZs83i/2Sf9X7vW375HRJpDCy0ysEc8l6
3VcvuQCRQdDi/4QqFDdm5H7qvFmHqk87LNe7ywePuGzqh23bk+8axmykBsraxIcM
jpRClxKhEwBsbDyXY0MSI810/nJPiS5+kXGql7MgWW7dY1z+tHfm8W7pFqp8BmrB
X324lIx9U6+4Llv7vTP9ZnEWMuJU3svaZAvhMN2zLeOz7AqoVVwDRbP3IY5cv48I
2NUZmAI2hUasUwn672dIryYc2KeU2ZjmH8eZPL+9/rMbLpley0hyRq0pRKnb2KpT
G99N/bVoC5NF2hj1TTgT0MtI3aJYoGWTwytYui8p246mXGe5d5ji8j+jkqObRb9P
ZkJIqfMRHjn6OfnKgHYayjUKMIU+R9y9MwGh5HW9y3zPFkxLvG0602EwwtAMUH89
PMJz9ftD3kdXZq++QcfIMVjSX9udaplVPkYHeaRpDB0bHDcBNjDbsseCyd+zpphD
VUQlYifTpZcL5x0ew18Bmk6ZgLJVhF4qndeZgcgwShNYga6Kt01xhIYeyZb/QI1m
rCRE6hy3ToY9VfFj3pUD8aymhRsQFI35J081R1DdWVKKSom7y6NQb7SYlGmPntZT
4n1Tk+peFJPRQTj0oT5twLj8TaTLmbkUZ26wztk0euqiHjoj6xEVAAiUPHc5qnVj
rtOgPmiEO0jSgeMpQkl255ZjCHyvIazdbkDXP1I5Ky+i0CkS4cGdgypS1jzojhri
sJ6N6ufmiORq392RLO3J4hVKkwVP0CoaUanytj1LU/hnhdQG2OrMKGGgU6uGcuQK
BI6UVuHITwwPMxQH8E6AxNgdXOdmhQxCcFb1YaVXHZnywXlabddKHmnPpm6zuPjF
W4NqAdWV6sE2SKV3BQOwC6yN/SIuG0jy6GrsRLnAIimA2vlG0tOoymGNxDwrTukG
8tDsudUnhSDQcEPvC3YAED4WlO+sonYwvHuSzbkuw/sMrjCHkHaWLDMdJkHJiqLZ
M4eVqibvrbuSM1OSKvJquW6FJiiLWBZco+G9U3hpG1IM0j/DbWh6qqs2sq2dsRqS
1pWsC0aAC0BybiUE68OlqZ7hYKXph+uadNsBKiTyqINYd+DUD8/wWPRe6X1bretK
RXXtCAWYBy97V5cjo5m1ey3LuTdx+rjrmEZPHK/GfF3yTGwrSIbP/3USwd0so0Og
9M+TIpodR9//G5gV8N6yrZrr+YR21pMSua3RdI45m5z633M94sepIG+hp46csXw/
kLr8HQyfKxhb8RYUnIwZ0Oj5+FVuQDgoVsbdWbeXTBZp02MPW1V2QNooTY8x2iLx
iDqPBxaT7YKSTav8vXuGaa/i4Un16CJxJZiTu5Ua0/7E6yoK4mSlgfSdCrImkrJ6
zIPRWmxx2UjIbUwS6Esyro3PYV/SlHO23DVahxFSeFvYoGqI64+9S0GD8Oo2vLIE
KTlegfjXEj1c7MZ7pMtSdB3VUk0DIUbCTFPaCYkpjOK92xOjsrRU4A7Jvt6vXWum
nfcPa718bDI1Oq6r8D1v7Rx0xeadaCa6WxpIVntmQ+2v3uAFSgJgNU4KE8x6/Evm
+k5GAvknFvvigw8Q9LRQSseMj3owqlYDRaWrDvWfUz25DBtnxVKXOqplpBW/uPQx
/6ptW4rresh1Qozi3DFE1w7uBUsypJdS8DcBtvWepLI=
`protect end_protected