`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 7872 )
`protect data_block
XAYzcToIY1VIPqVIYOouMwaXR6+iabrWSAEf0x/eFj8GuEaEd0S1cjNRhN4pe3ey
dScutQVB7r/7WEWDYSh8KlQIia3LXI2SBE8xjX/tk5LCgNzhno9H5DapHBuHJsgO
EulfYGnLpOIT24L07xg5P17sCk7kd+DRP3vcqem01wdq+TG+6eIXhe32T7uoUaqi
MHa7VDL4hKdIiFnAw7s/XmJXAsS2NGxT5i5XOiwNZNCRPgTJD2a9q3I03Lhm8jhQ
QmUKmn25gZG8jRJcPqCKqd0o1xGBaSNQos28ss/fiwX26fDtjvIQktQM0L0Hjc8Y
8FEE1/ZNyrSX4Yx2O58FGWR2kHRkKSqeiXi9Kxfq9ZMp7F1gE1iFaYHxogqvBv9X
C+owOcKweQeR4NXWjOazXHtPoSxwt6sLrFvKEm9JZnjkXfyidZygqHYKU1L5I/aX
Q/0Zih3Se5Pnh77kbkeUAWpFpHP3EmKC9p0P8dAMhJp4mxWsFymgdrX3jxS3UGg7
Nin+f1fXTleZE4UF5Kkay7maYVf/URYiUkhOHOqRXT/ZB4dq9I58QS0SxcmRKqCq
aoICNBKB+95yJAsfRF+34YktDbsDiCWN/ACxQsEJoQu62FdBEo63oEWFKkJXojmp
yBFoHRaGCZshFwfdkqoKO3bcPYFmU+gA0aR5gB1Iz2tmzVhpjyqjUs7Gdiv6zmcO
e2wwvNH9o01EA5ZVPMTk6FdIPyBSwZ89J2X3Lfeg6YLbfndES+Z1KIDkVG8foz0u
CQfELGDqEHCIyjxwuNkDeS3IqduZCEX6SeZGIOy2PD1T1wFIVzCVz5Kqd7PHrnFR
IPqj+GYrFyz1ulF7lWk4jNkA242nAuTQdJjbKgpVQCbgb4zM7hy+EQRfU4uvVjRw
xSqs+xsWGw/D5hAGa4DpkN3GZBipOJJni1SF37Lat/21iqO3eMNW0loVxJ8+72cY
31NyRsNH2TSbwtZluR4x5tqqBU9OhF7xunMexbCN0XDVCyfYTHHR1AkzE+Do0R91
MTYVs659M3y4yaGoOkV0Cz4ipasIj10jfNyMVRvnWPX82pVyf6qf5sZtDvI5Wj8Q
0PKBbiLrwDMmy5K6ACZ8GksnKwIlcaEKTEq/NyAVmqV5dOY6ZI3g7b4Fi/wSo1UD
1hSavrQ5olmR92yPOABN8Tqp7JVsXvOHZAA8Y3FySyBGCRalppipL6IxdzucG9eO
3Q5yhB5WHhSbK2lgW45oUfHWBLuk8lJPeJs+KBNpw91GDQqrP059Djv/fSq/Ov9R
Lw9DLt39sjFFCM3bhujwv69WaGyUvrSobAH52sg14aM4BzFLuAMu6KHb4rpDy7vy
Lf9Dei6PWs4FoeZZ9QXkP1/JTTRIr244W7zc/H/2K4P1TmbHi6urm4GeSihc+sjR
KpnffFC+sk96C4kcMO9KDyfx4yo2BPAeQLuCrvFBAAxGleIJHVcxGQy79xEOefcv
rA3N4TCXzkgO++d+l++KKToTqRY/fwuMB/TL5C3OUv0VDZAHwx2BlkVAqfxZxjEu
ckFnklYlsvJcsJZ6fQ/yZhD7ZS7R5RPEv3Vs6gbgWnbVYRyt7kDJ0JrBsi4Ll7Zp
KQCjEDLUPahInE5+3Jkul1tpbxwLiEj0vpZPMWEmYQlR/491FwaV5oyS06Aa33ay
2gLcjSfaV00KPSSGWY/IJfQG2VxlkJV06V0i3iurIWtU9eDiQe28hoXogGOhucIS
Um5c73AFVH/dv3DagmoW8HEL7lr350PHb0BVVfUnCibMiHqn5JAwRbhPyGBsYAQY
1G+/G8RTC74Cb4IDO+8UrjHQxk523VgV1Q9tiRuBFwz6K9aTtxt8umfoO+LR4TV+
tWO3BqzOtNUKSZdjU0BuseluohciV9n8hF2O5SJB8laOuOvX81sRlMRQXF5iL6A9
pCbeOrV4gP/RA5ipBOCnaJCHrhQEGDXKZPaRtSyu6WACEnJV/10grTWSoqWsuL8D
leqN9oiYB/FGsLO7/A2rX9AXvGtdH6BVV4nnnGEYxcywMFlGdPHsbM/hV4nRw0fQ
sJunskkJAyTYcIF7h2Jwxr6a7SuLaBnM0Yzu0vs+pKS6/NRDNTBaCWdeulQX1B8t
/Hz5ZYSExplzHGm37soJ3echfTj1IKN8gO8h2/YaP12uoSOD6bNBOujXwmWZwTDX
Y+MWSu38KznpbOuuVHBp5HPopPPZB7phmWtiuy6jJdSC8YjD16ALEs/SWO0CkJu4
5M88fEoZCYkq7ciab/kUnnjB6ZbQYl4ll5JJF6vovZ2TqdPOaG3TBwpFukZgiY/U
NqurDRRuIP4hC/rYlIatfKUhjegJRtD2NJzlfEhgW/GubZx8xQAVMUZXfJxmd2Ex
xc432t4zoiJkg+xqcmiODhEv3S0xDRukWqDInGm9f7UWFLV4ZNwgRMTA3FvXQ+7x
UW2ojAfDKXlO2NDKwjqUS3B4iP4SZc3HrtlWw7gtaYqUVyZTzPpVlp4RCHSfcM+O
2it0eyRAMSULrLwJas2qR9onIRr7pIH/g6P9VJeMQ7wJR2lIjCdBnF6VFXMlQpON
+La2eSHmy6tXdf9lngilozMt4/ym/PlTbzyYSOy7SBN+O8qTVnnW2OvSA3+3n7H5
BgsPAh+OorcKULRIDmPPARXB33U3ogj0A+Ua0kBImbowuV264oRrkyQxDMbCIUry
KlOmQkNu57b3+GcwZCG7vZkDlBy0qLqaaiKXGZ3FgcuqFCg0/jLfksrzrd+Joz42
zuR4fDA2s7yCsm0ndMAxyBaKL5jNJ0HU0jRMcdOuGgp0PcmAU3uzYZL0rO0dWKZG
g+HGJvXDygaCko+Ok6DZZdiKcduOYquJWzuLfS+5yiJlT2YC3yNE4Rs1066knVB+
78uEdsw4BwYoqPNIlKR4f4NqPUBllVCpaa+tjKfamkFm2RMY5a2cT+CFmS1t8oN8
JecCLRlD38WNU0yxSlDdI8+pJcoU6fQpEHc5Y7U7Fi0wtmcHfRaoID6gksGhZiCw
GTLCvD6TkAjof0ggz4XyyfaChszuH2LyfiYZEPX69zDOFjICknJ9SWQEYDb3yKOM
SkTP8jgAucng7igAfmERrXGQ48YsrjBOiTdkPwm+caWwQuBf0CrQKp4u9SF3nvap
pnzZkF1QBxpc4LOZV6okIzdZpXwNOQUMeTh7Yb0FC1P/8v7hsYgEjz9Whb5LsqHc
csCAEFWnNEOA7j/pUYjjq4yjwy26/VO2WJvj93UGTOq9mrA4YPoCssIXcCZkFJfV
k/k118s2UxlPDg7ddPB54S7tbCINEcw9BDNWyzYk2LXfEPshzyG/HkHVPCvob3g+
pJyLCxVnPYnjAqqnz86yFboMENWc6WIHdRTKFkC3iJ/1qG566U3x8tJHLOzW7h5J
7+mZfJEzoNqVH/bA+PxBThskiinQ8ynrz7aZFZG5h8vRzfrQIKHCEEu9cPq13EVY
I0Y/B7FaONjcrKDlX8jnEcxCxk+n0lL5NAW3hUc7LoVipJ4V7ih7X4LXCZCo2CPz
2YC44YkiX+/tKBYPld+bUD9WkE7Kh4f0gdaIFbaBUzqwItCE7fs9G2LZkYA5wgsx
52uyi1a6fdXSxlvWgYl3A2GVx9FmNs6I7SKkqfw4CwrPGLR7aL2eOTHTPp9zppqS
0lIRkZhwPoA7zsCRzEAbzey7cIzG10NsHPLYBhCfVRNJQ/GUTdir1rB9J6Naq9Un
Ew7lBX4WoGcUqg0jR2HriV1TbzdpqajMsRm6rpUnjzNfEFRN8BZsBb+PXzKMqXn7
94VTBImsYw7gQzgzTVBNFJsgBd+516Q9rLo9c2FGTgJDRYN7FwYKxjlOQjfHT8zD
g0ihqkt5RQbfi4JUO5kPRoUZhIKmB+60US8FLzruNhqT2uyFf7KVJWNfQt5RHNI9
U4KADHyKJyiyI4OfFXNNezfosLUUYYkiEu7EOm5F68xaxG7jbEZlgafaEHXbnm3J
049cgHALsbZzJFRhK203wcvx23OHNLEx08vt0BEVLEc4UoUS+xKnHTVZ0mPjq6uH
cBRsg/AY01EPTrpFUtEp86/1xubmzVzIsP1Q3vVirPFfDuxHGpq3hh0VvIjYspsQ
oTO0tMapx8xfpBe1mDtCUlB/lFbGSWgSxzmfI46jZAhrS6d45jYgprgwfUjwgL4R
kddCOROnyg68D1LaN1HMe9mHg/oAhP8t72V2HPW/Umznu7j/Sp9HDJaTTR7aQYtm
VZFcJJhxsvUOKjL9fqmAXryv33xx9F8S7qRmWVmAcA0U8iQ1ZAcguG0tAmJ1F+E5
f9NTcUX8qu1Q3x3a1DYh5X1E8i71GO6URApRlKaR3jetWzhWnWwa5jFlx4JJpKpq
oUy4d8/XBe52Ekg8fV8xOJoFHxw2OklErMBZoKe96M3v5tGdLsVtHZJHNXdSZX1H
nk0Wi0rgSxokOMH3PboUjcmhuxdtPAHxCxyFG0g48swF+V5AguQ9yTjirUnGsNl3
nimEfFFFNsizzc74MKRDk3HmC8WYyhnYBH6kodwQLd8xWjpL/yCxYBvrsYZrEQmp
KpMWIRn4LrGgwZwmCqokcsRLr9w8ICPYnxafMV/wvoYEGYtJtAqCPj7fdRy3fUYG
bOkt7ISufmCOfh20UEqa3SYozKBC0lZF4oLGTFI/WcSad338/PVZyT1nAhQEhvSz
mw1U1dRvBxTessRi0xKY9odrOgPUF3/PiW3N5m2EtkFp7RhK8ru/LfpfwZOPSX+C
FjQ2DIrpD7FrOr+6FrIiwr+xJA79oeYYZZ+riDkvWTN/C+j1Hh3wL2PdAR4RHw26
N9tCppmZ8Fl6jMkRj8XMVYqqkv3WsXmzGuUfm2JI4DNACh9WORYXfim7GpTLfbaJ
qSyTwK9ODYM1KaeyFoWauml5oj8uvqlkkUT3huxx9OIS28WjsEjSa/RTWi1zMS1H
fSl1DkpDq2X7PKc0ldTkQ+90TRFFPEBpRjkuVoAzJgPEZx3swKF6Zb08IZ3IcO+w
CrkgRFqA4TipMQ/oR99Y0s2UrgCeVqCYZA10MrHjxyCgw+IMycv6v4/cDJjIhgvn
fQJsDcKwQK/2en3icvB9YXCOYpX8NgymBuQCAmMWR+BY2qCSEpVMSmFoUKdcReH0
EC2OcqPxYOmiJxwESzLqPF0G7m+ps8f9YpcUCJ85nBzxEcQCMV2ZIeu9R88pedwh
d781cYefne7usTWBvcdJZRpttarqaEAKZlEr5DnZETVms81naUdTEcFIxr7wxFSS
BxrHYt5geytxPvzlTJDHjvyB4x+83ZWPY1jgmacqW3cGJrr6BbvRn1t2jno8By4K
9sdeTMzQZzrfOOZqIDfcqphXCTAPFMoBIYrHBHOiwbBTfg8dmRRxGquFM9wU5VOw
QTBagfmtlQlJF72MKniTWB0yGGmx55rk1X6yQggTYUjIcC1QViL69tpvDuQpaWxP
DjsqxkWl1j7ZNgVKZSDsnw8KM8npyYmzqAUQO9D3laTuJHdpr+03qXmhFVmbXBO5
lu76sOG4WW2e2OA3q6EGX+c+So1jUfroY4+Uxc6O6wl025OLxERjYtHadrbkkn0H
TaCLDJ7st90LrhTJ26DDJNL0OjUilwnF4bns01J46jFQmfFmwGEHhhN4W3mK3clF
9d5+RCzggRf7R0xA14R4QATCaPDtueqdpxHyq6vzCcBNLgNbW9Q3jvR1zhDyNZpz
ZFxwrTHmPzN9RWAtWH25SZDtm03PvoiAseJ6X8Ah3CocyxFdvliPID/kzk4Ds3iJ
cwY2HzNRNQOl3kcAfmVXAUDxiUML7pE6X9McK/1vTGag1uxuxAJ9kXKMOCipTk/W
0amdUGd13/CKalDvR5DujH4g/386SG1z6GWiAYUtu6FxvQbX5x50WqZNZ7zGKHCg
tMvLsGnUcooXQbhyxp/C7CGnLYrKuF/KLwcfvYue3A1sZKt8ZO3ecYz1tv18oVxi
I9t1tcf+MzIfkz9jn4wvOYAxUW7Q/SsT/nFnSAFToLXaxWTDAzx4enl9j0IawRZ/
6CJ954yalF70XHVI7coSJlQ/9JQpDq9is+7v5/EU6OmHCa2rwNH7ke+mecfK7WCs
x0k5Kax0LtWGrEHRuKK8/tZHkh2jWRvxWR1a+B8g+83azUloFwQJAk8YHnzP4UQ5
RKMMrpxdfkdfoGte1kPtOiQVjbfyBswrBczon3tEsbH+e6HmHini6fQ92rC3ZuE3
bb87e9QfZAZJPgJiGkvQ+ykXgKFBD+kOGI1FMUnCSWa5ClD3TlZtVmeMmcZ/jPMP
Q8Fynyxa9nCE5ax7X61BBXztPrIwSxdSGUMX/Aeb1O790KnpmSABKKLjANsi13uh
YqpFwnHS++sj/WuK+PRqaz9+0PG13z9P1mZBWzCkkeWM3+M9aVAKXuYOAZdILm+q
PGCakkB1wkYI2jXn2CblCpkRGeL1Q91geUodAJM3QlujGjcsA86EGq6PIg+GeNA1
ui/kiT2mzVytiiSI4UYFIZkktC+DS8PcyMwwvljxk+N9v+O2kgHD2amjGoMwOZLU
gOfLrPHp9gp746owuXpk3/nw+P2VAaZ1TUHlZUE0YwXvMiXXxFNiLsyZsEOKMkLL
0bNI4cSl8LIjV4sQ9hEWnRbNLv51rZ9ulTnX6e9vePqsCywBfEAOjL6tJA1kifzW
9ZE0HBPSPndLqa5By8gzSDgCun+tzs1gBWK3nTQv4CBH9uYJpsTEvxGSk3fv93D3
531u8Lfj9GGr99cNNeDtARlArNh9kmM7dzmXE50InGv6WSCkXGTSufVPkmM2GRci
R7sxJ3Ty+DHopG+YJE60ADLjiEZyHkkn7gE03XeL1K1KSzEQOunn06msrF4O/er2
cjWVXwwkEJX8qQ/oLK4gsN+W2Zc/F6fwTQ3G2lcmICtTIO83ZaGU6uaQrppO2I51
dXQCApBH6rBsnT/ny0hH9AmOernCppcWYV8Au1k8/Fed7jsUYeFrWnuGzuU9fGRD
zviRr0BIfrvEsWhroZYrbV5xQEEEw+HiBTxePKvcNk1Wfu2so6G5G2d7G6EZrvbM
ER5kWG9dhxWSqNldMzq4K5IdVleIr89tlPmbkZthoLhkJ4cBFu32SlMV4qmg/SgV
yoFrxC7DDEYLnqhwjvdWoHzYtxoMQ+sJuGTldCmQsJO00nOAwdw7pe6IxviG33qN
sygL5xUDqD/Ah1uZpGBb5ruXImTcRbJIayGEv+OB3hsOvmUpru4aquPPsxUATxtE
XymXwtXOtovtlvAGoHOf6gGGVZjeSVu5wkcHUDDzFpvVZ4EXbIpVFH7XH02/FOGW
LLlioIuqS1Uw6lKbUCv+GlipaYOteWf116kz6TuCrxbps/DZMLoHcNfZBUlXhbR3
g6KVGDCREgK8zw7gAV6Fr4HToVIJusNRLUeS42bIX3QrjeoiOIrRuBmD7AKfNa3y
aLAf/wMLQGusBQfHC7Uy4bz2baWUFOttHryH3m8tLGpal4jMgikDN2PUw9OF7V9p
FShaP1msGfnKNkX4DhvoK5bd/LwpR3cQFMv/IQDrKep2wkRc70oa+F1mbCfAXwNI
6f1bvMkMBttsXQY8k4897XyRGUG+exd6TNdAnwoNeXBicXwlFVRgnTyWIO0K6PqK
2ywUTMQHmg0UtUiMj/sE0kqaqxbVJOtyowbKEGbyx0d00HMPvGzJfFplEarIxmmZ
pUdcpAstWEShwNJQLazZVltS7tDpl9hiuDVhYFPE5QPPdD1HKboz+XouhEdQX5In
nBPsfOLQBV7CyuOFDFBV3XN1tyxICuPaE600l+jixwj/WkV3nRYENAbpFiv5LiQ/
xkDMVxDt02GiiEUxV5SpRVeXF2Pfy2ccrzCkDxVgkkuUBHvjPQIR4NE+dvGFb4aC
ljnXMUKvpp9lbC0Wn7M59JD+UV0znX0wKuo2oEv9ZFmDQewHVzeanr1sEvXjXou4
4CJuLLLopSc2oQNZY3Ehds4XvWJI1lzGQbKDoZGlyyjyUGMxyz6uC4Qadro05Rdx
dfhEe1jAKjVDofeRRrleeA9vsLIPpiQPE3HjIp5zxN2sRgiTC3CXoD/2MexLjkUV
qDNb1npHLYzCyKS5jdfGEkO+XF9znQm6vnqw8+sfeHq6vJVqWzlSeQPo7vAXaAeK
YDXfjASYGNsMTH475alEyoXF7Q+NxGzV/ttH0JoqplEkr3y3wU2/Ek/dqyKiC/34
/BEdWNL/U41Owi/WN5cgO8OHMS2xXbCeOM+Nr2ifLsvOmEUlidXNEfw6P4dtK/LB
XAi6Tfdw4qvUHCOWV3J4SWIL7F7B4Y/T0xAnE/JrpQpXAJvs0DGYLVekMmB7w8uu
z0qmojlP1VFlXqIVCOJeUJAJZEjT06ITqgYQJKP5ccoOaLfu+/0O+9T4igY3po0U
/akFTA+JUOlaNpp7Nhb0GaxJj+gfEDbL024EVxqQ/M0wadaMErfg5DJG7WqWDqO5
75jWFioTgPBpx5dZrrhetMCFq0mDBE3yYzLo4y7Xkt5c1yBRE+3GG3fO11ZzXEKJ
Ofdif09ve+jLV0gN0M0hDGO3sGraM0wKIjjqCQWWORjDeAU/aO6CZvvcCEEWLGJw
ey02vqqo4r8mkUw5lLrzylkKw4P9NoMICCR2pUXT1ZOofh7NzcZ+iYIDyWvjSV24
qt3uXJAH2jrJarMgZfbL0vV9X6LYPeRqRqVjKGsUuF2J4bePi9DvtR5H9O/jBYpk
SHzcLRDdhdDxpbsmsBl6wt2oYluQXlwtnVjnSK97vEDsaYBYmuwC4LALJ7BemBkz
SDS6ZHYFrkbJ5dluQum1ELJN9PRiraD5zaAeC6Ie+lYN5kid+X0ohUDjD9PxBRLx
k+dJwEhzTvcB+FkqGTgSWj94vS/D1wkCXoKX2peLzLNG+F6mzHUGaPcF/q34/cog
z0vyC/3H/NoLjlnlgYrGLQstrwG6Bx9HJzVwLngUe2UtUElGxjT5qrPbMG/vlg1s
bhddaFexllOcMaaZ/vXOjNhbnqIMRLNsBqOYbUyAY9kQRUPWtQiqs1hd41/B0HzE
7wYAVfXOlpXcSRhzdJe3E/28d7aTsSqs4exzNAg9SBRl0q0qHrdiicCPZIc9X0t9
WX/Ogb3Xl4SQX54V0GdQYNhMa9jR6zdojhWHFu5N7GWBkiEYPfjRQhYojq93oy+v
08VHbF73Gl2WwsQ7p1BCbxLwE3ZuMHxQGuxXsXiHEXH1FtcSM2xrEswB9SFTIGdf
Xi+TiFwaX48IgjLsNAWNtMB0jGAZpVkFXa3wTW1j2ZXzXtgcJM5Sfr0BChlTSuVC
87ciAyFKnpwYVOK6OyYriKZCzwtvXIp35NSyzbsgN6j74sV0FFafI2/DDs9zClQu
6nCA+z8EnLtCHFRrmFLvweetrRVtr6RokmiQudrKoFlYvMNBovzYIRq8CI99Cl7N
VeR8DVdxpmdwaMwi3/b4XEobcKguQKEU6ZAdonlNHo7AIrICH0WcaFAdnfbI1QjA
oLzLavolYMqAyneszVOjXkwA7uYQUipJNw6JbXn8p5V3ZEnW/tfqqh1zdGO3oWNe
2X+JrSlfieuQmW7D7eD+yqQDSWoUeeSCEEReCRUj0iq27HHwAD/NqvbBJ+U059ca
RrOUEp1psWZwpSn48p0/h3ogh91m3INee78t4Ujekuhfmq4xElXIdMU9A6KqHmBD
3RHzydtz++CwCOy15GCtY1rNLK0AAIWkGgPYQX9mFw5wCJLBo2TQyeEtElstB7nr
dE7959+QRCirCQNmB3UQaDCRhxPo5pS+GUQU+V/J4kI4V4b5JlYbyEE8XYlq/rdZ
YCmQCK6LNQRsG9YL4Q5Du60FD4s2ccKTI+b0qmsSCJnJ/OTS1UbutrEwQAxzAZ20
vJHyHA3D+40ZJcwokSGLRAaioD6i0mWw8OzCPJ6dryvmgSLxyN/mgLHudM09CjZg
/+8dtt7lquqDjI3hI0ZNH4Rdy9G0IpN/tfHVru2qd1euyGPOawcRP44SdwxBSS4V
Hh8OzZmTLcirOzPStwGIGWYNyrwqhMUPCqiFAKLGobpKosSFQHXeI3/Umg3NANqx
Ty7U2tkg9ePfxv7SIcY9/KHMn9BeY6M+VXE834KlXmg/Ute51HRfV03JUQqVcAzl
GJUPNEPMFhb4J6wwkB5Dgw3y1f884kcG9Z8wgFZjKu54O+cP4N4qEupX8fg8Vcs8
1ZROu3Iod2T5y93AO/gFnbHLqjEH3rP9Ft2MJLDF/UqlEU9dFD2vKUlVJnj7Hte7
+omp1BDnK5xrRLIHGK8QUEzRYmYFsfxdH8aY7O+2TgUoi5H+dxYeaLJ6+dnWgATi
hdjngc0Xcd6SjSOdRhSL3GaUf5qSP3gYDzb/wiJENDXGTtzNSMHny/Gzm52pImfP
9JkzyGgH5M/Qrf8EcEoM5yz/PF/5sKKIJzdAKaJhgMkDDBJkOBFlZK17smjYrldR
Yjy2PZEmjBDXYxFMHQp5P96qngQ8Wtxxtm1tFbhznNmCbUYqbEL58JPcFJw5RJjd
`protect end_protected