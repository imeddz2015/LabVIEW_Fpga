`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 37200 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/59UwEX+aE7FohaWu0/8IpTj7mav863zUNIsgIH2BWb
Abd9opeuBjbGF/waQMI2vMJTwD1ie1YueHc3nSNpEh4OXp8P5ybZFY89uyGz3ztU
W1EsuUnchJoQgbHZ/sLbgtGRgsrAFn+ZoIeGN1d6RAF2wAESJmYP8zw+p00RvjZ5
pBGEHX7wooDexzkaqKS5GzCvjiSxjKRojnbnJu15vN546bddK7AdAB2gd/pnJv4N
tQtMDjUDWOQV0xntXTZeqBrEZ1TYb0qnjDlgDTQHcAdnpeikBkwhkALZkn1GJclR
t1Itz9/NrpjKj8DYt9VyWr8HEIxJzayyENHEyJiZ+J9p7UMYlyCcza7UdERc+nQM
e761uWgNFEKYEHrRfdwqptnjfNxdD5vJgKcVImbggW5x07BDfTODA2kVckDqNp6a
Np4pwETXTTMSnK+9e8vXBenkg9ALGR7Gqg2IarNNuKU8ZdqAO1iotJHyu4MzmqSp
zpyR3ER0URyqg3HojKkuksQoy6KukpOiBDiCUvn2MKSC11dkU7+BWXfb4Ua11wsh
Rw8hnkc+xtyS269518r8T36OJUXKjNYJOjVLd+P2e91NuVlZrEZsSGG+Wh9CkxYW
85DKsFifkjW92w1HbtEmjN9hHQP9vfSrw7BiVMyvhojnToXv6OVa5SQeu5lyO5SM
uliHdKryspqyhdUEHtAK72G+oYu1vslx9qfSaltjsXjUXdHYXeBeFDbvpDuw+xkF
g8kL3Ti6dmCSYrrayqSGRhseHvga+Y0bwPRJeRXRBQMdgJWdyyi++jc4Jc+xxVVy
/DVJJ/RG0X3D3ZN207YlrwxFwFHTPGAPyIyM2XMBFa9cSStW2SG80VP30ZFyiXGd
BzNhVIV78ssJ87hWhtcjLmTa8kcDvNwZEd+IItebadsy8MrkR8pvyB9dsJOLR9c3
cBJrvmQ8E/sgCoWArUmrSLm/Pz0MOI9iNM6va/l3Spk2VAZOOvLrUyLUdwZ8l6Kb
YrPc4Zp5cKkOaXSEv/KtxvARtWCsq9w3RK6bqtylZ+qS2+KuVU1UoLLAAkM3/kHH
acbdw63Pp+MeZNDTQZreG9iSamrsKpu/LdkugBaE4GULOR25aYFgWSd62uazuXQF
yRxONj/XuJTEsbFFojeASirFU7bGVsqJbLrB67gZN/YdBhg8Yndr6Z68sqd4uRIs
z1X3xksumRW5Kb7DONLtHcGl93mywXmX/wXW1n0f4o/znIIOsBNRfCouNW1lIUJI
6oU9mRxjrKDsd9WEIeiJF5mnaDeeD8cM/8lB3FR+mLnS35Vgz8eddL+oICM6VAbu
eLOERdBGBQSkcfdn3VrhO+1JUiGkRRoO1wrfqGnzJS99vkIt/Xzk7c9Cy/+FZtwq
y1ZaT9tuaWMEk90S5w2EeGIxsjP17hgYqvsXN19fUl8BjEpYDsAa33FvroxOSrJn
zMoGyG0lZ/U8EJy1r0h/G+BbhrZP1Y0wWUomvvdUgHFI9rz5HF56+rSsyk9XIAg0
bIXxYiplm5exFYa0GSnUZr11r0MwY2Uit7GFmSfM1rHDyQmUxYCrmQtiVOpUps1P
kgfHrcUlhgTZ+YYurGZtdmWxB96zWQ9K05w27oW5tg9SVbqlRY2Xi3H0KaBJo52U
9D5jWy7gKrPObmyzz/IuKtiTR3wK21w67s3XPlfAWvveBc2nTrHkX3IA46xUs4JW
C9sFvOzf2G/agts3bVsM/EQRQ14nVJrB+Jmt46Gbj+ssBbBXDni2aL8btRt+on3L
/zMJu7RwXST4S54hWQ/hwdPPAwlbZPTLxo9xtL1xlPKmSujcpgycvfyLD3WAxqZH
qBl8VWZ2eRu8hJCcMvMthygsGMlNF2KGm8nUUdKdtPrjExDk1GagkxClSngtZaz0
N2USienChul5Gx6l41GrmrWaLf6xxv/vKFvPNI7WaqTbCoLNuMQau4DuX0I692I9
oNd+zpeDdkfIv1P8VpVmHItYZAAr5Crub0yzZ8102VoTEksD5z94OEUPTAh86Ren
0DxEnCqE2/X873RPimPoEsxsaFaAzpVeIOZbsws3v4b7Eqs6My7aYLJKqr0a+io8
eo3J3vstkHsRQI2+rDyUWZEGNbeI+xlNjatqz7hcqmHUkuoEnbLWVy67dNzOGT6w
BEMnfsUCBJGWkci02GgnaJg4bd6OGjdqfThm+mKlvai/f18Ws652tzYXJHYiiD+6
PVbtGKMSkj6T2BCQDxjapNP+z1BXBx7z306KhZxlOf3jnyhmvGxoOHIxeatFeerh
Jh9yxhDkbWqT4p0MDWhh3tC0g4ras4zysVv7aDDzrScb1hRj938JQai0YfsFzCAe
koptwJUxTPT88JZIEEVhHR3x6U7jW6HDK2eVQdKdMdVKxDyOatj7WrCH5941C4+e
LNBtvtFRKb/NSWGgxiMPZQHPZU2/icfszydl5VuNAWnhEyQ418aBD80mn8q9OXPZ
WwbV1AI18IzdxiMimx37GFe/rvtYsNf/vdjohx47TYgPWY3Sq6dbC8cUkBY2ZgEv
a5qYbOw4dTOv9Mi8jeBy8TrwN590hANPcPGUqShri2vCdfXEOd1TNizakU3bJ3nc
5vzF4xLfB0bAKPWYtyB3FOaavBZehPB6GITa7b6VUHZ3DVqSbewWBWGHeQq2O7Fa
7rdeAfaZ3SBNyxPUYubTjrXrUguutD63rauRQnw25qPYGycVAIKK/uVAfpoGWM0s
M2B5210QmWXPSfShj0dy9CTQWnbaWxzfW/pnsnbbNfTCxHwPjiZeU8z08NbCGApE
o2t51OMSDOrtWyItZUoMAsg/x+7Cu8dE22wWcYq1JHor+qEE2w1xtQv0AnjJ2Z1k
e0mSPTP8hJVBUED8F9UxZSE6z80YmbFPfUiAfPcUUT67SkqfidDZ2F4j5627AvZt
Syc3rSS/9XZ9oRSnHAmSeD/T14N5bLe+AsIXxrpLbnUWCV0vTbWFSEZwFj+1mi3Q
KnFn67jNH2RSmQQfB1/ycJH9Y4qY0WMWjbC1GCTP58jzbV/T/ruXBkC+/i+e5NhC
gTGwTlBRZTVEPslzk0k+WbGRG9HzzvHwiLRutdg6Y8ekXGlrncEEyWNP2X+7AuxH
ja+xfep9oUdNO2FJu4y3LWI86f5ZN9rvlvbQmKGmmuFVRZ2wcG5gQjrQIzsz9mQH
HYjbCaMHRR8p+N5SDOUIkgIX0oQY9mNXMY4ZH4R+ETAmlX9oyBDanUuykyE6+GYc
E4jier8qUCXDYNia5L5QT/xh79xQJlHR6Be3f1/CxkAqmTvGU99HfF8mHISM7xKE
o6GXXyj71+f+7/6w0y/0wOSrRhoBFRFYXReU2xWoGiQ4McTPKYz34tDdL8TWq27Y
6dXnC4gu5O4ziIUnF5ZV5qF9xlEyrULibmfpZXf1UInH3a9KkJ8M9QgPKqtW7e4W
Ur6X1oEuvCQC1HaES1ZcBukZlqMQHEx88bd+TSAgpqCdbkBFsyiIJ8BvHBvDSmkj
pBsK9Lt9aWs9rPWfdzSeL1yeGIewdhlxTkoO/8zATanyaTOSJHZSg7tLpv8UcLJP
RyyVRxSOmIza3pye7hlePw0thWqbffzG7GjaY47oQbhSOoiW+oHufa9yjwifQePE
bjacC7QmSx5O8zRHh6oZ6MuL1qB9XSBrp9UQ6NPLm+LwnsrYGceQMAVDCxzdl55f
ux6kAV2uVMlcexBktCxj7LaQfqHoilOZtDhaLy7b/CV89i4JnqIG+unKuEQiqcNT
I0+UXeaXhq2MdIEV+oYVpVahmZOdkkrczmW5ShOVW+8o+soCo8pYUZzV1kYaI5wr
J19fSJ1opep2tw3kJeyMxfYktoP7GVC+FdRM2NZob4wtgX4mSptPpN1U+0UKwo2P
/GtpuFa4xwGk54yTUsLTb+qLNjQP/BsyCBTdDM2pbc2mo4iKCPNDOzw77wynes82
WXUHwUPYR9zMJpSm9hTjLuhwsy1qTlAXA9lLN7tyctkKa6AYA9Nfa8Y0xixM9a1b
5tzFoaony9V34MKOmjaHWEOjbTHEUYwmKGCtdKfAL+X7XggTy6oCUd1DOl6R7S3y
6TF3Ml0pQYC4Ea3GGHnoUOmomoqAW3EE8Gwk7ZhEUGAfRdlKPAtqyP126Ln6IxSn
7FSXAXiHmcumwGkgQs7QPkHimamCWThaAWPfa0zXQYJRyCqd4eu4DseI1C3C/4PM
BfTpFfYjMNJ9/uoCb45NvHtYiGVGd9H1toIPCkXwedrT15NtTrBe01roLJqSzvEW
kCyt/hQzO/qC+GWZFGlQ9cfFsxR/+IiQhDrwm2C5kwfygJtSDv+rzBlH43bBzQbR
owrm/cVFixSU+1aBHATYRb/PU8i57lI41N1sDZZF5QrJ9WNnXXMmAxMz7h2c4A2R
LBwKdghr9cV8jt9ulLt1MBK14Be3tsmWwQfAk6Cpf+jq3UNn1hZjVjHCCAibiyUl
D0ljBw6EFnfeBtx2tFkHkv33syWw4VN8eG6H7bGnUz4fR/MiOzcCog1+rcs2vMzc
Fh1lu2Ks3qgjUbBr9uz2y92Bb3YiBnUw9y01DzuI8ait2op96Ndx/s3GpmyVA8Ht
yD7/BR/+5p1Iab3toWv4DLcrduFdZgjrMt3k/kp9+PePFqDv3bniT9hShzX+uAOb
WUQvJY4n0NeTpeG/mEV8qLAsxapuo9CgsPjE7O9Sz3r0DdfntOFdHenfYg27Zn3C
kwKGM+lERtwgJyGSyDQSXLur64doAiwZurwKIMoLCClOcTfHKze3aFibjMZe+wXh
2BqJsIqgwLe7t/9FeXHiETDyiki4ssNsh1CMWvn5Xj1nE5Q9b/99xpjIoUf6VTZx
of4JX15MQ7oyCQV++guuD6s2shOikwBGzMatPuM7/WuZjaNU9KXLkPxq0Qtf2etG
ueFZXBRciiAIigZK4xFPviMPMKYrSooUPHYfBfx+Vy7E1HledkOJOK6zvinEdnLf
LL9XLIMn0mVosh5RVJkkmgNQAb0IB7cC/LWstt+U0b7IqJF4tcXQ9+OaMN7IQ4VO
iB2d/KTaFcQBX5Fol35udH+L2q4QT4IhhoZoNxgJZUAjvbpHq4f5QaZOlxAsdOiY
tsg/7DiiBSmeUN9jMtsjBOjCx9Sop7/szaZaTJMs1ylODJF8O9nFunR54koCV3Wp
DB3BxC0KpfAZ5CdC7V9sILH9Iboc14B0W7YRFvwklK3MIVZZZVa21sbT6G7L3o0S
xzMAaRqKt0g+vNuT4+2z7WHAXZNOVbKTxtmkeeRIlhrI/tgciRNDDRF7PN6Yl+5e
e4JzzjxQLxnaZmHJW2WZ2NfofOLBQ9vo5FEYAGNEdBA16huX6N21ScndDgp/RdGe
IbBMiwSRM2z9qsCICrRW4yipSfaiz0sqAlEukAd82ZZyk1S9lc9tb4amOo0aTwxE
u5TSK3ONdVtiswTt2hgP+T9kB8zrHwwsBXEh7iszkiEtmdszB3HwMQ5flUpnKCZX
gde4n6dTSR7Mxs4y3DaGjgYl76khi5VDSHk12eDVf3Mx4NzZr/XYsB3+VmOcGZXn
fzBBl2HPgjQ5Pyv4tAVnhCpnHaYFbJmLNe9VtEsvtZtVUOMNlL+0kTXwUEaVnzQg
VUonCOj5Kf09t7uhAph8n4cszB9e54DCuu0OwKtryA1DAbFoTS2MUgZj3jSfktiI
Kxvl1NZMndmRdwqwDuPYk89c2v/17i1CJu69gPEmiL3W0kZbfso/759oI95mC0xT
W2fXrptQIuzprlgLuTYuYiV2n7n/F49ET3JaEQkFEU/owWwWvNCl8oRbnZsNDJGs
0mT46jsb4nSc9LmW1bt9VcTpT4nZXdNhg/3Uk7LEycakUxsUcgL0LhKGM/3j9nkn
s1pTbb3F1OAWM6ym9gxQ+jKaziX9g1RK83oiJgvdNAya0F29VIl5sgPuBgMi7O5/
DYEHuXvkDZeveCnyYeI4n2rzB5zuZk2YBTSApef43u7gQNYU+ykgTxL+M4Jb5Ykq
DocGGeiPD8x7s5zOAwUEqZXr/FaLLQyPdyFp3hZT9BV/LXVJXrp8Z3z07amdzU99
tdMmt8c05zvbgBqqF3mxvwbnnzbrsrYUMLD2FKPj91JqjK9J39GGzm5rpC4gIQ/L
q3QKNjEdYLF3RBVv9B+IeOipwxpvCngr2yAcy6hcIz5/7efeAw+W+01Jmi+l81iW
bxz9cj+jNe99xAIj8PCHyM7s+RZeCS4VoauqEAI8aVN4cmEvIsmvugc1PMZnkG6d
U3s+6yQ4L7kMaR+SeYzcV8Hijh62pjuLgJRe2LCXZwFbRGV7dHyp5UbvUP06CbYe
DwE+3dP2Ie8Eyx4nyHF0NXghIyae2fQSe1RYnaJdIeUcqlRo0rbtur/PK17H6FP2
Wg83Hu2EAosbLXoa+OmIS/886cixhYbadV1e1ZVqZybjb+c+nVi02V1PojWDGYx8
/YXUIjjJnnPk2/E05b0TMTIOUBQ5niA0RlhdoVmwFFWtH3SkodI6+mhIHY28GCBa
FU2T/Bdy3/aGAMvOaUTakq2AtkVM3NFAFDkCFdh87S9veaymlotUmBvc1d5CEOsr
nI340BCga1Ill+9z4t7fR5cg9JKwX+M3KkPXdnzcxoYTLjBoR9l0p18EbOlW3zJW
U1kC4D8TOrb6eeFfa+Z+JATjHEutT0+ubJlPKEmxpB0FV+6MzLWlxJ9LimaIOF9x
P8UJrj2Krb51YmMiaiEHBSK5n9Opsuty9ScBKbipM7EhLqQ/hrMtrjkhqxF4SuX3
tJyRrn3nEp6wSzl7JXmQpjs4eT+e/FW/d788eaSVujIAP5lmw0bvG2mkAU9Mr9pZ
Sp6j8J67I7WFbeekELUmPtV53PuxII528Sft4G/xgvtZBbnwsGot+d9SeSPRcl5S
6qJKaROPorh3M27TCbwGym4wTPdCEZkqORHEu+xY5Z9XJux5USeaw6pHWm2FiQXo
xHuQwtWqeh6nO8IvgTlCgmS5B9Zf9PX92QdgktKA+lAvN7Xy6OXWWE8ZVvXb1sJ9
qqXHxpbpTXfg7OeEAibcyn/hEPOmvTA3ICFvOgzxI036/0mwhwVw1kkbOL7Cn3Sg
MLkO2QtbiKcfqVOEYcEb0kNYHEztOcBB6JiY9qP0QwKbBwp+7TUQUrddrseqTd1D
IzWnfQrT/pM3aqzIYhnAS8yGSJbrn2nT3sD5+ar/dOpalZuXNJhYeZpQDYq3Naqf
uCZc3tlBWZC3azblcgpI0rru6jCrJOh8ihCpaPA73D7v+O7De84LkDzZrEiAZI4v
CyQhBCkuJ5zy/Ta+qKAzahTUMFIkK2JILNRoDQYo43WTiXWTDsGc8iPP6ZVklBLt
gaT2/YMocGWwy3V1ecA3ogrsfRDtxaf+7P1U55jdEeMM9GhlAjVQyNj0rhuGVOvr
1p+PxA0aIdjOA3Y72WsvgmRZKbkBrNl2OgmW87cq7amB3dCRafuJiYZpCQWIhJcU
AKVX/3aF9l+Bf/tTnlK+P4gUzNxlDwrWj64vxSiEqnhd1NYgZrLtmQCPK+fQXYtJ
j7bM1zdwYxpTBlB9+YwCWXYgx8r1ReIZ2cIw4wRu8XFiSsTwdc/cBtvFVS2hcboo
3FQeHClWle2JkdyiAeyDk80B5Cji1PzGwdA8AXDKMzujfCryA9oEt2ADzA/axD6e
qXOtgEJwtMyX9uQkc+qgLM61F/4fF2V/PqeIba+TQ5/jN487eh/+rXHz6JgG5tTb
ycToxzmnjd0GF3w2KJXzfxFKh1wjQtalaw3cROkrDltEOnWaxb0/TkWrUFnnZN/j
Ese/14/AsZIsAEwUSmyS9dCotVwAcm6SGru4OcGib/vdxJjnovpKGba8Zf9sw4Fz
kRSacjf8WvECrJ2rhVckmPl2rXWV9kh24l8wwRort0HVStI7gnPlNEdcV0hD7yTY
O6fZ11btL18mFtYFD4lXCy6Ag7G3O+mUdnU++4PSFN+x5Qr6OJHxSH8fbfv5qhHx
gD3DD4SnrEiXPedJqXv/wUEolosvBIrfv10tXnEpRbEHIG8Y3jCEZhJGSfHte9C/
94Z0JfCqL40AnLyxBhPKLRjH3MkPB+n8MfuI2HFOaxuRfP7j0/ZCxiQq4wwUBbWV
GD/3Cc5XxX2cWD8gjbIBySL9bXjv0R7uumZDdutJs7RLY8JebS+Vhy9shlNmENQg
89Tk/kgE9GcFOtrMPgsO7rgAtmWERkZ9791bTxNvDaMb+4RIOFzLjV2F3iZim0XI
vXwCr/5P2Me4pRsNWT/26D1Lyq7HSWDGSAvbGaqzIn+uIrfzgsStI9ySC6fbdQ8d
EbqlvgfyA9xY+wAI0hXQnw1EDpSPpXnGTvUTc7DB27BLQf1ll+Ph6vbh/0SXnULn
KIoKFzapbgitrgYjI87YefzhzGho43jg8Xvv8YjdB+PUt7xMu40z1VltS7JV4AED
X6xTRBG6CMJb5th1WvPa8a7V4TV6g9N6MaPMS9VhGJE5hjXhRzJ37zwscaGwfsJp
amIg6c4rideiZAN3SpTzq3A1VlVh4J8CjBsK2TPHG1Otd4x608MpBceVlRkMi3eW
f6LXq6z6rFQIYn9tj+zlBhJFvOlzV7tve3Ni/ULYh9kxzCo9L6U93hNSVb9U7Bxm
GOhC08+fASeoy4mwlET9Q051xPvgheRZrhe/cgcXPyVnK00Ri2v0MXTM3mJQTD9c
cFM9Gue7PeU9r8LOEwAh1hzXEgOZlfYD8E1FUkEDhWAkt/NZmoi90RQHs+4k+cIV
yPqhrn7LTT5DD2UWbZqzziESkomEbFsTyZCr29vz2xGoLNGToyPPhOlrVYernOSO
dfEKFeUPtazX1v2vkESFNdI+k6QHszJd9oM4gL4RzG2l+igO9K5FlxRIUqkNWgIt
ieoEOv6+ELyKlKmlhZK4/KOtEra5Lf4dc2u28/LufADa9r9Q0KPWjUFh7EcH8xPL
GNt8FiVvtFCPuTtIPnBOdSXUgYXzaBLZyRDsY7UEB4xAHLBYn9yeC6l21U9MAXAv
+pRFukzBE+hs+mihUdgqvVQAW6SY43r27ae0wJmuhnoD/d3c+GJFgmFDCPwuGD6u
2LyFTowyEYGYq9ueOivFiLzZV+mKUQeYWNJnVUSp4B+jghg9yVsZYmChCwN6xySh
rV3EchJcldnHr3ZlNtay6Ew6/xh8h6h5SmV9y0fL8+wq1JnnW3ytWYCUhXSZ3TYk
oHiL5R7YbIGPhrMYUGbayVU+QsodmkbDvmuCmOul9NWqYofmkCNGgqJRznnRrJDj
5o75zDbM34ayeMYhIAb8ztmFTdIOiAzbKaRR1f1o427GpzjDRVCU1ViQ84KE+Oaz
XGwUyt+WleWu2NzJOfI8o+fGdixkEgM82oSrE4iJoweMGuNr9gtsjL8USpShm3m+
YlTi2u3v57YrcvLiH3TrwfxCTsH6iBMwHCMrRx57/IXapqKcCEkfXi3oASyfkzuj
53xQnynLo14L+einNDSuu2d/vMVTkD4P5xZrkwmBZuo+G4QEfzF3TYBx/HGzcVvz
XLQfE+IoWnLrcTVYstux185LdhrAXvf3j2qIdZmFujNW6wWjmqEH/JxpoOljfl8y
WAOAE+FBFr7sv2/xek8qoP/ytM9ojeTwJZY3l6+fDvkLouS3Kc2dE4ongJ3LZiJM
YPVlZdHS7iBEwyngnEO7T9K/ZeKBUigIH2vVoSs8UV8ByHJ9nbVWPLsiZzLLdo4j
v5OdYylEduQZsUkFGIZskKWJIt6A1phZtkkqpuMyB4GNwNyTHRu5/0Au/x4Z8VDT
cwIl/s21AavKF+eEv9M7odbj7AWiLQyvV6tDEn738PhjHIYZjTCrTGaL1PMb1Pbd
+XyNNSK/LK3h3YCyYT4RyZC2L3ZvLdYhUd1hO5RscgXU3LOYkQU76iXpyfLtYzml
NcZhZzI9QWBSGopDymBYF3cBoDvWe52PQNWUAw4zUmHGkOgn5qV5j7kPQnulznSc
Hfdv/ticcftyiyL8Rnv3UjyJ80S4pEyrXAI4LtZWCuZJcTV55acxDRqR8QwZ8tvh
hfqnolbJDQ3axOiq6VrjqgSlMt7eQBTUyb77GqViNkIQHF+igiAyGcPN//0YcU1F
iwndgr67fNHzEZ8tX7ha0ogBeY7WFw7F33OiPlXodJZ4/AYB2/1Wzp+dFXdg59rw
LVYlEZXS8HImMGwGM5/Jvh6pMah18wtwUu36MFsq65AwQHIvmOoMS4r3DTZHalb3
BCTiGsj7lqzBCPku30t61qJFYGTmOcpA+RRei8rOnZxeRYIMWraXHiHOuzsjBDOJ
04GB7upxa2wDw46K8/XM0QELqRJMZaaiDqhSc3+Z6GjoSC2c6LJC6JgCf2Jo0Mtw
oRGew2xxEMIxJ3swjd6ZAjVyGlcZLdnRGHfo6xmEa0FKk8uGa2Q0ZwYcJAE1h8/q
CmmWAVWgcSqOYs0aJ945yPuhwLd2hXsklT55nIN2urzm4gI6NqDNv4eupaC9nfJ7
WEEtFFu5OFuUtoWuFJA5FTXWRI4rGU5pAz5Kn2ind3WyvBpZcj4tspvUyKDiEi0L
VtLf5UX/sN7LCvDyuzFkCMQc+2CWsktaFIVO/2Ks3hRzZZjnHZokFQNdV6v1GD97
8/Q/NHQMLSdOVUG3bJhJzfAfEx1kyO18veX6AqGjwwVo72a5HT0a//7SOv1wJePc
AmKLE8u1JA45Ws0UBpvX79TQooLf9vbdZ5dzczeMhFsY/A6nvS0uSUpvSJMO3Vlq
qCZU4NibLTrGhsC56zv2hIRwPiMGk9LEfbb/69KrLhKlXUfWJ4feqWhAce7NKslH
ETSqY75Focu6oGH8ysc1FiFtlVxLCmh1tC+qb0tBVY0CugiY0PRcIJzSkJd0x/we
yBEUQUeL0MqMflK4aM7uIVZcnxx6qK0bKqx5B5TD433kOylX4Lc8jnaP5oTXDm2Y
fBe5mu1dnX7wnEVqInJM28fNBsOJXS8KhGpZQMaNZdccGlpSktDh+Yed4qPLN4uC
1WQJdtI+Wx7yen18etIJs+utWrSUVsYtScPr9fzKNILs8qmB5sdpkaUxm2gmBWJA
SuDonfN6yZrS3AI19yx8Mo+VUGU8KAoco8wXD2jYBOFAGKKggG0rA/Sv2lyaP4T7
wXxbGCsuT3Ap4f+rN1T5UHjTSfgWvaHnMfJWX0olyZOBrnDGfx8O7FZX2trLluwT
ByCyHKqdsH1e7D9lIwErVOdaGQY60L6nyDVrIr5oRRr3WPk5WYrLyTwFG1OVYyxe
p+2Z5+rAhFU6jZuX5pL5ZeTxSsVJfTqp9r0VFNAmdospS8Zi99VIWUxSSAXlTqb8
xR5ehNkjnsx2IeFgPr9uikgl8oswvC6qRTgMYLs4FZvdDk6NJPUvF/Stmb+SIvXl
ESXzfbJp8DrF+vbjTIG8Rz/ws0W5+sLSrnuIjJ+JweWfWV0p+cMpO4fuP+AF/a73
c44Wbnga+Cn0zwk3Hh01LyLNtTtzWB+eE3RXSaRAsSF3pxZaZSEOErWvSgb6V/4h
SMf1rFYN5obPrZb4uqsYNoxmWpq3W8kr0klTMFExw2W5n+glEDc19dEHxmlwE65j
6X2WlhqMlfXVMaEVayY6WFaMoiGnIyORBKvI+99Zd5pLdxbgFklZGXpjBhJLssVA
bhN0yZeIgOlBYFE2RgNJmUhXYN7YMfZIBIC48ybpwI0zwkaJ+hHaFCsI2o6EJfQL
UwtOONAalZEfNivV9ZWdTQWnQk0287dzJK7/Ld00ypFsl4WlZIFlvNM444oIVkfK
CFVYeHFFblxElbFwkqoK3fYbG2SmYof3xlhoRoVmm5MiitF2voywdSEGpxGUI91N
fVELB6iDkTzXhegG3DwA7+jJse6oO9EB3XN3BpHa5RQKU4AhJhlY0gel5LyDuVCf
MoFrrxa5XaZRBAREimFHY6VmznE+cdWb8nwdbMSFfZfI7n4uQSWt3pQ+nVUrLCHm
gWxVTVmUrqXqAta1rn4X0XrYe3CGDFB2j4VmCUtYBLxnHx7Q8PRVz9dihHGq6h+3
mehv/RwZy14sD67K0iswruFjhjB7k+5AqO6xhvnfX/DtSlxx4sYsfqDd6XXuprHL
urAr9B/nOeD9vtffgT+ptpYTMar0VIW/5cZNkeDkC97JNLTHomSm1sUD4WyWkCCE
xnSfh93P8hjHj3PRYLlizSa0xqPAEpKRc/w5uF3XuiAeeul9m4TpvdhvfAU9tLLK
YpdIkGIMh4jqRZTDYas4sVk9hoGq8VCuCCj7Ba2s0OF579TwK7IWei6YHMrFBBVo
khNzY38hUmUqwvDA1v8WPDp2si/nE47xp2qvvOdi8zftgQl19g+5XWwISe3pYFhS
V9d3ZZv5HesYNT0vypYZm81jBlqLgkuC22hPFpd/64asg96Tnpx2lfyc+28HAAV6
Jsf7sub//tAH3EIIKPUpc+Bq6MMQ78sWFP+e3WQSpCMV1JDaUK/6SE5J9sUcpu2Z
EcMzFvhAU513OeiACd7Ad2gge7nd4TAjgDGtew7tx2gPUMa4LcgF7O8YEazjQ38d
443hREF4B91KZtgviS1PL4uVvxE1mEPH8prGOX2uU8MBylNaaxU1H6EpgTl2DncB
sU1ZZsk+EvNtrXVNCgGIZW9v55WA6RpKzgLDGTJCtKqkdZl7gl/m1wN/xF1jltw6
Ns9GbaWWZM/JkQetxjU8+oZgQsJrInooybXY+dAyjlsftKzcgNWhgUuJEouU3yUF
14HhzgurGxHdK/ULqbBHk42vofB1smJ8zdt8oyZglG2VBadOLSeC3qLG8bEoszjL
H2h/u8w2IPvfnOOTLfTFaGMq5rwSp2UKZ6bP2QSeTn0AXoJeVv2TQcZLhzw4kSFh
UK/O5zNFK/Mpg430ckaAZVICeV3Ox7gTQBOM32V6WUrCMVgO2p0FM4ueW9IUSXG7
66fmv/NMfRPmg79jsCf95Du5yIiFkTzQZHyaMWXAW3upSsagv4b4nm4yyhrrnGy/
8WWDrx5VrzDK2feOVOuSsuiCDb6rUbIYjy/a+uSALron1u6gKgxKLFWx8LYWB2WW
zdn0sLzlh/ZBCNUgMOoWkFaVWju/fmvjqrWEgnnXRraS/rJ1yMdWtW7u3Cy+QrVk
+bGfMdg462/AEKXDAYpuq1mocMCLpwQYgHXf6VckDVw6Q65d4tScoLpKf2N1ZEDz
HNlBQkyYwtrGE+y/G5a7j3dQE19SZ9vsHXL3DpiRopA01+hakEi/6g5aXl1hkufG
BfWtwr2dCfg/7I28dQREiB7Y+WvLjW/0stflQupt6Y3auySWeJ0NX7c7Rh+iXvXO
NZ0gpOEdS5T4a/8I+04dw6OAMuYEw26l5ZVTPgowgSjjgubc92uQ3YhjFKl9zsUQ
4SCPfT6eXA4U7WUhKdMJB4YsWSsJE6wYDSp75/MZP5p/8hiVO1Bm8S4RDniEkO2U
7RNuGnbV+o8RoWyx+U34wFesneKx6gJgO1YgqwYTNFsxxbe8V0/e2cY40wFx/1KH
Jbo13ZMfYnk2FGRbq2MDuMX7dubX3zvm0SJIPsci5v6dcDJ2VPqnO32trxCienls
9WjPmWs/Fj8aVBsKtoBCJoMmDS2+L4FsR8bKyscJHWwgwPxVnsetfyRrP3pNBbcu
tM1okruhCtuMpt59m3npNF5miBT5iYu6C87N5rVOSZgp0UtdTzgEtDCRaQcpNabs
uCqhZZ740B75itkCK5SWDf6eONPgWpjzPzEugSiUjO2+NPSrgROGlkZebjxVzaV3
LdyzZGUyyUOTm6s05T0KWDN5cn5DPgil6t5uCyZyrEiGCwaJrY6gZcHK7Yr8TZqm
zAC9YzNafHvuHoxY8BpSG4y6xEwcwkF0d6QFdNkKqG7Umoy3pRAwLb8lmXQSFZ3Q
gab0RKoqo5Py2m5Jee78h4CPU0XUGt9ISeK93z00Hx8B/UpMOuMbHsvRf3nHhtr5
cQD2PjP5h/MzAEGbyHYheNRdRGwgGwZmncl0U8dqF/GU2t3dIa+jD44cpfkHWHPG
vlhsmwKvwlUg8Z4oyGHuY22LaNivlbjXgt+v4c3MpK/8eTnK0Gk9BbZEN9KL3ADX
7/eON4qAXcLi4pj7Mt9o/Pfr2YCxUdF20TXJRTs4zbM6CyLUvULvp6NFm/EhIZxh
kjmlGQmVj9OOgQeuqH8fb9tEKWwzd1nuqHS4GGfISMloJc7GwzwK/Mx1yQP+od1Q
9lCQvGTPvYuNqI1FRv6LkHRhWinfS4psaMpg9NfA0sp61pGoVXZYUw5+0zMnZYxB
ZgeYcD65zaFz/52UyM1DFqzSUSDUepKOvDS4nOrXINI2uFddi6yXEmk+cvgtkByA
KbtjgedXebiR4nz20SGxF4siNGTSz5n7DJ03k3C5Eq5amQqSb54KYzSsG6G4Lc+T
3iMfEfoOSXaNb7Fb3Vsr+sLdM679JtccW2Y78Ob/xU8Gsg/jXdPBU7bJ39YTH4y8
fx1N8ygxBK7jV8PC3vPAnFnX7fsR84oYFom8R7ZWrT55vXtYA9Z/j1hW027HO6c6
STURSg/xhsk/1OsvKVlMh325pN0BUxpaEyGzHE8WgQCrwklgOvhQJFj6QX0qu9Sc
ETH9jPrxZGeetJKs4jI+PCfhn86Od04uk2w3lq7wcKGJDXmeqe1MDf+tYE53oHP7
2OwkispEfdbr5u7jeNyAI6KhD3v9ytbaKHV3+ZrWSdNY0Y/bqd/Yre4W6BJaSMip
HPJYakuUBwzksCs753clSktwrbav/OJ+LJqckQ1hJkUTvyTIOeTeUlZsTEE8D7QC
nMxeeDm0NkHQkgn792iaj/5TX42FWhHMwmzBC6FF8y4LHTWVeta4RW9DF1HMpj1W
gNumA40Ta+gD1Vhr7kh6M5HgtPyh81YH/DTAYd4lws5RvS/9jhtsBOHGZ9JTPoxU
kfxYrWiFamKfScsx6wdiaqhPDsiCouQsr5AtFYu7yZaIp6nQAc5ZPh+33AjIo4c9
+2ORglt/z2MLk7RvvWuG9CmnifEF92RcQn6ZrZUbit9rbunRqE3jR/1M5kN02p57
hSZoBMrvk6vZLkwIzYkY4d6Eyj+ryLhVyZT8Ua8w8o3juCW+DOLDBkqlaikkg3yx
IWjXyBTkQs1+egCxywNaCA+ZrjF5VO8JiCNSBzsdQGFbJzbCYVTD8uRieuUbALcP
HzBGz14FE6uivGAPNvbkVBSel4nFWjbJDOfkletFNZIXG8hRycq70e1SjOGEMIvE
c/Vcfa4avhG69wKSyPHJ2+g0LHJu6cEee8EUfaMe7VcmmXDBp1Bnf5a5LBg15Nbb
oG4gUJNFUAR9j8pPPte/RSmNNJkE6cJy4Yr0vJYGH0yFA6mUUdFxqYoOVYs3MQfd
sx5CgpPPiIktaXW3DGeeHSuguHGvlUaiURt9oOLDflGFEEX0xb6K9vXdUBJMzy2I
o9J6qJddpdJsbW6iNM554cS0c129ATp88B2ENox7Kd5axJWbxKRxl/Ur/iY4vVCm
JRKM3vPwtMdCzkT1yELqyM/sT1rg6cGR2twdtqUV7HOAtQ5snLg7YmLjJLaXzPz1
ZzATL8Moqm0rXA7YOsGN4FNsuxyxQEd78hql6z79s5h0L7yBh7UkhG+qsuX30XMJ
2jm5sfh3ifRzODzxuoVjSe1tPEH0UzUAgahxubJwALOUhh1O+1nyyZa9La2lRR9z
Qq/aDENrr9v7XSW3jC/0+Ei5k3hd9GZGEWODwbhheH3B0Aygl8cqvrQKUZ+FenVD
h+Z5Cg7Kl+9trDBRm/dC3UkFARoFv/Y2nenZBB01rAkexn9QvK4ZGxNddFKmZOaV
48sZ7cKgQGV8DtKkQUYtY3J15zNUeIpvSUk3hhSOtqoA2mHQuXXovw0OMDB4N8S+
DbtL25PIturdgzlMteK1ucbHsLz+1ELdCLZsp+r7S6Ti1Lspy5rYvl3FqTsHdx4M
naAJwefJKcO4Xd5n/Mu3ZgtpB25M1Og9hL/MKViq5CbDZbF8Vm6P4RH00eKdfixL
xQjWZMNdE2IXsCjDNvyIQvq6KBstbP3rnkgTpeJzVRQZcXQO7YzcP2fBca1XXDI/
Z/RGZXan9efSm90J8QdK0qN30bjpvDvHP2y9ZBzHq0OxxA1d7aNucGWIAUEoy2QS
vLVCD8xu8O8eeHAXDDtuZrb6reEM7biwQSpH8T1njpsS49ZKpeTTVLDuwmndmoe5
O5/8fbZb6xCxFrNKePpFV4FNLip17R08xTWSDpeP0u/96VLL34BdSrE0f5PtyrYM
E1gv8LXPMc04W0k0yv69tnUHcmM8GfZ6VcyLG8/VOeFSBwI5Zcu6XQPDoKrtDo3M
m4qDPic9uLcmKTHCmzs04UooAZGCCaaLGOWC5tiinAXr3wa4o0aKJssrWfBAkZhR
9hSU+suLhl5S4KV/C0IgIjJUqRNSPfqa/NELjCBbMnzy/vfriDAPFUgFUmrfMYnz
TLr88lFwauYAH/LV0OV5OX5tC9iPutm/BY+jNh2JICbB061M0XjRpaNDWvz7an6u
sX0KMy6E5o7JXtZSdrc4aGZKDt85DgQYM0cPrCFFr0YrU1t8Y8uNv1xpvwLZeHpe
BT1D2xVOwGKoRxDrcKneEg9egZGvd28vRCtfbOjlNre6PyyWSfFRJzKF3KlZ/8k1
cVhmKSb4bIwPuuapfGQK1kZwRfTODmAfRJ4Zbo2/XLumJ7MhLTRKxG4i7/bkTeTw
TQSKqna+18SBeKOb1wvucZjtQf0x3DDnQ8MF+DJ0objI8WabnFYSB0jonHDLv7hY
Bas4/M+7+pt62ph/Eb9LSVChLrn5ataumLmX84WPVf3mdiqYQihOQBWW//ynEjCZ
MrLvDj0WUUQvYn3+ZTibk8n0mF6eut1QriA3iKZ1DGiMUSz2vmtmBmfh7RHhPbpJ
Gny9sEbjkOZj3xUkAsl/gNfjt0f9aTdJF5bFToFs7Y6bTKA/cTftxmshqL6gbNpl
gSRZGC8gdbEem3dhvvO7/FoAyBPG9ZnWdY5do/TZg7dWZHAg50ngdmn7BORhgBVq
uIZ5amjE5g7HOwjQyU7d4xqL0pxMHTAEYsgcJc34btDVbzkirtiCPSwqTFWNnoiF
FGy6xxe7Ai4eBZA+BYj1rtzV0YQwvcvVufMeAPUGF0zvAy4Ags6eqhRo78pi2x+i
KlA7bBnseLYvYkkCLBLleoxS6/9mQiQdVyp3AeGgIpinis9WefKUXR7CmnjNLoc8
mvp6r+a+PFUw09OxxYmiJRprQUjioYw7QWeFZUJMoQEqDI9mp/N1jOCFsRqLKfF6
GbiwbmLbDMfPqm00hdOmHM6mcpdbyYnytZ6XeeiTLWh1AdooStnhP7Oi2T/epUfp
VsUQzaE8OC4qbii7z1Fj7pWqPZS9CHNbh2zA+PcjtcT+bTTlz4+ZPgygCXAaZ29Q
rbtA0TReopAlS12oQS92Lhz2KkhNUd0jTJr4JYq9aYMHbjlCPtMKoC+dKSCsuCG9
IABZ1hXb+cNwjsOING5J/4He7PKC+lR5Lm9a7+29pxPL9IOxrNdJAFOlPxDMOMWI
bChAVl4DpBVX9s1qss3Ww2NGkKuaG81v8jZ6Ng/WTpaWJnChDIQawtQve9PkQct6
yglAoXH1lQfleoXj9TbloKZELLiFBTo0n8F3/ipBnlFrcT2SOh+t2P4zL4Y3D8gM
jCR0gkqiGmLCeesSNfHM5QGd2hmF2lsoP36PA7IkjDVX/RaHiqD8uPmq/20TK73w
ttGRNCmcm3oVOuCQymRg7M3Kb3I1MNS3kUJRjIxNyeRUZb/FZy2mcspoc3ELdN2Y
yKK7nGwgj9KNvW/M8pKDDW52/44UNHIoA2VXmzblNNCMbUzPR+vA7Is+SqXT9Bzw
bnOGPSyI6RvEZbn8QE/acaxM1rNOsDXDHL/SXgDSyiAHq3bDp33DffTjsX5Sx3G0
O8gDozAIxtN7w9BkyL0C+uYztcE0UKH2cSSIBGyJ9TtvYlrndyyRBxJYHDez9JJ2
De7zIp76kJBOaZK0N0KxqvtuQ0xR5cBIMuTtOf1zLyPXJbkZSaWrBDqEyMxATpJ5
AZL07TAFKDICl28ZKos3S/Ef8tlMkIlbXa301jC/qEzIS1lH2M/Li8nWsq4we9PY
ft/rhMmBFQoJuOu6N20cc66FS5kBi8oCLZ4VW0apsvrHdjuPiP55ocuEi5qg2jRw
aQ3FqTJIrBiwsmVglZv54pHDamts6o9tU1n8r0BghKGmtkuPwmh6qomZ/rdB2xs1
Mo2MAZcMo7xMfU1RfY7jL3BBotrGHSMKpZvg9GXlF+APDYnfFVDep8bi/zmCFcC0
bfKLL2bbIRlIRbtVOICX1Gvt22B4yCN97jmKdWmTGfRNDN9RTigPJzsrJRrkbg5R
9+WyTZpqpKZU4/pQIwAlheXtHCuvWC5CTFmxlM2Sg/z0QL4YZhRmsLxjohB3Nqml
D4MEExSOBFjivQzQnc1RfIiuRsOi/Fhm4RytxrqfqKsSz1qtEu+Atsi4N7MR60DV
AysXdwDX6VzJG4cYSMHmYjzLgl/oJ1IH6xVUf1YdKedOJvLH2ntR+h9umsOB9Gt9
9DTQPHf6AvGbli8TitIDBwrnqUwVP7lwJgD7ewuJ+ABOxT6R2FYn+ZIPf83YXKeE
0AlyGTrFCJ4GDcwlxo5zP1SuPqI4qsPBuobBJuV5qMOq0QzN4deJqpDoPxJt99HY
m+kf8BXe3w22aBE4tJ1f3WGay+bRbzOOTKo0gGGjJ8cc4xlMnCUn6U7D2O4MfzrW
pMBqgtsOh8NDksLikZFHJQ41o8Dauctb89jm3Lk2tvdPiCr5TH4fNAze7Oa/CBR7
dxNP8Qt/YPszSJf66oZJY05v2ej8oPU8HAa5SoLlp8NmGQ8n0ieUXqT2vKI2vvs2
DAPVbAO9jmSZz0mY37HvH3PmcdH0FEDiCyVXid9/CtIVDvkPCI2nGgxz+aCmSrp9
x4bqr49XbUDLdXVpplatPgxDsxOwgjQtLrV0YfjnWmFfKxalqyvTi1BM6AJlAUwE
DzlLWNqN+YAvg/QId7n2TMi1g0bfQTT8KtOou/53uwtqmJj38jLSSEGf8EB39bIA
/CVON1lfiPn/pmboCVX6K+JBWVpqfTc2N/NvB0rznLSyjbZxN41JMLZ+80UiXPn4
zTpYxtHBPiFtYpxxBKMq+0nAxak985yEh1WS8YxK0SbD76L3GN8M8BSWMQxDsi8P
Bu37wkMuCaVvi8iplrjJfF31lnKzjWQ3YqpF2X5grqm5vng99jNkVx7dcOdnr9/D
kOHtbMBsYZ6lTNDcgTQp3fInYgSMQQoyPss8PJkijd7VwG7qRwC/74UlBpPUFKX9
63ZBcTHTG9a/1xuepsStPESG4jkFNLmfQjOvl5964j4c99tQinmg2lyB66OhVkPs
tI3unC5oV6eaKWTxoitCoO7fY4FAunu2Uya0iFQQ5TgT96jaafjNHng8Jz/ByKHz
D1xVBi9KD++qRJp65S6vChuCisGPq4yNLFco5Q3MiGw053qvTCJZUzVyAZ1pi58W
ktQj4Rh9oj6a3rua2NUuOSyBbI9iZFCiuZjyHf51cOACvvuKxY/djhUIwZYXpTDb
HslFprQmVlwc0iUzsky0OuaKQkVVd73Aj2npgTsCy8E4E8tOG/rnMj7MIvdECIHP
Zhwi5i+61dCRPWW0FIfjC+UD4gKp6re2Gei3UXGB4mbJVR3e7KMEGNQRbH3g6fHY
jMW0UBGoC0p6JteQ097gHF+H/EDMQpfp4yjwpBS1zca/gQNnLncythzACtqUoRyg
7+8GGc/bOb8MOpi1rrUtjCTuif9x0i5879gFuVcZ3lVbvYfyPayCLtArHbXeUANf
7S3F2bAhBOcHhiZFgCXKfImG3Ulygqi/VL9FZSQxMvP5/ouAy/RChkOXwO8B7f4C
ERBrYaW8To3Q8tDKOOl0MWV55bBHaWx9jAPAYNscRkKTJ4b2B0JQIyY3O06iq7Gt
TDzjDg5UNv6Rqatt/CtiD79LnuV/w6T02rSiouo3Ap5fb2//9cSZ/DHaOtG9cu6j
UyTDLGzhGEFHVbTPbU0zBadu9jUBMwY3bz4zAymSA+7KOv4o1N3sAX26hA1qR8ng
pNc1xGZwmauIMGiM8cVS9gvXzOGRkcJAE30BNHBrAYIxLixkkwfn22cWIuO6TxOb
1T5ja3ayl2kYT/MWa7x5u/Q2vCFf0WqZTU8eqbVDHIF3N+JvvuySAg5JdHq7HI8n
ThCvCbHCdwTSZ1Tc5TiON2vYeolVIVCi4GQ2JEA365u9ytzryqPrm6tATIcAfewr
MrXdwDTjlHawiZj5D1trMyRl1piHfVPOU26nGoZr51SloCv4GYLHjsn1R0DIKcwM
7N90wvvsX2jrxhxKmZfVjw0wOmHXBVGYlhuOizgXVljr/pw9L39TO6bbMH617h5j
VnNnA1sHMYJZP1OgPL48YALJ1rhhKosgq9dNZaV9rYOGjn0sY24kAWR2i1EGqFfN
rEznictd6r7x0FHREDSzQqw5J7MGYCKgsiMOAuRX9AW5/f4oL4IvMkLXDDcJ7jjH
ozbpGTmrcewNIZIQq7abWjg+uU08Ttx6XyYRotfRZkNZum55uuA/9y5Gm0pw6V/+
jUodUysW+t3Zhyp1e27rU3RKZZdqv/MJgepCFApiNB3IfR6Jq2G+A52mrLNTTpK1
819Xu6m9wIHZMvRORxcrlf/t45x6xMYC4Le7WfWkzGhzmzPLrKXXO7DitCZd8nHh
5hRXptNbOATXIlefLj7sCzJWPP1dOmFsiADxLm2e+tr6kGvBvX/hY4u7lTNiEzA9
Zk524hlAz81iT59xi7dwyQ7wtw/Eoce1MYov/ohhacbqWH3gLLMFneeI3kdQkFrz
QmIU8TAhQLxFRIGDR9W8ncYx3NZzookBfmgbx7lpXkW/o2ZYjS5Sw4saqJIfLct1
WL50yS4NAmpQJhl0n0N09atfAIjwbvJTftjT884SiMoU+IL9ETrmFOVW8TQmznmk
M2E5TkU4A2+a6tvyzp7AJ76d5W8BjUuKZczoYouXf9mnZS4vNIiJqInjBNnJ5Cc/
BOHEtWjd32H0c+Z/t+y05ZfQvp4gQ/nVIqctYC5FzqoDvxayzvtovRtvlYTLRA/G
0PGDHbx86pNVmGW7NdtAKmyJ1OfnaY9NvMdW6ggz9XzCAjgxINDG7wisvjtzi7x+
ZSSCcY+WF2dcerJi5KDveNTYjNeuj09EBmUs7GXi3DKxa752pG8kRnCGl4HrKO3p
3o1Hcqz+XZQejWm3c6MC1Q1O6CIGIfwGXaxBs9kg9pxVPurTuG4yChWLdPWeNQAL
SDnhd73sclC5dclqciMcgDtrmZTA+lXHAVxMZh9VS40F6uuBvejzpOMF3oF3Q85F
EhFFmZrElaXhm9to/bRhTx1AJpdWxeJEddjp2eh9nW3wW1qSCNDFKBeIbvAfSNx/
L/BID0+H48MuQazjf1zk0uaeeI4Lsj5oqBgEF8l06aRkwWgM/L3wgiuveMGIoE+i
hNclFlyKN8cEC3u+jvvUW4GsYP1iqZqzUvJJsdp+iblibedJp6qEFHKqxcMxcfwW
zaRxPPJSB3GtAPpp/aqKKHqehod+ayYO4OTSW1I3SghXnFKiRZDepA2IorOKAbBh
ngiMZn1lb4U3FRzHjX9OXGIRHC5zY4VdQU8MhL4b/3sGtALi4GgJbvsa/HIXcl8Y
153L69QpIxFZirvkw9OvP8h4rkhAgKlDCGYPfGYSoGOLviL0Q1nQCkpwb4jtbMOx
CJRPc8oz3AQyxx2voq8V94di1JLSPLKfZYbx1C/3qbVq0OYPjO6x5KacJxUq6pm2
IiCHjfQ5fMi19fjV+rLE0okFSQTPvv9Qk7fajzGazDwqYqXCU9JMh5RGDQlflm6j
oZHijTtG0lIoBWB5ubw7c6JICwD+1vyOmuOBbliUptFk4sU2v5imOs/k5xya4tbi
pM3OrXjQyxxWrpws/5FdNlaHTK/WXqLuO3sqLlr8GQ9EciZMKBNvTabC5GvhAkzl
uqqMZFWJRgQLXcFUqxdWlh3Gj8cKv+3183Ci9oUi0EJ2766gOvrwc9XZFnU67WlC
FTtxhbSXHJ4s2RgvL9dnvEyAT5vPPwn/q4hv3zUNg7HAd0TopCl95hlAyY8Q0TLj
chtBeMGK7qcPJepFH1Kvz0lBqNC3hlgcPpqkmqbuSFWIAaGGjxvLwegrlc4Ce2kh
aAqpMwk7dbGjN1exoQL77O/vXUhZ6hmu28DVTTn5/Nw7YfqU4h6WqlNLbJgVfp1e
N+Z6/f4YeEvwPsQBnfK+dkRLfufM/Cj6L3LH+1KOFkx7pZOEuVxqi4nxHTCc8HhS
+LwEMkJTFNGNn8512hlY4B3AR2kJNLIf05SITb8hzNMtH2f5F10vzxR3rhoAfLn7
L2R8faVfLpQPCmzi4Y3lLjd9PlSX+KORMlEgoIhDbEsyTHets/6csg535HEEPGiw
1iP2utg+5Go18K0y1eIKtiqpqFv5vSZBLAoro8OmvI7DW07Od2mtHgE6O3CAAFtW
MJopX/jkA7BLbypmxMaXn8YXQ0fIPsxg/5xehCjYv+yl2CbP+aDafHuEKPY7TA/S
koo9pq6losfHLDlvxbiuBL305zVX2XbE8umR16KLn/zXr4Rox3L2G+zGzrmxyRhk
M3hj4MWHhLrx81bHaAUG9kz8FEy+dbERSQf5nd5k6AhEhSSGPZ3vMgCYLyGenjKG
Of4MFuefd8bX+cVHvHQCe/IiSZWDw6zJRC2BvjR1D151ABkTdRyueJryPW3ZK06A
4hkSf0CuDeFnztFoURkqmHGSnhRdcAVjKNzTt0LvfJkjL+NgHudQgZCICFXmGAd9
swWhxz3IvcXN21EvZ5JcqkEjSd3bfEHAOj5hz8d5nxuyfJT+Lu84ghnD7MsJsdy7
sgyIuyq+171sJ8cFzPZdURYJRQV4CM8uccoforCAJQKR1xtjYkKzRW61ayFCrzBE
s2DxVqoIc+vLwQW2xElisMf9RPm4iL8qWq4gpoYm05ob1ArUZB//eWvOcMFsZBjD
q4KlLgw4+gCPh5JZhMFgdv6VGuWpVYMW0bDycpfOnjJsGY4tlsSiFhctH4nQq9G6
p6VRiQb0l6p9b1CECVS8ZpiUay59nNORTus0mi5+z6n+mbiJwUNoRgnwof/Rg67O
gPLdvmF1hFSehPBr3hLU+UI/rwhSe87HEwswl/7BqUvfKA+n6DJ5HKqj9S3/bFJ3
8IFJ4ai7OWaO38z1eVSYK7xzVLC7dThvR3cnhfZ28DiTigsBa+lIDd4TGb+3ad84
E1O2SiZJ4ql0ulgrUIZPzxfQoU2wdqnBqylc5CyyrmTLJVtFy4/NsUBB8IqmtpCH
MK7nE1ni5cpvQPYNLL3jmtqHIdARPH6VBUqwzpazR+meLu/rY+Dwb/VLvce+/Idn
JLBr+R3HZQIlVoV/TRiQ6OCz64SUqVldDEKYZlWwOt1ljaV972FmiADW2nyFbsAH
A7pBj64epRJdGQNsByxeP2aZjKzN9XnvKL/QL7xNp7BcOK/kreqmFdx8faTpRVNq
EuPKlauuJhKqimmIt4DJ4R/S7+pA0uahn3yaMYsYEJmjcz6wZS2deW0pIqezQvte
rNvEA33qtXswuYG6yAX2NTNaGXq2ZchIeJX7h1a8gqQ2kQK2fazsPX1PjoX0kLK0
igiVJWJBlJF2i3/SIYK2g60HWoi9Rxt1B/4Qx6COquBArXoQrI5FzWJHkeIXqThi
5Mj3Aynxol5TtWme+uvZj7Q4l5QRUPSZa5/OQbUQiS8nJC6angO0fLDJ6QoY/DQ/
AjhzxR36w5O379PAgocuGEM5dynPHg4s8vz117iR3lXLuu/xE0xliDfFpNb6K8tc
8GJ4CnD4w2yDPLkz0qeJLjGeKR2QakipIxkomeu4YlUs81mgiZFjJJE0lHTAuql7
SecPpdKZAfdHdeHdXX8wHJnco4mYbBAlSD8QaF3a/ZJX09+rkC5ufFGUrCzXUo66
Yztgr3YjPwd7W7MctRMIZNYFa+0zsdQMdVnF51qTou1tQLUPfKiRbOOJSjztEiNr
libm0bZ4lKsQuvSOnzq6XJJnyt7Ydoa3y9od6lo2QOPEtNb3bNaNaxw97pWmuPui
l8S1Vw1e9DTUIuFNbdEKYgHaqMabagKYSupj3OzhY/ZWFTZ9S8GxtTazos6gxqyw
//+6xsRCtCfcsUhwXRNuMv6HKdyZBGl3vDHgPlPlSDW0AenwpGGGmrKexlQ5MhGN
qAxI3uzlHtZj8j3QXc4O9ojHGDEwu4YGHdXFlCnnVGNG1dWDddUM50i7Yd2SxDdR
aB5EjJGQ2b1IT6BQNUSlt7gkLGQU13mqR6Y/Y4LrKAIO0lNitGw+hju7/7Rm41I9
i3DZERrMlx3ksrh0jMc4G6W9ogCicZTqHgjrpHo16ITYszGPKa8LxE4Xjxb00x8e
SqfAZIVjyd6ndp2faKbUdJK888x/F5MeBnAiYo137DxBdTPRfAyca6OPg2MfcVk4
JDNhyok/l0viDVvw34+FJfYUjJrUPh7upkNOVQyonfkHm69gP92eJzpo+GXO+Xj3
QMkb+GDfBP2XsYjtn5Oj2BxBux+/0/qEmPX0EnI0N3ZFJ5F89s3VVhI+pqzbr3HK
INeU402FYuTvmrb14hcJHDFE3wqIyJo6sRMSC0m+6E70og5xiLE08Bpxvy/+7Ak2
8FkurW2C1DvqGYljfVKCbiAjKTyAEDL7Q/ICaJp9e6NdYIV3Suv9NhkvLZeOuO7L
yNRgdOPXAZmRLsxvRyKgsxVbsGLKs2S9dVDhR3Gc9LnlxOwKhfpDa9hVDW81lhnT
vphvgCif++2G+FxaYlnrR+ZazHQ2S8ZBIiwsUvRV2xDDjMDWwvQ6R7G/pGZBPpu/
eMboaMgQ9Xps9DnJkK9ImExaA7pzVVF6nhe4w9/vmFF6YMNp/noXL2n0rVxyHIk8
UyqZeyGWRnAzUxda3RNZ9S2jipM22ojvww5/nY2iN42BDbKBoPH+Bz+fNzm9LzfB
yLNanf5Kxrt8ecstopM+Md7B2nYS5lAEHtkCiKPHesUoiMYIlmAB+km/fRlbos35
hpYEMGT93HM6Cj7iaBebDKFRsoVM1G2xmnEC5ZoeB/3fZpKZ8FeZpeo3nag4s0At
vuT08ADf90iSN+ftVNehHmqMK8DON1oRh649Zk5LN0Hh9J7DmOFOj2AsRaLXBU9Y
Mh0LHa41oGtHTOQyIuFDKIPmas6Oh79rBFApqyOkg40WbACZQ4xOvlSGxGSFn/Yp
VrCtwVBkbCpzDDrTbYiFC4rRFq3bU/Q1IYwyHEydScplPwz+KAPvcw6II3chtjDw
bbC1R63+je4USUk9IVE1n2Pqg2CY/tIcbokZaw+WoldvvqrF17D25uIOykudQa09
b9h+8by66wCmVjfG24AAOtgy2Fq4lNKtDYM1rhtBrXGjx8Tenv9zcZfnFKUZr59J
pdsT/gpBe+7EoTlJmO+P4ryjBWQRr3G056wQKRyXPPCmriQCTSduYfurnviqU02X
cJeDLi7o+kl1AvdWD1RheR9A2H1J7kgERbRBW3Ubj7JlBeJCbBm+yhM9Qp2NeuT9
HpwqCRe+seVHnx9iFn3Prsev6eG+l3Z67u6vq+NdyEG0HlR1g4Izayfr4H4XwHUi
1QlZ7UQIpXfQLQiUUvsqawkHClw0pido1p6QBdufnka4OG2voieLgqHtQ99y5BSq
PJOcLUfxojWjLhgaoQYBZ225zdoCCqKBf3IZbBBEHvytP2Vp5Y7h+0wk4udcywbu
AiLkeogOSVVEyIKNKD/PQbffQZ/2Nqvc5SjzAbMD3OglVVy92DDH41s+l1dezlF+
MgMA1Nwx0+suf6MGKIFGrQq7uIkPSkBiSXbo1wJ51zpbSDuQKGQJOhF8O/Boejgv
kkwJzIMPgcgk/i9oVK+As6Dj3pSeCcIPLy8B2qwwXQ3t2RMMlockbriu08qQWvPn
idBrcJfHpGRWSn1PJbexqet6p+om+xEqjMSPheydV2JfXu8C514JfyPdv5chX1JG
EBmvrkkKF3zBM55H2Wx3Ukg9t05MYBmOLpj1U9pXae9pVuGlmAAlpK7XwDDXo0Ij
eP1iF2qDHKznbbMthuDLeUyJuKe+JomMTyA8D7epwFF9Ol6tWx68Wvry3n1it4Md
/7Hk2gRnhRMusZsh5s5Zk+x/fAJSWRXkces4NWI05HkgG1CQgspASq/J1yTktLPC
ymyKM1HJcfrEp1pXaRraOFp/M2j5DAZQRVykUAZTfmhMtUqMnZXRDa8KhJmQPlvR
gs42wnwxLnTePLbn3J/cFupbzjfbFmGurWwRZnCXtJ2HQx19Cc0cLePWZKc57pJ0
Jxn0STmsAXj4qsfAiFKXBeMoEn6WYiqicjDHIveTl2W1UZvgXlWrj1QjEufcLzVp
QZhX4aAmOxoA0m8TdnopoG96xhodHj4xd1k42uCJVMSCuzxRQ7OpQha6oGiPOAUK
BzG+Pgvfxh7n2t6dDaaqk3tORgldeHhvObWZLWBTSyD2O/Mtk96QJ6bisNAMmV/F
RI7kL5CzXUgQ6P8c3umNLqNrAl3HkOgvcLNYT/NrDxxkH73wZJL+Z34N0iyj5rIX
vACEAgqipwhvI4lBiLA/OnjIinhKhNxOCp9BmHdFH8d3euLlEKTljLLldYt1B9XG
cUi6evrrq8YbQ/oCzTifsr8Q2TKRmgXofeXbAePaX4qwbox6tgSK1c6ku4TOgD9T
JQLBEo9cqazcBXpfkxeaeeLDuah9ayQd0R9JQgLmuGlDP9tOUwsAH98McOOWs6iB
/kuU9jGlL3OPP8Ze9zdui792XkMM5D2x+HwCToxoP2ZZVNSdJoarH/nOzAkwxclT
QdA5GfFD+HkUsP39ihEQvoG+kO+/FiG8SJ5EXQtOOWhkkbXM2RboZzwipXEdAGS3
Ifw1Blwjqh3yH54WAH4kHOseQqfQ31fqPEhQBo5GSoCGUkorxzO5KH2pAlpxDF6+
8hzYA/W0Csvgmtz+dZBAvBC/cEopWP1dZJNYnWNMSDuOf4H0ywPjOwl+AT7I8DzJ
mlp5LP3C/PlzxKd2DJNLJ9xzNqI3rMpAjuxvaoe4I228nEzzP9yWu5cAxxItJeCs
IIf43SQb3Th7JNDR68MqOTq7/K0+7m7gfnVok+bgT1xFnT4A3OVsrcoYINh7pV8d
DFC1uHxRosc3qv4xgKQD5/ES2a9Nx4U70IyEUxPHVBn6uBWO6pmtc1rCagEEpdQF
ns4OAQXpamLoOY7Hc2FJ7g+XzSGtjDoUq6A+Hi24hpeZXr/3M4LM7fTd7LRZmByj
JKzK9jW8tkzPx8rQd1Ti0ZrLstspEALaqr7mBjutmUv1GpZ9H8mptwrD7Yg8uKvm
UEEpSlIip/NlmvGQ3edoLfJczsz9Ws7FYe/jnAGch5/D8LM8IAfAFEP9z2fXws4r
KYoUWEQy95jkq9tgTDP55E6pz91cCV3uF8Gqnr2MyhqAjHfJLTmF2tYlaUWSVdxV
h8Byembgz+VKexV+0Q4tjMrU6QYFEvGH4KFlyl/sOr00hsklCBgD/gcNJiC4BsQ0
9/t5l3zg0fQ9zNKcJN7VLbkQqIC+nmCZQ/PUgo/PPrZUn2+WJEx8NDYpqOlSHssE
3DCJ2AaYIyn9OPSrRNxihojQtHvHgWWKKettXxmH6M9banB1AYaalA0zchBwHmVX
jAHTkMXAG+yIUzL9vWmdWjuAImMa2yIVctr6xqGaJJfNfGJtw3mfka3PtFz5yYAS
+oY68hexAsGOB5JA1RrBMsvfaGJw/gvnaYHMncQ9NOjNcVKxKwZkxqEx0+hQ/Fc8
BcyzVcBL/RW9Sk+Rh1Nn5C0+TFCdRYHTil12ntQkxybVUj7um6ISunarYT72HLvX
etBaHJqGNJIOhcO14jMyUv6z4JNs30w+P6PRkDsRiIJ28hsS2QnEAkjzLrgVm/HU
u5DYWMVAa/nVNPuG/+mEUw7I06PwaBE/hF/prda7CK40GkPs6qei/uwniP4p8UyE
5UlIuu3RB+Tj2N8MirVg/4ELcVuf1QBGhPWyz3v+zwGqrEsl3YhG8OgANva1Gv0w
ypd9IOt0f+3RB1qOUO8T0pB5RVO5EotU1GBMtx/unW9FOKjQ/9xDxnOQzaobYB2W
AwdjYwa97vSBqhHmk65FvD/IZqwpuSoZZ0J7kqU2IQen5PN9WWIEg2ZRSO6YZGdM
Hz0um+MRRQ9X1ja0opt5MebDqNw/AQfyr3oBEhNyMSniov/a2mqEGN6ERZCIF/57
/7JiZNPKMNjlkiLm0RZHVOxthQeeMVVUs/tHsZWhP1qGqSupFPWAmh1PKRTgRUb8
YARjZ3DoS5JRuj1fI/yJt4fO9yRjhEbiD5av+Gc/4Od0edayE01XXq7VK7Jlu7dE
eS0yAJl0mAQ5nmKNGCNTW1a//+gfkT1TteeRb8d3oCZ6J/ZbaDDGHqY3YTjdpYSF
deUSqqpMvoAa4HBk72emaspcVMoguOOeciMCF3mLMzyyQOhn/iSaRXOl3XTt3tkz
x9s2/xnUsvAxZ/0Bd+lNnKGMvlSD/GO8epaShY1nvwN6B3rn5Oiui34Q9+T9idLE
EHIwTlhi9UtdJ9EQM8RhYoeoFKifxwztu2EOZLJsW0lg9+YHoDaNjpwbTkt7Chfg
qmuDo1qQv8yaEl9GwUyGkGjAigRgzUAf7Qj5ri3Ybf9BUKhzhCQvsh+u0ta/QVbg
2g2MQKkORIwnx1Muy2wdRDwPFRj6oFOmUNDBbssdzj9THpurvN+bKcU8T/oe70Dt
CjYky+VCzX8yauRCbt5ezkDi17wY6TARoOCl8jNOpWOZULk5hNX5ABk7VaKkZXXZ
KzGkc1Os9UHZK/wedBiMYW8kTjrr6JXdf61lxT+mqgamtxJVeyJnfH4lShvbbWW9
s5pwscpZiBnaHIOcqkCsfGYWZqBe3E2ME/uNsi86ruo63tFyOd5POsVkk4IW1KLK
tAree5rPdSpje4XX6rcMfVIJ+9V9772GbNGMO34o8H6iXORLZ9UjScfX1OMGVmiq
3iBeuBmop1LvzWT1SIScnEdRZFoPNc25ZQxAFw3AZctvX3F0OM81nNAMvm58SQGq
3LaGkUSHaWtxEQ5YMsLAr84u6hzBlUEs7bfE48ps21sTHZqqgzqxh1iQZyFVDCCi
BhqPLyf1cWXJZxfw9YsVzgYTUzHxQh6S82QRUUYsgrMBECr0q3lXVcIv4/uAEJE5
am0creA6M24DleADpaLtcalZYpqLkwNrG9Nwh1CrV+8rhNhYbSgJ/74lgMVQnbti
llgbiyWz19dRiAD1hkVlX9RvJoAFiuVF+XlpSAi3knO8wiePXyXUKdjLFVYNfC+U
jQYz9CEMGQD/7BR9mUN+PSTBEPXyFriCeCbbPx570bFh7iTXM90XLuC36rdZNE8X
+AuO6Rkns1yEvCaFkq3v+grOE5JiRL+cDq6C0TtrUtl0iVqH3CTMHddPMfAUt3O1
yVm8rIbSf9l3YGi+xsgXO17BXn8H66QV1xsMEG6ysNdLeRVPXdIE+dV/k+OcpvPE
fXiAVSIRTyoQBI5wfzdI2Ctas5csQhk8HPoakK8byr5PvvMpK4YpGWa438HutavV
gi+epmYggkoz/1BXnZopt7hkaep4Xssfep4OPmAoi2kDR3DAZ0vevp3EReNdil5d
2jKuLs/u9VbNlAzqoG+tq7os03VYd0Os5ujUkwKSclY4FbImV2fhdZcjsaoD0CSA
c4hD0RhGR6pTXe0+FpNyqYq6LkJD4xuM3KgKZkaj5Vqd/GMXVpX7AMMhC4yZkwKU
/RHU8zXUKE+f6iGJHOpGEFaIjVjzMPvqnmaYOFKEKklzWxHqYEVWyO/h001T4S+5
8/T/SfPqfxcAtmm3KOA5mqjC3Cv3tju3G6rC5/mga+Q/Z3Zwacw5cNj1rwveRNtm
rEG+fnDZ8tp6f4500xamExEaJKwYHSebUJw/HtGrgbSY1PoRj5famXMGGp5dHgp2
Ef/bSmdpYewjErB2nC5kZtZgHdcY5V14OxaTbtN0Y8DClAqf1JQfP4pDnajMLhSm
g6Yz0+cPaudYM1W5fJdXX3iHqpAkESGxD8OTfj05uuOsYbymo+i5hXroeYMXk6cX
4nWQ9tJ2bZpq+WZIfWwwW8aNQKJKcMYdX5IcX9QfAtsMtKZUSf5SyeAecMDfYpiB
6844mMLGiVP0AcgXt+N4v6P37YNlkZmi5gZjt662LJ4aXjTVfWsesHFeKClvUWZG
7dOMn8co2vUh/YINr3HdrwHD+TefmjOngQ8Mw+KOJvB/LFxHH2QcoJXFXHocRRar
a1VGf6G0HjActPX/eTWGSuAMUJEhYBf9GJf3P4DIrPft/nn7OsPrpBBZyL2zPUlV
n92bruH+tWMB+RQ2xOfF2R9uykeI651B1DzjRL8Z2pyLWPsYu3WggxHBuGJ8R/Xf
5wiFu4eI4acAYCqt4AZAdrr3vfTR/BqyHmz6c2o6Wimi8Ki74WBf80EZTqzEOPfJ
uH7KA0YzTHz3uUail4Y6xJKNp14X9Q3lPHet8FYcAToHupApxpoYSEJeq3qv3LjF
BhVRwaHvRG5yKn5yl3xYcY61titJxM69o8pPn4o+7LW9DLXlFFiJiQEIBRX6cgI5
i5GJFVNpMIGuiFEBE2YH7dXhYrOxDTNOQJOBqx2gIkKKvVKzEoQ60oQM1anFTHGm
qMxcqaoOK03A4lPY2XuV3YWYfqWqKgGJv/AQ/X1OLu7ksMHIL1AXaOj9iPSTzfOi
l2lL6kB7tIraYC1BoUoZ02uYtx+b8eUNHB+pYyyuiHp14KbM/S3eZVx6Vu5aZgKC
kxd6HlZiMNhQl/mbQoNoHy5s3p+t7K6XgQr1h2Q+ITYZUycyVBOttnvtYfrcs9Lt
d7M4q6Dlw50hC5GsmSsKb6NLWW131lU9tQ8vEvNuCbVjer1mP1nKogyIa+XcNdWZ
mfpGQHYKwttIlvHdPsE1/mW9LLl1lWjVOLH6C3PenZMQKFEQ7k8PHoY52vJgzj4C
Ml+KfO4G0FlSgKRVvUBpbxwevmj0dOwIyBiJPHJ87/E/28KMLl8dFv6vZiYahwym
+3w/M3r20Gd00yin2/NIHfkcqVdhgKrYHyCn5NmwKfvtgAcvzP6Y2Lg1rSb04JXK
AW5ExgeptcWauQYv5Oz9YIT09g81uSHfZYUYBKLQ++rrmMFgxJ3cplOT71dfqie3
zMENacInQ+r8hqTQfbE3io7/i1iuVpVCTtPy0Z2GWtuFjH8rD9XWf8Y4XoO1egYl
xDmxNHBO1YZs15iwh1FLkgmfkzLfiziCO1SgvxU1VHq7a4r9nkjRLCKKu2mKS7rk
AQerZnBltE7VHQl3jsR1mT02GR9T50RzlK7eDzN7vM5Hbc2SXv9oYuSQF/bG4Owg
kxaP0Q9vJHisru4VDBGlI7ZGmhPuZliT1YwdijSCsO9g5cYikQ0G/mzgOr9xjt/9
LglZucmPX0p8Aih1Mm3N3pY7Lle82/NMQV51dM+j0KWPtnh81VAcc92vccuVpxwC
MaEbmBgWoR6DQw/OQ64Y1Bz6jJNERdnMxYKjdbrhQ7CTA28CxWVlspRzKg0k5Pma
UYvw4h4MSez0RtraMjQCqOLSuLz4dnWeZCMv0abIqAbWw7NaYQcIwmSZ3F84RnIt
O7w7k80W9cCRrZlfuz3yNjd4het7vmoZLoEmdnsUtGiPXS8NXkcuoFjb+eliLL3L
RaNRICSDwmpk3OwTP5GnSF19cGdJojzwvTM8LV/GKD+Uj89/S9MP1PYYxW8S8BJN
VAcy/xaU7fRXSwRNrwqNIhZF5teHztR5oGjNnXwDMV51HWHTRoB892e/K04affB5
TRxap7BiX+oZ3KLI9VQZ3q99Txw4W/CTZUOqBUGExwBOmw9HDoLtSP8eoxKKi9YG
hx4LmJe/XU+TP9NAfsm+uF7cOFAA+NsEdrd57Lw0NpKTOdYDZep0PTIlv35HMiq6
u/sTQ006wIN60cwhYhPJEhjkDG92Js0OuJIdI078iKInr+bCTCsYJFlB1XZ5S8/d
5mIthYDd4DgpLQybezjYxLCUn/Lvhck7lG0xHOn+Dscv3IxXZNyvXnjJPNl6pK3h
uyLAfZstPno6MzSko70f0avD1Silizyt571NjcisRYipvo1bNJcuL9aS/VxMFhAJ
5ZTTULwgrVYeWR/c4ybKoQxAk/+H44QBt+FdrlO4RrsvhSUXzBVV3tqeyQeO98XA
wxk1Zk77XhWh0eLX2Cv1YnWjlJI8VOLMY2pGIAXi+mrph5zPMzkPQpQLexTcftM8
4WeY9ppqbUkQwsl1M3spUDK8dIBLCb2/987RuPX8CraMw746eXzzdpsKoaLu8pIu
WQ5BBkCXdgdvg7Ur6mR6MCEniPewBSBIVGuDKGoh0dyFXtBsQ6snfgV0bmkVKYln
x6AY8G/9l0bYZJijHPd1OFyIHSim7NTRC+svCXuOo0PxkHRoCeT6lcBkEo1pXEmg
brtmQeCcIOgmxafAVwpb0a5cYWb/3Fa9hS9kGT4XxqYe/Geclr0RWGWNdi3ITB53
RerEUAdyn2XqUnyv3YW1u/49pRUp4PLOIQ7HYvu0FokYmFSpb6rksmPap64uZDYv
Z14bbzEELsaOOHukuvpLIf0TYSPo1U0SnSrHHnKY2ujPIzJE7z1eaVNRfQyRvvaS
mtVxCr27kTtEDEvBcy907fxHxzYdTQwXKgp76rQGtaCmqd42GIy/rwP22UigGjMT
ZNMyZlwfknpSeMdh1aq6lxtzaOxsBdFjVTG5N0bBUs/mEtJETJkNxzAGOuzj2yJ7
A1RU6BBB7mo6q1l5An9r16yRdkcD3YRU09yUdvonv4dehwfLylk+lz7wg1V+CWLz
mqJKGc0hgNyb/waPmJwCG7GHQZFJqaddLzYgvV5i+EsCN6Wys10yQ8TcAZ9/mO/y
j2SQUu0IsYS8RcaB0+v4eaoYgSeRpuPt2wotWv13t8QFQoLEptOmuJC8PIW0B+zg
wLeRyzZ36zyiYwwjwO/Klc3ariPR2zpZdtnTxHyJNj99o6FHzgzE/MFKKglC3DPa
aWgot3nHKlH4F+pxQ0EjU+S3z2LWagQa+ModKneGKwJd3XQA8LOTSa8V88f76kCb
vuQWevGkYpcckAPNgPk3yNZ5gfT3i4Sah1SzabdkUfdSKXIWR1age9kvN83YwZao
ZbAFTEWRip/l/ufkrmpgc0vkNgjnR29j/7coeViJiCIR77WJGtFZs4uUOrmWwCVd
hYvQeS4UWcjgILDAE5+HOBBD/H0nDK1uqXIZhBsjvW4FU1B7hwENg9qSQiG8eu+Y
iyxm1bxv6kbMeMuFANJ6l6ixR/RXFt5iVoGdUdnIJxngYjjkx2E68cs4DigaIEqU
ca4AWU2b+1PoFJdQRICRTBHw0i3/KBrqjH/JVEk/eWC26pvw4E6dF2tuKMzUdxTM
tR7KyZ76IDW3kh01+UAPnYSsGf/e4oZh0L8qWmGXLPNeI7fhEvA7oCY4ChyKncG9
Se9T058N0/4FUjLeFCNEN1hQ6lmZjOWzacTHKM2fe1lUjhdsBHLVrJ1K4LAbptrK
F4RBIkWvVj72PHcG84LcA5IvFA7NfMY3kCHruTI/V9RorMCTjiEGwovd57SCYYnV
5BnY72sYBpeQ9/pz/GHwHPJ8A5T3X1YmUc9uodaU2IO0vGBYC8Hu1PZ/aZVoQifG
ka+ed0dppkOTpVHyWP/Xv7cITfrrLKBGZx/avDSz4ILnNKO8s+oB7QPZm/jI4OIY
OlbqYrw/8B+RwVHxojTsZplCOGgi1T07MSFFzk/zorbHGbOi0KqKJhSZ/Dwq83z+
3262fkP/fr5fpeymbFkJ81DdnPHguC0H2cfxz7Wj0Pfto20eSOKzRNOcpeUexR6Y
Bdqf1NlIc8un/RsUIGFkaWNM9nRCl1CpYXdCdgMAv0WaHvRmRUPUERQeQoBXk8Hj
08UFpMrZWhrbG55MJm2sj8ISbjySxgNCN+p4hR1XQWn/WxszxDKj96dHecFrheEU
HqtJPFBnCZEL669U0IEMEJnZA1u67B+kTp7KNuIOS9NOEaBwbDtSRgR/1OjMgDdZ
dlv7ZtbX36jaJk7vCByXvgbHn1od58qJXSrVkZ/D8uMcYoLSAfqW5C5PlEz87n0z
1PehohTZW+y7NPmDkx7Onsr86+m0pDwvP4+N4o5ZxMGc/e/MeAiIJDPa1DbkYZw8
JfCF7rt3tQar24YVLWNitzRTELcw5LYpEGAAG/+S8XlW6TXyVoNu2Rhu5meR/UGr
Yw1AEjnq3E0U4n1k1vIetrjtU1xWENzX2FIwhBrOOFGJ8ExwOoM2vZU50pR/7BuI
8svQpL9envQJgXpAsg1zuW3QEvTvTKhpcr/hGu9N5W+ZRkNOGA+XcEma1b11RLm6
7s+UexPGngRdDciRoFZNkWKWonTAqO3uIeboqXbAAUcEs+AH/6+rG5Sros3YlGxv
VVqiUqbghYuB+3O1bQAaMPRdLeF0CFmfeBDtkDFZ2L+psnUU8WQtjhe3X7ORgveD
x3AhhlzCUTvLO9EtYzVr6FKo8/1OasavXXuoKViqdbrJSlo5jNFyJbES5Wgzcfyz
S0nqt1wUxF+mWJKwbgGJqL8BDPXJnScNxmvhaPrNt7apZy4zTvDkch/QQhHx/SMT
9IsUqwyGmzon19LHg1ezM1r0s6TiMnS0v8YyzhdAdSX0TgeRy9clMyK54exXkbWr
7vy3c4qxc/ep0r2zKmWOO5dJl3pzdPgNE+TClMAmQ6RrO+Imzf21+AVCb4fhAMUd
3y3AA4wAvDNqVpUted8jmEeNXpXAJIRrOWty+2WraAm6QCowskMKUSGX1MxQ5KNY
qg2cB10jYNU8PTqbCpXEKYiCYXelzhZKiWhd0TH0c7eGZNVtltM6P7ZBqmtdsae1
Gq6P5XjCq3yWz7fnbD60Ph9qBQKh8fuAl+StyrY//+rH/UWLyiRs7llEOeJUlPEE
sQ9PzVBN9mcOjV+cEyVH0ZF5hbL3RM9ZF2clhrpKKJbmkSaXAspVDHCuDvgtahHm
vPG1T/AFOZlzyuXzIq9/VPkcduaSq0Nr4j812c9uudqLLOHmtXBnPKA2xJwBE2Kn
Nrxr1PwXv4mUpgfn6nxO25ZimOjqQFbFlM7QVSAC15TJ+qwds3XuT5j0XpBzY8Jr
qtMn6ZP0jaW2RTfYyJuOJl4R6zKP9ZY3c0hCO4lpbk2rSdMwxQ4TctAIZFIQjNNF
Ul/IZIB3loK2WnuueRocFFzjal8UFARhLXpUn9N8+KeKyjR2jWOkRc1cyaOoRHcY
XV6C7jZMGr3MzC/9S+9I7WDQT6fJzRS39HXm1N2IEvaz8LkpQmBYVpQd1EkA7q0D
L33g2MMlGfttopAHVJUFAXll9pxdThQsDGe+qC5SVHG+D72XUX6fiAmgnj3T03QY
FqYs71MtcyvZk1wpwosivnXr83AmSu+L/Io+ZpxVefTqs7C/1CxVWRiObQ65VFiC
Qd0lWCYJycOF+sr/mpXQliRAZoQggwwzVTH3r8apR83u76f21uSt70DiNB0JuKGC
skCg2ppHEggC+RY8aaqa0Z24kxN2yErVreY9UL74ps8A0ci/ADrCn57msKqGvpP0
HUyBspqmHkLn2UMTmgyW1d29N1SexVJiLBUs9M/hcQAPFIAtds3Xy1IH/X1fgkZJ
Xc8h/gMxF0dVld+qjoRAI0ckTgpOCXcMXi/IIZ+q0rQ+dCHiryUf8VgTMcSfV7Nj
q+rkIv415S4JQU/mF1ABCpamv0RFHR7xvTD+5aowOCkAQnc6gQ7EhVhGkxfJA3QG
Eqg3D705oVFYLPg2hB/MGClMzz4Lmk22TonjzrusUaqPWoqy43JBOpVjzM4mAqVG
wSpKCg3weSPm/5alwKkrlRavgwlVTgg+PVCyraXa0Ylwnllo7iVR3teTQ01pwOQE
FCrd8ZsBf5HLmp/bzD6cd8u13QJknFT0eDjdHJs7RPqK40a6wocRP+lzteLcYIkI
TAvjR18b8h0HPohTSlQqtm8hMRnjh/602WXau39uKO/be+peEqwFtat7uqxjDWBt
0ty0td9VwJ1XenYSzS8t+V6rIhezPMpdnmneHwTd++y5f5ZfzWwfXSHTetnAqL3b
Xnd7CR2uyAhW4YJaHGDj/v3OnWjGXMcMRh9c0BKM6ny3E2niov7l3g9mqhw9XxSf
IjMzXPL+GOve2A1U2IJ8XEofAdla09RTR2xYvcfJM9QDaZb1DmHSNvnNJ886/4qN
nzXbLUxZSpF01WwBZap4pjOsXIbOkss39Sw7xKjTNzXfrIYY2tfN9uYtOZjvfce0
l1UIE8SJlY3GXBl6ykxCVoMNJHvAGnwKIx7AIaxvYBxooJULbD4GtYsy3J4F78cm
ddTdoxg+8MDda+tJQswKmdvhmdAFR7liLftnekxrNs6F/h6zi/O4ZY0PcPLtF6Bs
zn97tyagmXpfPcU+cSU72S15ldgzeR5NuZbvF8fOQ7odvicbf1/+1EZMh0IE1r4i
ygIThmYovEKwyVqtGXWRGrxhNkTAc3mPGGHpFGEmbJtkrO47vrRjrRuMLkwgNg5r
VGdHxz1BU8GxwSMGBiMepG8OV6kGEEeri5hqFiRytuTpSp/8SAtU0SsEWENw/L34
mxwfoxuFpQRtbEgfkdFd107Y7CuhtIi+VLg5aCD9OtYmmQZ6bCIkzupnN76yMIVv
jG6EJzHb4z2VlnVj/x+I0oR0yRDd+0IhxoEFerNnGlphTcPMk2BwT2HvShrS9vnV
Eb/5Y75kpMD/cQSKjOBuz0V0IEJqyCcFYl8LJ4zf+FeDJWlNl22XHkUpYt6lngjs
HiCVy/dKj9/gq3tpR0ZpyGGXHwLgedpk8U+UX98hwLTtWH4G7PTSfP6RdYuZwozk
ZGKSu9DB9x1h2Gpze9KInEpF8UVw0Tqf+vJQjEBlrUkAFi+VN1t2523Ixk1bogWI
nV3dsOraZy7j1R1kBxemtnITUViY86fpj9e4TS6Pkt+A7Phl2OajaOwBNrRjPU4+
kR/hWm8jeP2w/10y3t+YlYtqZlAzhlBpog8xcQbz2i7yN3qkbSZbkbyqEmfWc7nF
2fmfvDXU3RWunwT6zQQfw52YJtPrxm0nQ/WS4adfjZOF1FFTxghBFn3AVM4FpSRC
cejm1fMcephtiE3LlF3WySHhuQfzeOiclPIMENkssxcMdQqIKHHY0s66c5xTXSej
yfkXPClKKpQAlF6nkRpmOot0lQxjXdaPB0zJIxIteGDojIJNAjsuYWiNwwdLjlIv
FYwOZPiEPM3jAtos/Kr8vQTOgZJhS0KHtDg3Qk9Am/LH41H0aQa+kLPiI1D01/xA
wNkalyqdiTOhAibvaZbvnyle/cUrdusZcYs2NEyI6+90JGghY2QZFQz/RFYKRzbs
+rtyyCfOIhkWXT9eUWI1Tm0Psa5Tr4ZAtYMepzEWhylpgSDQ+wiz6rCtYy9xN3Yk
lixiLfhzze1Z3hP6Y8RRwinLg7FSy2VtNtIr6aNbZP2Vns4kjMs9Yn/6ORmJPGYy
BOLjAe2TXl6Fdimxbu/KPmDtq+/xyLHgoIGYh6mPK+2Cmxq+lhl1X+gUW/KlH4WM
PiZG1k+5mEhXDsx/YD3/uh5hj71xRin+lIAbhEah/vUC5Yybg+9/Wn28oegtHUOb
TaTHOIxmGz18CyhcBiPh+bFVqm0CR7t8iASuXBmrSTKgUXbBu7s54CXqxhvICotK
lrWKqtY6x58veMdsvNrRc1esWrG8EC4O/VB2yAJFSHWZqTxRrjuarVyyed4B8DO4
usDFEX9v+gVFYLTfdnRckr3pRxSBAQZQLSRIopsg+VjHBR/Ww3Qa6yfSI7Rxk2OQ
yfW7HXKNDTA2sNUOSv+tO0nrbDyHcz7uEe31du0LzpTM6XlfsTAAVsWdFVDFsf6t
EliknqKt7Mj0OT+jMCPPBCLramoYjife4iOXV2bncsjLFdBfO+GB+6XNfomP36+7
o+GSr600lfvnWO3jUf3M+s/fNO7nklo+s4Lc0tA38Y30+zey1l5phG1ASvH5/4KQ
vVCTyU6Y5yWtLocQ//jaSk+S9JyrfbjntypZbQMl66qjyip3mf1TiKIka9GHm1VR
USd7AU1rzlESCqFtWUhuFANWcPVonSKZzb3m/kmQyPYWQ2IhimY8Z8XOEGckn+ru
xvvW1htU3DrNU+nooX4bY7a2BXQ59mGAY1PWoMoK5rvxCRNcRjynO0SKCFigUoOb
P4nYBv0TYjwHfkB29gsRjlLe0VjPPVtm6JjAJRICLhVuSo2kIjSYxuKSbSzEEHl8
7DCtIb6RwBnsJxZMxBQ9Qg+QExBF/F7N+eNM44JWm6hVa8yu/U4m8I6xWShSo9/j
901k5yUNeFd0VXiNhvYu6s3qZt/4lhZcmvGdoHVe4KqAB0CWlCDSDD1n3fubyvHp
uqygkyS53bDNKpTJ5HVEusacmtCi4hWvcQY4o7hw48ADLXAYyqbrTjMWVMQ4EU1d
1sW+cClg3wy71g1Bw7x8BjY6GxTBgjGyqFhp+q9/vcCfttM1OsMuTXyqbONs1fKE
ySbf2OqyW5jFvS8eSoWX4zhER8rD2nEFPjjJnWKvOYLDkzsYwwto5Vn/Nbxn09LB
INqJ9ppQ3KAdpZZzar/PefvUjncE5BcCDPi7YmfUDC3FoAcj0U0gyQkQ8hGrr0OZ
luIT6AUuO3Zva/qhyye0AItHGUuWbc3WTlF3g7ed5bZiU5/PpPII7fw5gLl1VYRI
iWJ90riX3AH9o99TZXWBnLz9+12ctPvIgXSg9bSkw+MoGFh9dMQ3ehEfwtiXnEMn
8dtSswjli+crkIKbioGHbCkbyfrhXFO7ofAFd4lNmqc/HNUXCJZw0wT+RlHdC8LV
lTGFjb26RoRvKhRhkezgAxMghB11QJf3y8+ZgnvQdeTfgBrfFRP5dZK47LNsVimw
DzFRaLitYiP0IBwbHrhkVzjVz12gSzZz344ALiIR/gRDcAYDPmUH4+WDtDjgsqUv
QxRVJyMQrbdkin0TmDW5RIlmX6ckiwQc5YQB5GeltTQkPocfQnUs6PTZXcoEayKw
w0X9805UdcfpH1QzCPlkcKBB5Hiw3KOqjgl1jSdL1D3OphOkkx4XM8Xy62lBYMJk
Gvna5T1hGetu0mchbTz24CGfPVwbFtqxmVa4hURnLLhpGsmQvI+qE5O2l1RR7cMS
SxyF+S1Te1kXOhQdzMYUS6+um+9rrIRLbBOQTxlrjlmQO7X9zuMHpm9YJQMrbPNR
VjCSVQ0Q2hBubNZgb1bEoZlDx/+0XE1Fr19TpQ3tL49Fiiv66WArD0H4Ggid77yL
X0tdfKYou7H3YkSOEujQWUAOvEpvB/z+ZR7vegLPiPGji3V4y2sRwg1Ik1XU6Udr
btr/GN6iWFPXgCx9zWEvC3BrdjYB1bpWjRfS4WuBh0f2S1X5JeS03+XhiZygFBfE
gnLhG6tmSQ4VY80XX8GOz+V9pjfPWYfL5klccC2FXQZ/EDSHNr8CjURHW4oLZHsp
qxi9R3GMA/ynX9nlR4E04GjGfn6VKZnLGlSJcKa5XIpi4e/j1+jK+ceEmpyaTCHf
E0V5Ks+1nZgKSe+hO5y/Weeh5L2p2VLuQ5DhPZlySHhn4FHGfdf8wjKmUQdciBc+
P/DPBfRbmwQDAfCEfYQyVr/bvmpRkmSJdJY9lf5snDYdCLtHtUCCSaiSeTQdL5yC
4xeUGGBzWBXsX7wb4sSyrm5kar7ycLep647q3pzAjWMEmVFYrO48dIoSqR+QKqvj
M99mEjfrhT/5aMNJw+64Yf+ty6RkBg6dL5IiARPE73k321InZHffQ7KU/Khn8wo6
YXZQcQ6JZ6eqCns635hIJml4vW6Zuk7JDNieOAJXhRXyfcY8JU5S+FBUwpx16IUo
StoQEUdsfXj9SyBgRnGNWs33mqqbnJQ7Z9c2VW40REnzN1qugAr1j1vRCrpfxECo
+5wotUS+KPzxw1CNFhSMhEalHskwrtHDGqa4a1zAmaaa8h9j/JDJ6PmN4g2irjha
AKrb9fWLHGYMFOQkkTYWSIEOCvFlGehXNY/KJldAJ4pCZiGFpbRuyuGr5/oBkeHa
Q7NN6hTGAN9842oNgFrmYgVtc0LfMJkRKaowH62qApM5oqibAwnig8FSeegF426K
HGR3JCUppRQAtGYIVBfMTfbDW0eI1VQhd/wSBD49Yh59yXFMtNtSc6sOGQYxYmsu
TroZxs49/9Iy8gNEWWBoWH51XEDesVe/2EO5OZqUhv9p0iUeYpv0xMrFwRw0aF7L
D9/X4xV+qfpEdGXem9IwJfuBU93H2xAijvOhO+gAS0CjKimow7LuyIyHZtIcx6nl
/h78EniZ1bdgyhETUyA4PW0VLenIO+GDRfox/31PfEH2xRpooRqteIX7BqLn7KZB
msN08T5dlYGUPTSCPc+aiXObqptDxrliVVLAokokmIjH6oyyWDYn4eJp5CVdKuCZ
0zWcKZmIepctVILLpGcVcFbMRm056Un92MPzr6QBZsk/ysvdc54HOlANrPzAAmWs
iRi6rU/JHeHGhlRVq1a4TfpX78F8TJ8bllkT1o1a6S/4/f95h4+V5jlxSb8uml3O
qIphHYmmZeDD8qsYLMZBRb3erkhLWqj5/8sRxvf6XEeIDbty+B1OUxP+cuQAyfUT
5sdy0WCJ+coSf2yRq0jCZoDZY/lApgbSqfH1dOfTqJS1ZI6xgdgEGcDazIxt4NFk
zlbfyQs8S3pn6G85CBh2kJKL9Tj6tUaCNBY1JDLlfB0zq/SQ0sPFWsqQcCjbyNWo
XEexVq/Pq9r1xZBPStxSVhXlbi2AuWGSc+Trf+oCl/hX1lSCRmtXckEk5AsdBZd1
j9yAFhe5rC2u0ueOhNPbEXVyAm5Kw8PZi4FT2q4dALoGd5UZ24FZlNlj9iVEhPlZ
nd3/oiOUm0MwOTUoLJ8Vrq60LVmpC6N44RQrhjoXTc3y4YrntI7o5tYy4LVOg2hh
yIW8HV2ItqmTEiBOGvBbFBcUJaURAS5Si8SOdgevVC1gQ11kZPtsPqMdfAn9T3xf
DyPJTU6v0fcf4RMaRTVKB1JM326ZVDaKvKVFdLbGHzQQg40Z5sTk1qk526N+r2Qa
AblB9dDRL5PWHwNDPx5Za2Kx129vdhajQMfCrleHwfuDfiWRODZbd5LohF3+CJsW
PkWOMxSfJixxVPzaFBd5KD0WpghwWg3kkuvY0nn1hOgo6MrTmcS1fN5/bojMmK6j
nx1HDsTV+c9+ZTsJ8lfZwU//jlqdFSftnbbsbbusL8q+j5fgzz/JEvm9OdyH/wm3
gbsb0lC+0kqVLmoOv3gsLjRFumZXqvAIvv6vlsxGtFsTxRFpYBZFhLYQ1FX98FbT
LozSe0af4+Jzvh5Xbhy2+DeVACzc75ARi18aO4W8LgEHdz94x61tGjSQ1A1/BnZk
aTDaSZJzLYoHdZu3uL1Vhr939sdnrbHz2cQmno40/6z4gf0BmLR4MEUrVsRF6iaP
slKyYniLO2HIXK38Z+Rn+3ekPwHysoof+iMkzXBg0RrGx1oAQCG9vzh2DMv/zVdR
gITi4E3+tmYd5db3M22Ypon0QjSC1LFKvxes1/4l7zBtc34udlLnuu8nYv6COdoz
b6SRYseI++HEUu7TiJpHaY2VMX9xZ0P1NlubK4fsrlOtJuqAbXayj5i39/DDzyPc
PLkryS4YnIIpeQFPGCCkHl5X+ocRk4/X5ux8pVSdXWB5B8JLfXO2/XvClgJ9r/dw
pj6T7H/0uUTTJEKsGJKE9OM2zffFappBFl7EZxXe1QNZCwCJM6JRXFdkZJy3nEvF
44UD0woGFndsZJxaEonx16Jr4MfyZ0OuH3cAqzY82TVIJmR71tE96OG7kVGSMBzy
hxlFunzVFjZpSUWUFSvGQC0YsBD1k10scCql6LUcG5upe+FFYo44eKFqYEwtezEH
akXsWcIITSgYpnc7mi1Fay0lqyyXED6xtCDr99imFXbZers2nYYivxBjbhMaXjc2
2t84m40Dvfv8PpvWetioK+xqJdLlMSFSo7d9VdcvSZe8Zys7OLSFvTfh+9Gl9v7M
P0KoL/TTyIE71dylC3qV8QIiB3Wn3Uk/r3+t7Jlvms6YW8VYprhYGrAxNkBy0Cjk
AXA29hdIppjP5HAGf+3z73Ob8mlh6f0txE1DFDnF38ySkx5U9jc3SOURkbtL0ZPv
YxjLurYy7zG8YjqAGFRpTh26JArZJ7xQS64LS7L82Kf3ajg1yVkBUZIJkdtEJWwi
HPCZM6FLCBPTGWxYjtIR8ZqLac1FRyDvkxZkGcXiW7zYKkwkZjOw7bskxi1rL7zS
y33sB7Wz8lhVdXpa3qA38e6YDZPmqFfixU9NN9ogQzi4I6RIN+WDMO2n4bjro8Zm
sUG3CAX0vYfHD5uxCUbooZAnmryw9+c3n65C11fqO9nF9RHbpqfFBWq5lSYVel8W
m78u3r7Ozg2AHNcBpo9cnxHKOLx8HafLl4wp8ipDa0jgwQ/Fyde/TDiM2x+5Kjc3
/Fkh8Y2OiBMsYgxthEYlDTT7/l9HT4LX2vybFbgjpsd0eW31xpsdC4DTroC4W5lk
EndruWVQ20+DDHYdLIcdNLKtsOR4xrC5DQy1E9Mf3om+23cAkCrTaJ+8QGtwVZZs
LAPecz7WC4sKDKtHQcM0h+jBs+/CnPFaLeuvMTXBGBdrVOFTQdWu/33cPUkzpGfx
+5MggwA3lSy2KTx8IarZCYS7dZitlL0Cu1UjQHMdkhSM+ra9YGGeV7vshuX4ejnn
urZ84ChMg6u2sh3QG9Z3/j6l6huAtSBQel6+942iWZyNybs364ZDQFlG3L0REbIk
IJVh2NAV25YfUrFa9oUZfgKNd78kn9q9a5DsD7TIlxvC5HCdvYkwO2Llaelv3kRf
KGFjp/9LuMEvqEhP68CLzvPq4y1lxhO7PALyqHV7TQ9Gs2sseCm/9Wpkcq3N3I+4
tRGZSFfaiRxUs6HzKqj8mgg/hIcE18rqFBOep8OgXG1+ex2AFSVhFVZI+CIwzH6d
mw+RM96SGZy3n1/bQy6A7NIC6yPAKcNd0/rcaSTZYOS0V1dbgMhW0GnY1nPj2Tjv
L4Byi5K/CgS68z5FG2AxYnu/D4YlE0WVnBk/mJBYLgoMAm1ST4Fth9rguMCo1wfh
+a3yFQoSwV22ox7LwgjCOTrphEfI2xhFUue7M1efF1dPnjT2hsXivTyo9LYIGIXm
bygvsMvmcaiWIaJdnUqDVXI1VEoNgTLO56Gtd/c8ZC/n0xqli+pB/+RbrshWRZXW
H+3MIz+wcdtzwKJaAsrAmUSDGnnzTAH8q4zns1Mq6sQCaSSEDLm6XRKeChma9cgF
1sfoZlToILFxB64HpfdKIrmpBxfl0KYE8P4M0nvD3jJxhwvYrmXMiJE0J8aCRhjD
by8YJT/3deS6kDakmrELihLrPykl587kDQZnCax+Kt3LTLQG/2slncHbNViIb940
Mx9P8yGy8j/IUoEfmuypIi8gqEmYbjnF06Zivi+9hl9TDJTQge35RkkbxX5/RdD0
tbPiVMhLxzdSV6dkOIMYCbyz9VXT68PdBGZj6xcTSNBweiwDBAjiipvbQZpbMwNw
i3Id5pvVhx1fOTjE2SR56fz6n5kCIxySYn1fmB+IzVl/5C3aY6aFNorbq8MkDdqT
DH++7IQtYmn8Bc9/A54nFG/K22iv6hGSy4mRbPTzsnhNtSdvqzA/xc71VPYFuwHE
2r3C8L/eZqv2qLrKQYFnEWG7yaQ8VrHNbqjCgBePgFt01UDnh4Cb6ZEfs4u+scmz
ejYzCClwZ9CDLBzBbaMIUwlLyGQZh1D5lfDI0eCAC212/Zzodf4v8oIAfnwTi0XI
PbEMsNL5+2koYZdiZz+6dNllfb+lLKlFYmMm67jX1in2uVroWxvQvPWOMWUKz/jE
bQeO6ZwmWD20jYMVboF/KSUYpWgpJlZ75oEdQRfB7mab/tlKSYGoai/zHg6m95cm
Am7cfyAZrk+rRmzsqQR0MTOERna0LImIKLFXvLoOe9zzoQ9okyZBKYzV6Qx57TA+
cs8z9Cwh/qbvhYlU54f/y4cTc2EJPGe8tn5Jg88ixsUpZhqEP1eOJkH9opeN2bUW
TIg/uOTyivJANKM9l9dhZ5iJogc7ID8DQ8sKTFBkCiyr40kDGJ339fKApLfNjA7+
fCe8EGOPtGmeI89ZmVFRCjdK30DXGKL4ifipYICYOwr1BZxGP4GPc/5ltGREMzn0
Brx1DAwq0PMi3kbPHnE8IKNKjcIt0XvDd7vNI/3mvIIR5VFFZM95PKgEuDSaAtWI
ZfXqXwUAdlV0HnHW5Wi44JhGCpRjv7957sf8ih82lNei/PNLQhyGT14otpZHXP+b
eMlOYoKSvamzfVlZ1x0iBi/kEDQUatqwpB1us+sRQcqFyeSOUzlPfWyLCJ3NDB0t
IO6QvxNqiR2Bx2nIF9bc7IXJYPdvM6TETq2YqqOklra7sFJXHB84SQGfuINd3HwW
Pa8QMfGh9SSZl1sIwSXEIzuRsIOLLjOS3rn+yBdNWIZOvSyztUF/W05hTZ4y0Lkx
miicrzM3SjP9tfw3D1rG3RkxmHuIYa67XT3G+kjPOYJCmNOMCAWk9PqREdV57d1X
ceLaY4mDEWORXy6oUt+/4SPnq2JBqU+X4uPQAr/vDe+EYEzdaEiW9oluO9cZNXU2
xFB9DGE7uU8JBkZfhEHPQY04oPbOxTlMi1QXWikzLY4bQW8jtfXScTBLM/ejsprH
jyQrcfUAjfqWvAYIgdAf7QY7+IksmXiaXUejtGjVXH/TX379DrMCiOMFg1w6k2sL
kdHZyDOjo++n1FKliTsI6ZdEe3fC5RaFpMsXHck3zcJMiaKh5RvkAG1ya3XAdX+T
FVnffXYBmQc/nV3441UBOSe7xydsR0sZK3mDNllXVz/teo9S0mk46VI7lJUjrJRN
enVctjcC0b28QZiHOn60A289C/3IYuPgxd2jf1+KcGAN1XEcmf+Jw9S1EG9vxSGy
aqmNrbrrnRqL0FYBvnsO8SVQGDmw6R5ZA1EhZQZLhFn0pulRiRDQZViCxHLZGk+F
U6A4GXq088KTyR8Bjw3F3kxNx4NEzslg8Aksj3FsRRHq+LAX+xTbmUNpYkAZSml1
6SRXyPt4EecgqCFU8ms4mMEepf97dMxEtstLo5pv5kbDav7CGpMhIekBuYWxDfJa
NHNuDV45IDgF7E9NflHvEMo4AB8RVkIHlhF43WdQLQP2SBzH2qgS86ogvaK7TXD3
6dOl9F71AcPfNu9qM9C3wo9i/S8Mam+oKhMEPK44T5z3ObiqlNVElIBEXA4xn0P+
pUW84zzmOJD1xicw+okzcUJJW5vWsdaV63Hq6W8cPRMbPzeCNwlWRZKfexOllVtq
8EkkU6b4s9rrV//7OL/eqIF48buMzI0EQy7ErqnNuXyNK6kxTQwEfVckgm5kCH+Q
cG8Fxh05RV6ZXnqiyMu+bMSdyjnhsAVqMUaRG7uJOXMfQh19ovgocoiWYRG+dkW0
yEmNq5VU1ShhrgQ8OVIQwruI+G4YNNcbDMofs7soZptzXg4QqZaI96EHIJsNapXV
GGtGGe64rz69GAonMfdtoI79ucTV5N65SE2QCAfReCTVPEnMzE52Bu//RQC5+5/2
BbugeKDMPtzmDBGvPLGf+mGROmhcNrrQ1X/xfHWTNHHMmiVGJNgjWx4k5QBugCsq
L/nIGr6UI/v0+XGIn3BevNIBKBVBGb2hcjXVdItT6yuY4eBAhk+05uHpCwVgPfiN
DNjNoR5al9g5PSsLrI+QcwanLH3TACbZjlt8t5vLr8/NuP3SjQhsFzva7rr2GXy7
0n4Bd5Nr+TWkuOG2mobpuVW4xShNjLGETvXLAOz+8ZiWpgAHTAY3pWSQgrZiSm5o
7ZIy7ovPrJvSfD5MSR/+/hAMKeTirVZZ1QRd9AU6ozt8q0MFwQ9RrgGmLKM+9SkH
WqUsQ3Oz291XXy4Hg9Rk/GyAX2rlO4pPW54Eof+RTmMxOyPAuy9KpS/d/0+vw148
ysmMVphDIHkVrimcijPleVYUA72RxZjs6FC20fq5JU5NwUgnIuql1vxRA0cFWub+
1tqu6MY8CVZzvP/oorUwEUO2mXmMtTbWXHsghDj/u9Q8+4YyaHqBzCR1CLVm9nRx
nvj5dVYo1FQdJ3/cqjkP7FN6DM7Hj4GmiW7g97S4nxjLidhxXvCAltzpIRR11Sss
+IvGwLltujvgjFkkIpLYWrm4u/ZVpn0IAm2LhwIZfelQfxulbP3WHqinSwXxmdC1
XK1XY7TJ2YniLyj6wAzb50XpmjnWdhfsQXcCqrjoptfUZ1TK0Hyiyx4a7kXlUQ2J
b6ZyFDVPfkGuZvpiLqUDPearnn0MBWw0DtBr3WPGc5NvAw0F24e7LXPGxN84WTDS
SK/tzsYwGDKLWAHLweO0lXSXjS7olRJv4RvGMrd26ZsijO3oiDvSsoSCmqB7mjpJ
dzsDusPhw02RrWRkyg3bjMR4qV0uH3y8eoQ6emEnyPXhDiTaRV6LKejPtYwWb1jV
2z+KQKSGM59atkzAn3w80i5RpTJHEUMVgkb7A8b5hr0vQZBIX4NgrfSzXa8AU+oU
5GrVOfBeXo977hba3hoUI1qgnW5O6wPE9mkdRBLtps5KYr7fED3XRso9InuUI7fx
CP257WDbtlZwZVFnaHNMIGNyzwe1gFWJZDmLns1IDnA+4w3vfwXSMXPUYJ5ctVYV
z8mULUmQWRbbgyvtRa0PULCC6FOjJjuXtXloeP5rqUriwwUzWQlaLvv9LpMgFNd9
NeUkG+K+lwvz5pJbHEmtoCT5V1EvnmuRdPdDzojqGuAGOHBKdpjFdZnhYxDu2Wcf
yjnuPmPzKt//RZoEcQyhPBtl/lUvxa/wv5NtqbrxIclowSpy5YhDO9tJ3hW03WBf
ieDIqLCXUsZuUzJmNoFJ6YbirF3KrffOhYD82Oj99Vr7PamWxs8AmMk6F9VXZop7
cYNi9K4l2pOYCFvhMdcu/y7yXwgQGQTSwlFzUkSkQ3RhFE92R8ndRBEvO4zdzHVk
+ispBiTqez+CWaTDqto2y8AjC0SYGVG5PN1dUaE0znN+/mPmEzoq13GfeK9oSE71
3v6kDEZbumRqEdRoTliD1a5ALV4ydo0LymO9c/Jpc5rO8J4pKbz0dDc37mHrBw98
6bBtU3XXz7s0jAMF4jeQi+i9Q1sOdNtpJd4w1bpughzVw84hSfG3JN+hyUTP30Lf
hIyRHw/MHr5Ck/mpw2SWDebuorCyvgQ3Q7MTswAP0DhKRP/u8kq08VuSAvJk5sUL
/ahCAnWrgchTO1MQySXdybJqG7UKXiaDpjjO6wAFMwc08UXU32cGu8MDJayFTIvu
pX4ah4CfxJWVTArq92caczNScaOx9sruKcVF1cyjpTJxUcTZb6fOdH9UOwlJNRC/
7PXC7vjhJwocWyi0Gll3gc/qIWt2Ot/rChguDnSHVhYpkAn38v7YZxYGIEynoRZm
uSAnx9YJMZbYyuD6TRSFktuXIWcfyjin4yMp/k0QSDsakfP3LqNK7ZfyNvv7YCRO
Q7ytIJEYd3faj7lkEs5Bb593TwJUqLz1kek7fNCB7e+pPgcDd4M80R7QcbL2pZrt
o+0yX6DxBHPZKMRRQs/nDOFju3bHVOd0Yql5v+YEflVwg5ZN5v21Kgf2zjmI+3TL
vgSQDx7lUqmGRc0ulQYiHK9ZPs9DcWkZfQey+23le9E7c3rNpz1qCGXGzTHfH/DV
ze6lZwgPurXR3bLtNxSxl/2StURHQ4m91qFJOxbXz399uZ/SbM1tb0ZJSj1QJgc+
0owypV0QbYV8T4+RZj/qfJAWwa8nVrKF5ZkgUfgliZzFNWSb7h4Cz0GXhdkU0UHQ
rO5AKHgW3A5n1/y64E96xTUXh95/jMzWp1qDC8isz1XWOFZDff+ZMxPF1ynMdwL5
dS3BmGFSwKJrajrX+r/BIOiZt66TLoe93ssA2zHMVeWgu3MKuI0ToglaeYUyV26R
OlWslWcsLumnceiMdLg9yEQsB03aGYJlLhtPZOcAPbDNx6TMrNHT+ZvBN1r8jT52
DP8hqT9dzFtzcuUsjyZBqSg9vd0OONo6KvPcrnw2/i3+Xd9phX7KmgwjMuZaD2TO
JdO/eZXsJ0lKspUpFCjpY2DMfJKIMZAQiWPVgmMfqf7oRw2SFuBDNBkEs3WvkqlJ
rIqHE7gMht/O4HAFJdnaie045eQFgG8pdP5C7euu9emiurOyzQju/SxoysEbFVuX
j4m47f8f2WK+rZAd4daINGmEHk/ydhyAhkQvMbz4XjdzRyvgi131LJwTDYdETNy8
LzIdRRkS3wzo/Usxp8WbOZhhF11UWabV9RSfNw3XaDsukZNhdxhxN7toGQtpR8tV
mTkjVfb33VE0+tgriy7znvvHz0z5z8OnZQS4qeVCUQ6WBU179Z5Fv/LtfhYwp/qu
xoK2K8REJRl3HvcnSdZ2tz4pTkaqujBDoqE6RXQAFP4bN9P6V0CGFr/NSfZTir8G
TlwCbbo02UOzhfzruXSqC3gdHJPjsvk/jDwwakTT1Sustsmkw00ysvHCk9EI5toy
vZVUgkBrJ71xwvSugQchgtphFUoOFGHl5uGZQM8Nmh6JQArtaQtJTqPXaNbIV7ph
9Q7u/L+FMbvy5oKqPWMsu0npDUTXJl0rx4GkjLsCMd0PdUxv5qRCHhhUMulpIYut
Dznqh7xpEu7vrZFTjH1xH4qN/DmA7uqjggXpIfoniZNZLcoIzXPNqPHsvyKpSraH
h4RcP17taCPQTjXLgh4nMkmb4NLPGn2ztpZbu+rqgfbxAWCq3O4dhJn3G93hdoj6
WCZNnoWZYB2VCSkhtGVluwmQQr1J5LCTpwUSAGdiuFftZh7WYj8pOhTC4FS5Uh6e
e0Vpq154YaNyLuvnQF82kyGiGMnnoRsoWfe1f27eRUr9dJQQfaUmXgC96UfrZFZd
hOeeALdanaMw9umano5rAhqxVSErZDYfnyiNWVAClBzYu4EMCrb7aVI7ztrludqz
fzQJ41SBRQhaN2k4DAILe3247BvpVdbkBCp2lz/iKB+lR3dUGtEbPprY0s4gPlxU
0spv4iUYVlVMLAVhdpKBD6Yb/p4lM710uDe16qzKNGE9hGhpUYxcNnp02s5xyQ9n
7B5IVQ+CuVjIyUqndKMI+cD/S0WSmxd9qhMGff2F4Vznj086HIPM5Vzydxua6l6w
7327ttS4tSRTMWALMgSyOqW7bsBB5wILBsH+cnpJkbE3hlGqHB9GKe/SVv0HGERf
L4kD4M/3/U96KHkuE/TZ7kqL1HP5jx1ffSl90QxmA6LmucPpe3zKYtuZp3b588DY
l+i3A2qeCz20Cm3wOYeR7DGQXcXc4ywNzh7HlPsvQo4LzRw/xKLiDxUdHoYU24I9
sY1nCBjXPMq69p6VVEczglAPgJ6LpAuDSapaVs+qlUm36s4oqMRkwpod7pfsw9kL
26aR0M1HECCLZ0m4xgHth7k9A3soKfzQrXYYX85Ovhx7RQfMj3vyA7SbC5P3OX2f
`protect end_protected