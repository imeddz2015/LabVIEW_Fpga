`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 14720 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/9huKRhRMtvnNqb3Z+UU7TahEoHV+T8U3P3ufru7l1O
3DlgtZzb9QxCbOjthp9+wDkjygH0eUfDrEl1ovhZG61F9HnOdaJOZTe5kl/x/QuM
doRQpBfq7hBqVvgB9l5JEorUv2W8JwKRmuXZrtAcwoq3+7kpCLgGoQODe8rZbPjG
jY4zLqz1kNvkDxIswWnpT5Ou5Hfc5MuHRSysyC8aCLwToixn9JR5HMhSvuM+fmcz
7BxWECWoGfp9ZY2MXEbJ6qUoPDBZnjw1x0gbuSE92FWbot9MSthLXi/RK0RRai6z
pOyt2ZBY/ICNhsU7O7YhVhFv97Nu+tUn1QETE3gpCd4ViarGTyM8yWp0rRR8ybQE
hXbj4boH+zLsdt2bDdTUPh2aBDSpv7YTbsv6YxSd41lTYokDi4KNgTYnpLZ9kG1d
aJ3iJfT0OHqNszqPhynL8W89Qv0UpwqInBjvAUFMkohR7zkQxvyZXEZqZbezTj2n
IgnBNjmtvEDrT9rbBB+/grTTAlowgQwzxp4uJzdhLz5oi4v+x7YOLUkIx0C8V9KI
wVedwrSSFPSnPIVxrnrOTtCn60RyCsTrToXRLoNdSyhyuBz7JZ8bA4OD8FB6hw3v
Dnvw+j9LfisZVY8dyeGBMGPul71k3Vl+LSY1wHrSoeSv8Z4XMGyeIh7R29TZr12H
FVOwnIj4IfP8myxAmrY/gGnGF6dPqDeeoZZh3QCM6H6bk2yW8y1qPrfd2+K9coY+
vLUXmNjb63zW5Ykm+NW5WDVjHK2Akl8+PSXieGWy43XYIn1tl/xtYwxUZUy3tDp6
pP9LzVW8SGiQWZycCR0dwluIr6u2kUf10xGKW71wKf9H2ts7RRFcS9/vXNK+0N7p
NXmMydoRGJFhlaw1O/xNLn7EiyFofyS5+2TeEUnv5YluMiZCJyfPkCWF5IWDFxND
cTHv+Qt2QoZ3SmAcR1NN/+ObvCMIzsXKjO6K5ivbjTTFjN6mq/LsTcS/TOqzv4Xi
YkG6iUBWgE83S9SUrzDaYX3rcm0lg7k3CyHJUn9uEuGHMKyEcpG1Vggc3XT7Ln1u
0avUjWfQtcf++mthBpBCny6kw1ttKXZU0RGt7DEQ8QBEvok03nyLTH+n4aM7Bi1G
DeG3mC/nOXCzK4Y49xpEfk+thddap7TdCPWEsgLN1hBnXuI7kUWGB6Or7EYK+Kvv
TdaYbGmVPlvax+vnRqiCafQ7p7BLSPRqxiXbTb5rsjesvO2IkzjwCQ+6qQ5N90Fr
x+gFWR7jEwZO2AQVFIQHVyS5esC/BGa9jwQroOVr/HNMAE9Nz8WJhNeXLMjkyHAb
7bBOdWGDmo9MwcPCf4rhchJBXdR0oOV5HwMipSS7AJbZfo7L+WtQnn5xVg7uVr66
5wlVvdxZbWp58y05dynUExkt4QmcoBTRYT8AJbeI/wHytMXpElv60Sn+aQYENNSi
qkf6rSsc2L9fyhBIAz06KE12V/jhV9AFlMP0fuaneHSvoATQpSCmc5Gl96Un5hHy
QZyXLr5vUII3hHFPoxlpPv7Sj/b+YQBxUlEfuuC2vytiDo/jGBO//w+NedpF0ugR
CWatZBVa0E5qTxi/UBRmNeIFvn2kRGrVrnZdUmu0jYhv4dopb16oZUiNltu5EFb/
Sl7QfeBqOUwzl20dYbN3F6Ef5g1X51evl0PGQsVJv3vYVlDjlMysg1hoSJUs0aHt
KBlCPts/zGyOJaoFEFTtYkxdy7q48WozIEkl5+7x33nTKdlXyG9/qee5JtKBjKGY
aMGHrer6M6f6y0rSa4nqyisdzxgr7pt9J1tK0CqkSoA4sywebPvzmrb++fSc/V3t
WozfZm+G7KgaltwoBOk3HTE1XDGirybHUD3kTYIJWzQZdKbp7THq/OBgnJK2n2tp
8ga5lBTG6JlUfBoSpbVgBiFGFVUEz042i0UxhY6r5+rA4x9c9xJDyRcbxTOsgD5K
9moenxlwHno1G5+KnZgjzctonRjHSt/VIb5uzr8kUG/oGa6qirC39OtjIgoLg1T9
u6p/qOPGtsHw8JZKRI7ab9GhEKIMojcnMnV12gkElPzDlMVShkI1sydbk17OMOmV
CTjYWRUjwjm2ybTZusNHFPH6u+vECqn7MHKaZjj8r9fqc0RPKZdjcK7JK4H0v1bE
3BYTWpu3ODLrg1jeGr6SkSYEJr2eY2FsekpG2TqszqjYYeWntaynETXDCLuQRxRB
btLnwQKWPqmHeux9AcViPCY0ABWKVqham6FChtoAMd2AfVKwrt7aKwCqsEjogKpf
qRxbZRx++LAD6HKopG5U8CDneNVuNSr5X/LIv++vzAW62CE8YQV4sk8y1vYFdl7O
luIZjkQtPkzoT1LyMZd4hyZ/M3+rXEff0wUbru7CDr11jrrzEW5Z60sDutkAoxIc
8ETXqSgcvew/bEA7mrZVGLRAksbNQ9T67jXC8TLHKRp1wRKAM7VDKkFnNHUb9n0o
aMIor6lpxg7DKgAcHRyheXS5jSuAmPd17vWEfnLaczNRkqdT3JLexchMv0UAMMis
qCgbIRYKnilUUixYkoKxmrdI2hfhJ3lR+ztVjiioTgGrCdEKttGqp/sN048PG7zp
WpyZWHI4Kjqf87Ggh5zcyQe4FHuazZkjNHk7+fP2TqlKGx2MWlTUaykMlvA4Xg+0
CgMgEd7g8EISncDzLN/KsClQ7NkIrJ+0u0y8cbzSZVznhCADOTTO792veDb78X6I
ika6F65/cJgelhVNYeq1B1msZiHmK0/EDtvc0PRVjsz2flb0uORwppceN2eoJvm4
MlWVoDCiYImY9Mqs/X9Q9hmQ4vnbaDZAW471tSAg7Ji/HAdjwQejsnP/X+MpKr4e
1TrV1S55KG7ZbESvmYLchY0zmS+gIfD4m6glPZEINp0t8DDwQs2yj7SkskkSk0sH
QfTV+l36Sz/0gCVllX/7WtREvqMLFF3frLNDPibbVWQMoB6SGscNyWO2QQ6iYd3e
af+kJsm+vF5AzZPjUGrcmNmNQfaXzT6Yi4kkQF/DYeoWFrCUIHz/gWgl20Q+wb+B
bC9NdV5KtpgIHqRGvM7+hzOCiBnpBOp1vf6n+E+ssGG40kAvZ05x4m+EG58P6M80
v/ExqbmJpE4Er9hgT0MTtgKLsS7Y2wZ/qOtAy1QNvRIRC/+pgXhREccz4zvlN4a+
CZ0f+zwKYk0B6g4/WxVKYHj0VM8RqrMYMjoQWP/A4oJUkPvf4XRZEB8j6vbzNGjV
2FUKnhXbeU6kyUV16nVVWs9f/LpYuYMwV7BNKUVMRyN75suNK8iRap2jf9nZwQjN
soe9VzP3z5BXLIN0o5CrUI6yAxDx+g9xaQwzRSpEs1vBZu/U4Eyay5aTSGAVtKdO
ovdC/2iaRHQk6hwNsB/+yq6Rw2vidIFR5WfVE3LRwcjKTrXzXrlptYubFA3c/aQS
nIqFEbiFZnOJuSOa2g2Feoo3exeEq7NGUF6lGMrpnscVJpoL8gLYHFGFro8LVh2W
Z1+sJYeMhXOGvTNZgGi9HkEWJlE6ELPatN/ZPIQGWA9waVw7nh/JiKYQDm9fwYjc
+vtwvb1+ley9KxEyApyeIhBx6zm4wjwjelyRTy1tA00ZwD/l/1CCLSJNu8NcXly1
UfXBoLiVxYb5XYob5MQgnDcZBgMDhZgJm5YYWES3uBYaun7eJKiPomQx+Wown3Wq
jrcpMyqDIbnGM563i/YOgLKcHMZmi63ULQ45avI6Zfl9ibexSaEiJVNWANjJgGHO
lhkszfx46vszBwlWhU98faDF0PFH62tMtJz0liOuwQB65EZMUnpd5JOiB1jH28E3
phPLJPuJejX48ZnSksI+BbQWETMvuoUZJIsfgxvv4SFef2hpDwVW1JjsYqF/KN/0
eW4Jn7TfcEsuDpSaOdMld/uzN0Q43KKXfL5w9ot97c0UWAcep2i5kUnPI8fIVj6w
ikdszMN0Uf9Q8p1gG7N5ymBhYZaz/NrWZ6WWf8VGiWC0dH6vSLh3pRsh7i+7Ux9R
tMJnmeI8F1pBD/dX+QhUf7R2CME94uipQ+TuVWgHpHYHFvUe3UWQs/pH9MNF22rW
fyJ6sN5Ae1ViLKeHbZPBwUgCipZqDLDznhnObYPYEND0plY0CjyEE+Yb2k+Uglxp
yre/YwOkDOLmKpnM5e0gHF3x1NPgF2Mpq6od3vs6VTXBxNnLb9dS6lz1NRAneCDT
BpVMSRliJNIevp4a22Zv3eB8pg06CGyXpbPxdP3I0CF5LGcMozXA6Q3dxJxsMU86
5l7yBuLTYvLUfIsULw/iKncCcuwMcNSjOTWS4Roc3sJCuHCgVqbr1luDPxcZz230
1pae+HK1TQmUIeQ1dETZT48PeK6UtQ24xVC7isRz06DzPKzAEK7fGsGSSSqMPh2M
KGz0EhO7+CiYePAdXqPjaM7hkupdoxLyE0M7o1HApT7iw6/GLAVJ9sLdLDTtRN83
e4Jy/ZrRkAsjiJcCdrnHoQ1N3g6FcuNLw5ctI4thzyOEsoySZsN4rLsF6gPexwr0
23sZNPeoA0NMDyNt7EfDKYZpdADmWhNRdWCj56Ae4Ak+YsHfen8eDyJ9IMyNZrqV
g8ZFKE7Kkz/PjZdWvUODBPOdVbtVbrq72LJtOhHkyH5EU/Xje+9a4l0FofXIjE3r
bQY3gv6LY0NurX4CeR5BAH+CJnjdf8V0XThFpYnFvhkMJhuw0DgLA/A6fhBCCA2F
ggKFNaPL3Q0b+LlWbrg29fE/WVTJVX1sF08qFR0i6Y7PUTsNy3BLoQ+Ot4z0Sm6R
C7oPeM+v1Wj21cKeidni2SfXgQB/13UxX7gArrqibDYS+PoeZDaDuQSCqttyiOsi
rkEhCRGxFw0THVtHI/MZaEg2T7RjACHXJH4jmIFHRcmxs2uQNxUqlyHoY+3x7soK
cY2tDCw66JLPrQhTcqo0HICX/isz0+FW+QyB5w42vNocOZe9zibnQVPYCtQOnrsC
wuDtPDkRK9BK7sqwojHzcNtvjHrBxJHJqoTRvm1I59mjOpapwKon/hhVSE4y5D9P
aZQhR+VzchHT+BsWoNCr0qPZJFGMJLL/GoqkaDkSp4b7mQ1XO00f2rjZhLJefvaX
wac64x+sqlF/J81WwSghgTI5cQaaMl6Q3zMMbdj4NmGIRsF7nLjrKip4ecoQfMPf
eZvk2ydMeWR4Xa+0VZIqi6JiVHUam3woMWvbwhsfWW11wNidbO8HLu5+SCShlaqY
pSLb3S4bmLRLR036O5XcyyqclWXBSGOaza1iG3zxbfcKH+DsxcwSIUxUZ+aVFshw
7vBaqnNx+US4lwNQ1cxe84CutZD5QMe5S5G7CBdydhZ8UpzPcpnBId5Z8QmoxEX4
cDPTJcfJYITpegvdvX+aG+nfa3maUUt26/TfqENnML+ZAldL453BPNnsF+v1wVm6
qHtERV1J3bArHFjNz/Y+n4HHemz6cGShWxFC2K2DAxnEBh2FSNROWSI9LvIfHOxl
XnyDxs7yAs4+sv8d/YvAmT+IBpZYaJeh5OzmZ/ry3WcYsfWHXJx6l1p7nFX0IE/i
DbmmR4LwI4rkxm3262BUBPgqeufg57jkHR/iZtkvE8HQFVViB+xE78eUdyxIgARI
JReILgG3nwhDlJB4Eh0zB2OLlqTW/xgIHtPe+UHM4zhGTDx1VRmwQvAB4pC4ah3w
j2J0wu+tj6hOx/6pRsZH1O2fq4vd1abCBtIsPd4mbUVbkekXS7pYn2SMpX0Jfcsv
ay/DdmNSEMtv9BJGyCGShMJfHovlDrf4NXXe3ohU8tQSGW0aWQ8WM4o3iCoNx600
AhBPrktp6gmbaJD4l0/OkJ7eJEEbcfWNWtGqeLX86MRgjB4WwF+YZHSGrUFo028Z
1XByTBGd5EhE6IQwWpDq71vWYqWVF73JnebkM0pgbNGwan7qZRl25RlbQiZE3B2j
VQ6bTnH6SEh9rhP9H2/5pXFeLvlerxF7PwilVTC3HXZQ86zFn2w7OxxxAMF/LTId
2FBCN60EMoGyn7jvgw61OniLgsmO6tAZK+w+xdU9sq/TV4H3J2cWbYTyLuA09VoB
PMPnFjjnF45NixlzgPCiK7OtndktUd748CYvzpDVhnp8gCARRBAdr41VNCCcqDrk
91wf0Zo8i4R8ISvIGOpGQQQyrd2Wc9+RmjAb7GkT4UnxV7TaDY2h4lWIymGWKDeC
PD48JSmIem39bfk2an1ZNtMIJL+e+v7nhniP/lPQq4B/yZMhHnJwynFnqaZoWr72
C5s60StRpICrOw97VEcmZf9PkPzyK0/4WNEQOMEvCom7ZW/W5BS/0rKKmhgo9b8W
4nwh8WIcy9euQluWFGUbS7ZGfJuU0PniXWT9qUZvBzSm/8hfb+KGXy5FI95mLqsz
yzijsFWvKxhsEThgv/fwa4Jb9Z8JT3DVVfqSsJc7Wq9Q2liOExPE9QYMoztaX/NY
Y3ImfUT9nu0cCFjLeYuOkf04Yi8z6wzs9B7qXFhw7C2vQfqWesoKCQPlHAnkgcsC
LUSat1WXneWtixihihawtLXU9BwU/cLHdw3vd5st7/LZQqfh5rePmT40DqytvTWN
xMso8fO0bRWu+y0gThOoYpYy+Kt4yTvIx0ib0i0MYXNWfO4euaLpt1QyV1yw7GKZ
fn3ZD4+5Q4X24PdI2kORlzINWS7+p+zfEJH8cThXQi0JCroWVHtYvDWZfczHpvdl
OQFxyoychuGv2kUP6uDOU3v4cfdHiZpvYVNcY+rvKgCNKsnKz/SJPlPYpPYQ30oL
8C85j5EXTd0e5yV7tn1LSA1jtCA/8PQVe9h7PZf7S2LVb3aApd84V9zewQzU+NZR
Gd7dLh0UJYwv2cuNXBDGhAmzd9PoPsP2BVLO/BgolzvhO6zpHPyCQSfeGq80c7fh
5yBJp6oYHCO02TB6vir4Fqv+msDRlKQdysbKMne8UO+I0ziJgIZjkbstpzBm+UNs
Hd/wsBuFolu5qf3Irsdd/FqTEAvvtraFKsbK56soKIKx3UT0ASKEzgrsKn/BDik7
PNn2nuXHX2hL77X/rr0pkpsMl11ov2H7JM3ypnCjQOUygHrkDjtvoFQQjhoiinEk
1nd8fCHIviM4rLZPh4Y8qLeW3Ear/JaymLuFMTS5YpQsObVgdhI/korG3banVIci
zu4/+FyIOPmmdjA5w2sQN/97l9q+k5I5/74b0a8imRl5IkOQc+Uc1SDe1ez6vizy
xpQjNkw7ksxqt4ip9+8gWqgeqev6LDRbMeIvw6CAPESSlqawbZAQuF7scvB+ortZ
bj4lYSdIx06x0jektAykP/Z4mHSk7iWXEM2uSZIWy7X5Gv9obct74+G7d8v7i2ou
Oedi2l4fBMvKVYJMf5xka+IjeCTCP/opFvXNtww+4p1JlwWlYk9qV6s9vwob8fuw
ol7sTkVAJ8J/yi2FVBy/TYv4bcWVlprIs/DTd+zrDbd1V3PeqH6kqISEzxehy7Fj
hMAKdoRelD0vk8i0/jiSASKb60UAPgNR83lJmLS25tc7vXQ4NXzkJtU9zH63icdv
78JiESAX1EuBJbPpmHLOnYDoBBDMwD7sz89n7D9KUFJ6xd+T086BdLjlHPMF7yJd
rmrvfCIQNh05JiwT8fhsukWBwz67PSohLmZOaylAYx8eJN/lfsigtsJHCPsIa+Ko
kt4GC4rzEXqupQ/joZFAhdscsozctEhMNTEu6tn+wIuWBEPaQ6NcpjU+bor5HyM1
lF0CFPE4eJ3Rv0EpiGNft4cjLbMo2UdFvQGJk+yLVQ8ddL1qKXJfVvrHfNqlWl5+
8HQDVEzUiBsGsFOgUsVSE65QjBtg3NWl3saM+m9cI3M5z9tR7bsB+TB21bsXcCVj
HRUvxUyVofwJian2snG3pSETRlOl0qJItX46+qv5/mC5jlXiaw76S2psHAO68n1H
JdVlEWx0CLMgG4AtUNaUTRHYIFIoh3lAYngZFoCGY6iyWuUyNyAS8a1oUqf12C0j
eoJvnnxAyBoNnlbx5sQMsrovVw7XW0/o3EGOxNv5XdhXufDWkH6bnwc86CbNS1MN
J51wqevzlSwYodSBWnx0dPODAOgHgdOOmC2Xt5DaTRbWTAa+d5G04Z8FDHlkJ8Ac
XU7YTIlQ2jwjXK6mmRgwdjTF0SBe/7vOqs9SGQd7Rw0IQ4j3cRlcvt1SnVaPqEqr
5iMdHEdcDnZyNfPx1bmWQHQU/zn1zAZLPeTEcIk3hrBMzx1oVq0hJFCJUKplmvEU
k8wJWSQ49PXI0MU2tl+0KwwKOk2UEji7sbEJ7dbD4fPt14QDAmZDuHkxcxIj5ii4
pBtgHbG00kS8vpSdxoJrJ6RHn/FdcmbAqSqQbZhO8j7i4AbnPZTjloIbO1HI/ZZb
zorQTpKpbY+ae6IF775yfgbkU0Pl5RwUkt20aIu491KAxFa05snBqVelxIvYJ4s9
T5tk+8SM2B0O540uQNgZgEJdxhEtuSj2+UFn+/I9k+VFenOUOWtGWgYZvvryEkAc
ImIMP1baQN9TBkocp8u0tbgrxteM1i3Eb4Zh3Oz4t14WR8AU+AOIHoALt/lHeTZQ
rpHEPK92peax+VIUvqOFSZyN+yBVK2f7lRAqjOgPSC8PSfFUoI4JaPm3QRwtC4ar
QDcOxZalvS55zIILFrEoWbh4yAZNT7RjpCNbPKCT9GIdLpt2hEdC5KwyKsayjO0F
L53NetWdNgqIQanEPTQ94q3Ka5VnfT4nm4RpN/v9At/Juds5ZmYCheouhuXdJGGk
Y8FcQSmpvL9BOZzo4UGh90GkPEgKTMqRBwX5Gjefu8LqxiWcx1640bNHiMReOmeN
oldEZoL2dFvjos6u//3GdRE0aYkN0I7svzD02081Qb68WfmbmvXoNU+EZhnu4m2t
n3dazsYGET0SOfqaZj8GXzuhm2MveYq84Fp1N50/tKYvD5PME1ov1kUfyAWH8Vey
2HlqiNHq2HhOtbS5Z0Ljyx4n/5a+N8ZXK4s+TfnQhyco8SOQWMv4jFa6pLYtIyg1
1WRjppXQ+LqfbV8RRFr6/8w4henGWHeCUFz+a5CuOuYOnrf+cdSZ3PTibV52Piao
znPnRUQ3lHvuLN/79z2JULbIUFFFUy5YLwiKu1TdEA+15aM99SwLWy1YsQ6U/ErB
fd8+hTzFcKTsDhuczhFyvqH5a36EOx3IUffeI2inozhkEihsYkmHu97Xfx5g0z3K
G8+KY92GAhW+rf7ElFvSAOqsdaBxm4VDfWyne+ahnkdJY3JNA1jPEFzTti/VLp2Y
Pd4ZH5ckm8edtfqYxeaI3di1x1cRuSFdGNe+a+6zKQOdHhnZAnNFmkNDJ9L23YqP
/RmdTMj3XQX2xXEp9SCcY1NOlq3MVKtjmxPQPQ3m+HJPyiSfS1scJ/h33RgJNsx7
H3olob/d3/+gxObs12KlMCOOJ22FfolaGiVDa84eHKxIo6T8D/BJhJISrWLOLU58
J47mCWwpN2j8/ULl9Y5JHu81lDG2E67bgGeScb0yyu2odTZOr+Pe0AaQNp6jzF8m
IuDKxF+qiY2rtzGy3maFPJqlrUbbfzxOj0w4ZlZU9pYF1ZyaJfpUuq/PaTIlpzqC
zhuqYAhcvdGUINBGJLnLkFiB0/p1NhPdRVrTruRS3+MqGB+ykF7ItXEz66wKJpeH
Jrn5r2CD0B/ieEHVZ3D7R1dP0c65dO2un/Sw09NTCIG1XlBgEtPjXQiglSJnySnV
kWR3VfAKpXK2TQxy6YG6IOxx1QbVP3mbvJWkCBS77SWcslggsdepxBZWzAqFgMyw
zz9kN/E6p80A0Rqz7SZYQoz4utdOuvyFBdrMj2PlQblgAOewrXJKhnynkLrg86wY
8hGfnhxrBInoeUL/ZjYC/vSvjLYclmC6lghGyVvYK6pYmq6m5ZMYfnUi67uU/AVW
eRxD/T6o/hXS2KZkhgGFPP2U0AYQXGOQh4HGrkfy1ov3h7ab7KEKiE1LfTUsSe+n
kHhKwPq6esCxI748I+QGh3vymYFn0e55nlMxzGVpvb+xO2iz1UKbFqbh2RhDBe1I
IH4TV91afnwVacmYDkXIeAk3sLxM2E2PHteyRwMKO+liEkj6ed/eO6xibqESqCVp
CQohnhgKKVLt7pkenp8M3I2ZrYdp6oiGNudQONESCHjpz3hOIMyyhSOPHTouHBH/
2UBLJ8cfoT84XkXwFwJ9l+QdTSJBtIw48W6qvnhJgzzP8W1KjhSIM93hXZtkiU7P
47ZQTwxD9lBPRumdfXL/hjaEBXYV9PUhDUgzPUW8zgvwtLF79Sg3nR45HZ6zdzN3
L1iORPjg9jxvdgqZhKr6Cgk80NB64K6yPVYOUtmKVwaXrGmrtIuGQOa59bH3JG+Q
9mbqgYdDsONzlaLJryoA4jUSDyIaHY7SHal3ThIwRsPsxc9sU4/jFsPnGO+wR/C4
zhaHAWTL3G3Ff8cwFAUcldvkp05od6eWkI8zAg4tHkSLvdF0QWY0hkZtPjAN8Njg
BuDUrD6CHPmYssFy/5OyZb2hVvReX22682zaLcFeOuVkiT3tPCSe0vtUa2vAtRc8
Fscx6JM1UJJOAcfwq0nbjd1hiLpw8IsQitTL70G0mayciKwYpX9spNCaYcVdV4s/
bvSsMGh6xuIP8AmMqQYw+DjhZu6Fevpr2bqBS7LX9It3ZlX7ySAxaw6FVO3iXd3+
U6zHDXZGT77aghHWiqF7IkV10wsHRQ7Xj+Cr56HJbBDOduej9Si5cWEUllV0vZTS
CCSBRju5H2uBYLi5CGTm0dzNjYVFmww+tGIVX+4U+ymC+g9WySVTOHKkpUkZOqWs
a9jWZNxMt/OYeklg13bkhdhq0BtR7kTuP7GK7bfcgWpkofZ3AKf7duEifWoPmhDd
4OwgffuA3CJZM59kRwvQU45pTzSW1jiUv8m8mpuxCj4v2HmCeesG7FfAK+TgPJ3C
cnZiZD9rD0z0G8VaPyf/9h9O2zs4uYTdeG3e2VZAfk28Q8dZlMCkQK4G4cPTSORD
e8p8MjuL0VfMwN1WVaHkLY0ywXjeFJiajp4aEeim0amSc3owBJGtEKCgN8CPcwCK
mDs+dzw0INwpXKEnvrZiSEyYc2nbfYMwAYS5G+Z2/rC1nJJQBVdXoKQgmouFM+6S
SwNASGrwBNamtYq01wUDcZq3rBdwvv56yZrcHD0KMP6IPAP2mWjKLFY5NVhYo1Yt
w1y3Wns7Dx6hKVrVXuG4R0LTMjBmqtwW3FFEmLcJN8KlIdndhtWJMnP2eyHCAbIu
dQ/gzCVSzjsnt+oqs9Hv1gJRTgbbQ/4Ptk/VsVh5NK5gNwbzXl5VVP8r4veKIX8t
uL6qIITh7z3v/hIRcUokXLRxmywXsq+GXaQ75L/XWU1czqLcMMq39e1HJO393Xhm
/w+ii/f6RgGLd9j/BLD0Zu2vlzbpdwIP5cefpL88PUupQOw5XJ8DU2iALBDge70b
sfGGNordYFcm32HorDSZuVTPW1HYS13h9Gr5Tz/cAWPvQqC5RD59jdpqF47SQP+7
kHvJ5p7/zNzj6X5F99ynVBd6XsHIZ/jPbddwXGwL5DpLW+P27pBSCQ8JIs7OvsRK
HvI9nWc7Ep7d6ngAnJyrUr1QZ6yFvk9MiLW4jXiUxQXuXBD0rrJXm5ZQ/D4/ZmWN
xROR7276YqVhQXOoepmFzdRa0pFgES3/LXeM3WpzXad8ygqg3H/SfLBu2Svk4yQq
ZuxNdiPb8j+l7wmlo2yMiaX97JAvLaVZv0Fj3MicvAfslEX8GWCFQzb7y+ENuldf
wGFMsjd8/oOItROa7cRkzGqzQSL1qaeJu5KYqQV0JLNMlYX6Gq5lOhoQ8uiiBuJH
Yr+wKz4ZoopBVuHuymIsCFhIJ90GPnrVjUxtRxIRN2NjWXPnkXsRRz+wstZLNI4O
fTkCizFlJIgfwf8WfvwgprUQFfOUw7rPE8sdf35YafULvxoZjlRx3NAjuTgING8c
poM1rHvE6WEV8L4mIKuE9ufXNQ22zkR84+uxuWE34yRCfX9TFuXpbVenkxcsfUvC
r2ZyzLBUIxVnNqyvQ6+BU0SLp2/AiAdfftEIC7n7IgvqIb5KkN7R7qTLlRh0kZd5
s3BlGl6OprXXybspEsD9dzEoYvGl3P8i5WDZbbwC0DlhK7tJcaoVbQJCQjYhEu1c
mG3CR/ExdCz1/uyyPjnInS1TMWJ1rfj2x2bFxdVnHwrlosfnYU/ZLHLLGRRemFvS
mV2sHB4PD0NJaYXtMzsZXyAaQzm9vYydjA1V4TWE/Z+LgKBpeqm7Z4nGgV3gKELN
F2Wki5FlTBdosor2jQMytnq8kF18Ak/L+efdmgriQr+ETC2qYyduuMj1FwqzjmfU
vN1tgo3Ts2TtPEJuCBHJsVIwJRc0h/ryAIdxix23Oowi6VKfABxwd8hfTqK/TKfF
3I3Js5TfsKunLJr6JSWcNVPoRwdkVnoIUvFbsvPTYq58k0bAgFmdOKh3Kc8uXvdK
Wt061UuX5dCzs3O21CXy9U031VGqLlwRuuuAZGvvk8E50hlqf515hmQZy68OBtrF
VB4ZZ7fW1+3iBdRtCKHjPQH9IlNfDXigS+Oy5ATLvAO/kqZaWc2PxPvdtsYxiMYc
rtllX77GQOGCFVYgDPJhXVoE+39BbnYW7mQC5gHQAKyexIlPs1+2TZOR2Uqe4rsZ
MG8xTq8Or9lgHI/DxrbrdZZNPuduy9gZr4Pnrh4819q4k7czgCfRwubaWw4qTiGi
rU356mZ1xX9DjDtz8d5p+Tb2D0hpcsNUdb5Pa6i3rgZyJNApDRpgaCCUFoizfIPE
lHdqTpKxqYgirh4fmBuEsnZYb3gbt2dRuRKVMLRMmxc7UVBAMC4IDimNg0wRVXFT
P9IXFYPcaHm5tEYXBccOwVBjtQoOH+AX4540/1JFGX1ddrt1Usk2Ug6ISo1V+J1q
aID2tURZCMQsUwdbEOe9JaM2dSU/UUDFstYNYUHDyoUNJxyJ0O/RGEpcIkQTAQYR
W7sYsP4s7wnBSUvKdpz8oUb4RnmfvIs2Ftbyo7fh4EvOP4Yy70IOxe8XfjqhV+bL
pKvgdfCSqhA+qOtP+Qa6bjRgbI2UJAomP0WOuO8JYFsCVX5z1IRGbardnDE9Z+K+
kPauhGYzP3KWfW62ivmcK+v3Y4NGJJv7q4S1ygV+yf/WgMwlKmcX5XMpHoUiHo10
CMrni4mNLx1M13v/3yzajOW3OZEirGlJZtgmTx7o1NMMK42x+FrmfKyjP0nSBupa
13bmHAUHY3G19R8F1JkSmgjfFRDfBr1DJcNGYfs5EU1tcBEtqMe4YJHZW7jSR2se
Cjr84zxY+yY5sC4n9t1Ne7j0xEYX+PFe44mVHN4nMjlTvu/+ox3Tc5dhS9NqTwZB
ywWwzO5Aqfd/p4rqPFK/JTbEEQdNu3qnaD/vYj3OsoIVMlsp7PK3tCP2gpZQG75h
Tgpw4xHo7aZTOxwHvuEIOrSqDyB6VBVzj/6ddN8xj3sMcyv6DqzlYwJHwDejSyFU
JgIUYhWSMKF1oeoxc3PqpTePnCFDm5gfL+bvWJZGDmoN7ZtRN++mPObKFuJvufXB
LHmOUgnq+a08UAkNgd8XRz2N4GkaFgGjiepm+5UcqBy6SXayMvSRGigjvtJsfFNu
Th/MMok1U1mz2Ug5wCLvn4DYwxZKVC7+GH4H4C6n9offjgMAkvUixqIfsO3q8G1w
KhrMUh3LUk8owBNx/Z2yMVrwFrJAxiEGt8KNVR6uf8wzsAw8SUbHpr3rz4ElReF4
TDuRDUDrbQs09wuHAY3PFztusUfdwfSAm5Gv2p2yyqsndzLMvIBrLMMuV/ekAuHY
mYsZ8uAw9fVVhfCKcyxOi3ju4twHxGHIAn8LP7o4meqvlOpoAYva40+m/KQpMmSf
w+zOPvV2LNTpecey4dIMzZhsLDIpiZi+4hOE+DjPsilsuJDE9FsIOJgh6NJ0V/WC
qj1hizeVOztgWGWwoZRXIeCc2QnqMrgCMd8+0HhEyd3kLAeYpJ0+yeBpVf9iCw4F
UZ4osjFS8IfSv4Jk31SFdokKv+8iRZkG4v6H+oNREX0QGn3tMg7ax5BA4QNkCPkc
mv1/EKpdSYMsoF6aaosOfl0Q4UdrZSQfYxZPoR+fkVEfgVpiLSjIgLrbCLo41n28
vDVaUxKke6IiwKEHriaQD/ecQhA3NHR+YJcpGqO9h7gdmOOv65cydfcakEAhXZ3X
ECfCWYaq58q/ZkJiwDjiNt8AW7+tqcvhJCqHKgsHdAp8jAt6cQo++qdR4rYvPHwH
Jsyf3lXRrL/RDQROjeHBsTODeBYFx+8wRkC9ihsk+AuPjLv89GhmOgt1rpZ+mN0U
1fyR9PZebyRTL3Wj2KwUubeVIkc65Y5EJ8eeiZgBXzOrWOEyfiqdmHxb2AbUSd+/
qQ+d4/9gLm6Eo61qUNpM/B/AlDA9UvqIUeqxczOv7Uxvouypk8JCU95O6BimY40q
jvgXL8liWTH+gAJgAlDSWPUke0D19zoAYWFHJeccS5DyoGOYJURSs5xK0yI+7fn+
7A40tsUKrOmcYyjJ9nxSVOLE4LmDLpFCinJfElOMF14uD8bDz/skGK6Y2FQ2FmaE
VpfG9KenBc+r8zm8JoKR7vmd4tRG78grfuXrd23XXTVaquGOGEKIXEgD0Iy2jWMe
oXO7SfUWpHdLjq2JvpYB4Eo69r9hdKR7P1faNqOR59cgTbnAxlM0pzkZkOoQ/bPk
s9SOhMv2Y2fY9lX6wh03ojtoETviowcIQnrM3Pgu+/OfR1wHkWyzpX8Jy0YJSMTJ
X1AAdkKA2q4sBMhe7VZgFc5PpPvIf20GCMo/qFm9qGRGY3lU2efRX9h/GNakauAd
vnPktPeFMd2KszILYIxbjcThBMVCwwzwpkPrJKQEMp/B0GXfTLb/640IvQVhHhMP
mtD1Q9RcOcelJVjhmEF0tqMbEBF7O4rUSQWoJjjQMLNNSGhtOhtHsdCBCDwil7j6
jCwq1k2KC2mkOfdyWMZCamkzoaRlVrickURyVl2Ft/g8BYKSPtJDwF3Gc74EyrR/
yt4q6Rsifys/i1pQ066GvSJGjL+wohfxvwjPgZSDRbul2e4Tve/LOy04qA0wxf4C
gSWqJHsg+hHW2eOX6irxI9+wHqh3G934ypblxo5YBJzHFGEau1zMJPenbsE52HKQ
/vpmXx+7RhHwYl1CeHNhw6CRaCDPA/zDroNozujpq5HkUnuNiFSXi33YB18Hey2t
LTcszc0LJT3WCrfH/f2kNHztt5Wm4z8CxA6ElTNlM6NWkd7ZHsZY/g3F9b7k6iOu
6hKIlgvi+yTXLElPpmpqMJqAXEpTpJSXMD89dfc5vQUaFPM9Q+aWzUg4V2DS7OoM
fdAO0VBQlzaBpOdxjd4jz1LkCfWMrW15Z3qzMCiVUF4QKsJzYoFRYzXcE0zZ8Q0Z
ajuRRokanM53SkdOv8rKagVu95MnRZaBfl/vrFLOH+Kq1/k2ObrOwbVP95R26P40
QziB71IMQM1Ndh1HlyHNa5S5YFARsgX5/L93sdibjU/NHW4HnKwLZ+b/pJ6Yybmd
ub3y1gEjb/b9Ab+179kMIbJO7S2KttqI8DP9HiQ0l865iEDxKW0CcPI89rYDzuEa
z2ZUwp8gONIxJf4QAAmIdH1x9qO2K9EGfPEJMb3ls3D8Pyl/9ocCbZZErzxL3VQ3
WIyaIFUIObvqifaVLNLMbEboa9yT8VqtJEG+NGLqkcprublTWm5tofkhkbT9xAyA
/XgRU989D18w1nesF5LJ3C2VHpZgwQp/T+tLlXDUZVAKtnifQCBh/w6I6xJh2cP2
g6SUAonYIu4/zOevHMcTWFVCmI+fiqvF69gAGy8DS7IchoBZPn/yQDBlT7KKJTap
5bLvv/fZ/AYeentn7MPgewwVXR1V7LXA5CBwm5QJzKjWdjz4Tiy7YiZeG5Y65ZLx
bem7Qu/W4HOvQJ/FkwAxn0YTVr8Chm6r8BfEqllsZhdNb+5EsWdlXpXcrNRhU+X3
F67pqzYrF2vSScYjqFA/F1FOJl2sJ5i4uqu9OsZWAQ5QJ9VChPfXKNzBKcn3U802
ApIbyCb5Z+JThKMBmHqGe3hftQiSu9wZhrCyIAx8Xswxy7fna69yQOj3HHAJ3yqm
2si34q3PSzHIqdoTtDR36ewnxUiTTFRSaCxEZE2dACzPdzttuKV4H013YV5P6OYT
EZFClDBPnEuoCnHOw4eedlojlxGqXsBqNROouopfVv+qYBmnUQlknNEUItNn0535
SmSRk6fanVVy8Q6CD7mEkcACgz5Y3uKcAyKuVOuOp7kBhPRl/pXaVG/XGR6RUzqv
Y9eIHFGfeO67hJmzZ/ePLW8pL1f7/b+g1xtN73KJEdOEesOFYq5uvPnxA9ioVBbm
yqyBaDpUFDmJM66lzRivcU2Pr3RmocHOV9eziMyaLq6/4g4cvzk5hVCrxX9GY0zh
1J5TE5aEiMr28/CM9wBMEUg/4taaSw0lkyQKrFErxM0yiCsHlpp28aCk+TJ/nre7
QDstGzP7uBqpDOg2it2fW0xfNWGasXQcqZILphvF0niEMAdB/mdxDuM+hTFGtnWs
j4vJZuHHl35/28NcPyWJHAud1sCd08xTC/zR0zNUI9e5w3ByITYg/scFIU/K5u4A
/08cQsPoppEIMONZL7xTioxpUItQRGHETz3mp9uNsRYVLDIteptD2jj763IO/HEX
Qe4rDCQTBFzyPAqm2S6flAEUb5hGwS+Bj02ksIBosQC9N4ZQOb0sWOt469AlcQN7
rc3B29RuxES4wqWFcU3vYlUsc4B8GIh6Qfz9JcZwiNlAmgq2Ay3yi10Snz332d5J
T141IDWqKVE3V5a4TBE5n7Jy6CSm6LCTfwc40SRC7TvoiukfVCLkXugqLgBoSo6J
+UtW8RPOAA/dtqQ4SG170/h1rJZsyayDEPD01aj3BoT6VgdBuo4hncbxh25IFImt
+HCqPWwPyxBCmUfyC+FCftwLsw+Fq6zI/Qynx4rXrD3NT2anKlYmzOHaKN2Z0x/f
g408Xfl7zF4b0pAHhIrrnp/wer9EDyoUNvKAvEPorkAsg+rFS5kTsVuX4vJuhqWa
lVIUaHBtr0YyKi38xVhehqU98XysgTrq19z54IslOl+I8l3xYF4PrXsu5N/L18iS
q9dq74PnGqWhx1+hUmYc3D+eyPI/MmjMwoqVLWx+YuiGxZ+DH3wqz+o7CIinnaGj
PltOTPXP9lE7ZgT3vjJjq2xfUfadsYyAwzyJSrXZCCnfb+MCIGXEMwVFFwhnwNpm
20BGUB3OOOj9eI0FFQnebqX/QGfKWS09no1NfKBvobRHFlqXELd+g1ab5KciOc3U
OxrcvissbNLJnZ+ht81O+Yfm/w1DTvJO+pR3N6UzhgmKtrlyNP0b6dqLtxmzCuig
cqToPh5duf/3VyUDvNfbK9b5Byc8st/TRGw8XLIedkCv62cFTvIfGMxCFaZxx9kT
xInnsMuwBkmc2zk7E6Z2HOlnmBeh+3H0zAhyittSj9GqX1/t+KFd6iBhCgUnGosb
KtGaiC6vb/d47GFoAFjPyWdQtRtFiAE1iU47MOkgA+1m75seFrq6YOiHMWoGE3UL
j0OT0A0/686X0HLPDn2aa9D5BMoZyQPvDDga834Z7dgcKi2sod51FFKMUZ3QJeW2
jgahS1KB/wD88H9ZWsYGeehmJf6Wev3N4XlrbjWaz0lDL9mZthdbuwUbs5IVDPMU
Q4FReDiG0fC3mvRWxBH+M4G3Htz2WMeGm6Gqetgwbd8X2rcSIjWFOUy86fxVMqh9
VhWqWZNdo3rucGX6ICf0ekW6j7bvuG5NoedHO+kB7yp5F70+O7FxbUgEDgnwhwqj
U1uFKx/MlNyR08vOIMyp3VjED2X1UHThPIYue7HSBoyiHekL0x0mYNOEzmZT+Mua
8JSDTwLrzxFLTP1ADBbdmBOvpoR7mSyCLxZJX0O/dka0FmicZlwpc772Ul7D5xAE
iEyvwHlB/hJqDT63eJoejeXWpcxFLx22TKdWPLzbVavSd9e4OCIq/MiChuJB0wHi
0nLu5wzEmii03/c95s/vnPnKZ+XpeChIvVw7/rlYiDFv2lH92QO9sGyXe7K0HXZc
3Au6tw2V4S6WzaahgoUkqf8l+5twOdESBLuXsLPPZernhJLGNR69mFq5hMIafZQn
5HotZgD253VzuBL2UaTSayXKiyFlB9/mD3VnVJaRajqS5WUOKGvPYLZ5lO8vrxHJ
enfQfZukdvVA9OscpC4oo4mKWJv9oBTnBoSx+UuoTwQ1MEMndAhYpPSk+FoE/CxE
B+Isz7pm1oDmzl/1uQLj4/V5JqwJ/b3DYJtMBVIj9FlbnVoSkPMtbqEUX7q+4D14
HOAi+ILF2Q+QuBG4rZHnHJMGg/CRs6+Dn7l85MfPUN2ITL3U1CGcATgo5OnzSxry
DJvNenqwZztAPh5B/veS7oYmRJ/2rDy/Ey09BneJ44BctXfKlr/JXyN4/zlnoEQt
Z2RMgnpP5yBusd9GuBBh82jAxiQ/XunG3nuW8HQIpaubIpfHP4gY/jhY8sKfvNDJ
3Jk1qvOCjZmPWlSYqS/figjiHk2FBpElUXbLuw7Fxi7I92zu62zpvRDw9kKV2TPD
VowEKisCFDVnVWafzrqlBCEJP79SZE7aOdkiqNMAZ8+dMvTftJipuxcwfqsdOE67
CC+H9J8rugcRGwtpEZyZiudLf9XdOXrfNdZQKWSBKR6JczYVoLdiagD/DwgK5cQS
Rmoh0ikdVk40mViAyaK6eMWEKQ5A3o7XXaGNZwsDyhWfMsVVjGQQjB5QVH2kSaoo
MVeIpwO447N3MzZQvpIYDEWmEE1FhK68lmF+ChVHUf+osBsruQC6IfH8pxVCGTFk
S4jdKYZHbHlDPEvAGUuN29GHpQnvonGHcO640DipJslw2/eLW8Zim6vJgzoFqgUz
lK4l3riQlBKpoXH+NEghTUoxevN6u2gNxaESxlcY5O/5U8ms+tbMjCpSn9+TgU0H
EakcdRjbLr+0iQYpRm27umHavBtMiJci7WyfLOqc/hcQREmeTsfYDP0qcytxXjpH
No93gyBi7Pe/n6FmsmUFrFQchh5AXrVDNLc5INHyunz6c9pvejDTXiQsWdougTwf
gRtxEGUPZG8CSZCMOlb8mbhSgpq4eufXk+Gf7vM9FIUjsQcC6jSxN+aLQL+DqYJ0
ONXu6p+DtJzw8YTduIymXLZFksvXKp6OEdmt6qL5vKV5pzp+p+nWhc89fvs02G2k
MrlkxZi/DiCyjaX/9MN/dL/XaCsFlgIj390bXdw+SmttSahOOUBMdEWJzUOzFAlH
GScrv9NOO5AHK9BaTqPlwubk3UNc7D8Zt/BNDGDl4Lv7eEZFQ8MTHkTwIts5uLvw
tieo6wTS/ADCASBXh3f/MET3g8kLijJ19uIcUCHAt7I4SVmrZAHySSB9jA5Ja+cn
MiGTWssA/I/uSl/Q5PMH02ruqm9lmLqJ0mrt3hKsGbkyFiXMpCQgXqEeiTtOIFU1
hHLdWMk/oAxXv121FSTua5jyx2Exd0sLZcuCGZtTJTR1uqBa7WrgbR6SW34m/tv7
Ax3IKI7RkiVKm/zgzFlrvZmkdWHSY8sW4UrYB8U/tHE=
`protect end_protected