`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 16192 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/9huKRhRMtvnNqb3Z+UU7TahEoHV+T8U3P3ufru7l1O
3DlgtZzb9QxCbOjthp9+wDkjygH0eUfDrEl1ovhZG63gA2VNTWdQMGi7u4+JVXKP
ZbuocRpqqJ+F3SMjJwyCkaZTt9WxRKUWlWbepyVggX9JpxVxcAuJ9PKX4gBzsFfw
GzHqQmDlIk2QXN8FoArHZnWz+vFPdlM/MapuzHC3ZkYs7Sld3Aiv6lgkRePFBFmh
wPkRS3sls0Y5nB6dCilujK+w+CQ638lpfdPA5okv30m4F3Gcwhr86A1/H6WK8w13
cINB56HH2CCIOV8JyhUEwrYdjnA913rPLwRFCjTHbZ0W1jt4WtMZdUeKfoz8nTmn
WLb9i8qOm6qn0iCgL80R7s/Qe5WX7Qt82OpAIZ1OpgxtQCVqMNAV2Du7VbK9G8o0
tDYDIkqRVr2s+YDNkLWnh4paDV1JDLuXOpg7G+ruoo3bIgHiVba3EWfuHGjzRytV
7uL2my+koMjlS3V3WNgRpMNGQvsIJJwXvNCCFT/bEueK3Ia8DYIQ02znBwM60FPh
3EYD741Ds+aTRUYTRfJuGfToQCJUR6lMdKXBAMSDDdBuFoDEANVcOBs25oqcX7s1
huxmve26VBLRRAfRRk+lxNaFUlcB4j3Qht5urf+woE2pj7fBeDLfw3TNbqMzmNb3
X8Ik3Zpy8yONw3Tezp/+84Zsfn7hdoyaC74iJ+ooyZwDnrVVjgFR6m16ovxZ6N5M
MO+E4jl8ZH3tvXQ1QI/CEgKjDLmsjYPKyya0VpruRaVYsx49pVuUXBj+jc26IN7q
AFQL00Sjr13vl9W0K4bqRAm8CKPmA0p6e8QYlHL64Pm9IQDKsVIAmUrumMf7Vx3k
/pQe1T/ETvx8LkFFq6+Hfj1o21HiRI15rvTVML8WY6CVYCpxCdAwv50FXVtN0X6I
67khY+AN2/yCc/AtBHbIjTwwKRUTzshKWkFgyk/psYRzEalbwTgTSkySj1YuQQxz
JoryEHgZB6tILKiyN1QSU4v/aVh1Lp6ERNe0d3G/qAMChRWT3+3BfAk6A59rTm/2
uXo4V4zjWKX0VRZUCcI2R6RDpVqnZ8GYda158zE+H7wogym46841/B8hR6N5Z2WG
wOjnIrbRoqS4GK/rMZ6e9tlG9drrxrarYDwDzKGlIpsvOLnjBbX4xUHckmQxv08W
w5hyGg81W1Q8zbqhslq9H8o6UAf2ExC2/fbXuufKQfaRT/rlRDrlmKeywcfkMlqJ
8pXqchy5yvUS2lHAzTJWJe3hPssZIi1e1ZCyhuktm4VxXFXYe8B19e8qdRwCGn2F
T6YVc9TynETbEUMv+nh117AOVOV5B4lQTikSLh4PQ2eZur8bgopH9eA/pbwTe9Da
CKPnB4kVeN2iW6geQxF1gYnqfFJAdXcmVo0yCCOAIddzRrpGUg0PmG+fxUBiAfHT
uU2qN0e7sNaRuH7IVCRSPCTcHVaruHuDgLst09lgnlg4Z9tsxaWqM5/MvbSCValG
WTU4i4NTUXNo+hczskY8CIcl9Ox527kHQGVkZ/Q0FTcx0qPEbE3eVXKibUPF5z+3
AJWF+WVwTQStmraLw7KV9HSlhw+F+Zi9dvtKzZJOElA8S7X99Y13yYx/D1bblfHL
lkOZCCfEQXE82eNRZkEFAqu2gRq8qygFiGKa5FhzjT8KSqwwILLZ1rvAzW5srECe
sjoIAF+wVPZYyqQsNQ/rt+N023zBx5GPeWg7sdUADg3DCNtoGs/rJIYCd8kGXQ/D
RanokO9+xIEav6csz2wHZ2+LWucNa5uAqYXMiTLKQ6AhWDrgbrqr0Ee+czxCfFRH
J0xdY00CQ8VCiMxUyygCkkLKzAmADaEVDobUjkY864ObXci7DF2W0wmuRGaI/Bcv
9PgO8MKwhSKXOS9UsevAhXYJpWgwQ9D0ENNwwxn1YvwwfldZOwmWtyRZ5NuWwkDu
TOUXmJugFAXQMJ9D+NzczCv4ztr4YRzUxQSgRQd/6flYLxdRkpXZpMQ7RsHgMCgL
OxX4e0gJhZwYaWz2u/phUbFWmdzEdxBWc9d6jtBchrEJs5IUBfgiz7kFxhN9+mPA
vSFRmOrUJUNdeBMJ1d2Mm+kW1JJeQpwuXWHXbT58mwXzssUZJgsI3A8iubLHE7HM
TrOumhHkYeF3tBNOcQMruu6pG4RV47TvcEbIUHq0GJs0QAZ+IuGw67epng4W9Rm9
XYdeNXraC1LB7dOvLbh9y5MwlIBp8sKkpawDd0gb2pOZhhb3sRP/IH/SvUtuk1kV
4phqB4BBRKqqJ7HRRJCcmb9VdaFl2OG3ugYmBxSQuDavrWCwnHt8INfIHS05YnJn
FDQmZvha3q7FAhCPdqHLaiGujxBzPOQyiYCeM+VxVqNny1N58TYvY0SuN5wbEoQJ
un8ouDaHtEaT94kL+6XuINJJbAtiG3Af7p0s2pK7jGT/LpViqmJkTkqpdIs9ic6D
4Mu6tRBt2dOHbwHJ6RNzbidCGXnd5aUOgHnG7jemEmXgg3cgzxXPiOdIMmKdKxb6
s/nBvRgy9XzsfztcWsau5W3CMxr86ekcso62ldjuX4QkJVm1mJOSQ8mQAJwRMeJW
UKkeYxJwqV1ngDsY7Cwf168sIdwyVWELCon0l7wyMgfQpBUeoNBpBY3nZm2ZYPlc
0K3gUWavGqiv+iQG+GJUaZwSLD8V17322eZuHbtcnrNZ+If6zbn++mBBT32WGVhr
FRcQHOXgZq6jNgdPw7raKnnaPaC5aqQpEi9wcr3eopnnkKukUMDUym3OGtPMTb9i
tBHQFxfyoG3XoVH5HHH+UebMZ+coB3loXLndFLrBwwynBDyUnxFKW5AAJ94G18jZ
pM7x4zTq913tlu4EzgqnohbxLtGq2YCJ3MlnMFZbLZ6V4uNq2VCpHXE4ux4c6mAb
IBCdMuRaeHnHuhR3x0daV1ARqF2idYYe3M/XQhs+PsxCyJxFN1S/PUC/XYrcHJBj
vwpmUXxMUrro62UX1pFoKgrEvbEqQof5LmhSKW+vlUmEi1vcpIv0jurY7i+B+iIC
HFxj64V2h7HSLURJCKbhb1Jmqd1Wi7x1pVLkc4slOxbKIAYCNSu8OP9qMv3RkJLz
b8usO8jnT1aT03C8HewOb0mbAkNqia7L7C5fPa5umaMIAeYwsJvHHIR4tzTByNX4
+DF7vzhSXLlMViVrFDi0lj0QjA+FtD8uCXrEx3ewSJz9fET95vxJUXYdajXdtQ+3
9sK8ytchvWDFcJ70CFgSTQJQE2Gpm7whahU/IJWo0iFavw5Z5u4QWuALn6z8F4XB
JHFCQuNNw+iUPMjoFt1t/K0Vs0BRtWKEhUd21+v9j8vbzah9YCezfB7Q8XPn7uEA
x7HdC1F+eT6jXvwtDYc6wYhLNgZ4MdVHp2k4koKpCzX5oN1It7bwskPTSDRgOCr1
uhuj+lMuTTVWKGiMq4NXybDe2JlrWffXZPv6kd3TwWxjmhZbfbX70ucZ2Q1He6sL
JQqsUSlTDIMzDg4j53VwO352M+tborDtb5QZjigWAYImxhRD0glGUUz2H7sA7A20
H6+jxRt2IAxPXTO+dsOLWm+H2S2SvN9YLLPbLi27SIl+6Cfe513lkdwHs6totbD6
fjz6XnLec7WkxsZhlsYGEB1myscs+LVsVbVDR8ZaxyqFvYJfycHZhdg6PRUWG9+3
CV3g60aVKtRhrIuRxcWl8F3veP59ak7nlfzhf6ArRxbxeDbZ8yq3ZDHZ+lddEErw
iP8MW3AmzjSkb9jUs4dhC52q6NYrLFlegFjc1fgtvF+2gDrTetMRiNtR9TodKFJR
647A4atRntQwJF9PzaKWBE7t6z5DnKsNbFlAKHZEVqwqtSjO8kLyo47xRJmIvNE9
9b3iz3CZv7ts8O8CsWnxu2lWixecPo5d3jAvXHSGq/XcZWhruRWXWg662BhzfVkm
iGCJxbEQhUwHLF98Q+bDvgQYbyg/k7kOP3nyQWgAUgSRxeHS5j9/vpfmFnMmDvNg
eHJUihTXHLDqetZx9bGTrHtrOT2jH0WRI7zR4xei/9h4kw5UvhpyIT/UhUiaj/T2
XVDnta09/uvH+AVDPM09aZkoYWv0ZiFx523uZcsUKiTv1Axns62HwpoEsYQ5KzEx
9cczd03+4A2cS0wRitucU6m5W1Zs21+BA5v6DmwSdyOFYL/LOrpMHalCr2cOvcFC
A4BmvI9lLPuS95JUzZXIfQgpDbsn2GjKR7tJMZz6/mWhNx4e0oVNvp50xIOCGTwI
VzlDA2vYhMBX7VcqgWSl6gbGTK9OjSdZN0V0DRyDy4SuSRb9reBeiSDAGQX3cy40
4/Df0EjsLDkCWHQAjdULqwEFlfypxmEu9nYr9uWkzqgNcxRqcH4NBv1R3+kZkQnC
DN9gkHpWHqze2HaM6vxC8vcsCoJerZ7ODZvrDQ198q1lYNeT5GrgeEfQBbl0gCgC
nL9OTEFey+5UZuaHHkqWIT3Rt2iPRVGXsYilQ33pk6s78Bba307Z+ReZaRttVhNb
FlBF6wtZL9gYeMFICbB8r2eNHFIzg0lneiI+NrbPEJzUdkFi9PYjY2H1R2YmWgic
KmseiQ5X7ETXHgCITRBSWBgsorrlcM5AypscBEU8H3k8bZMceADnEH46HPIbMs8o
Nrcm5DoQ6cz6i1asgHhkWt5NE6Ut9HNSgZ6WC+3y0YRsw8ljNA7ofA3lpsj5eMlp
vW/IV5hJRDuIzKsRg3n77VljadBVYZzauhUW64Qw9gnr3FGqc257YrQllTzb1XIM
6ouueP5bIvG+QqJbItjLWvhuc5x932yIUaqo7fN3ozIwiC2PZ2zcj8JXKfqLFGdc
bJYm136xGxTEPFt7srsqYe8USFnLfonG9c1lROWanZKR/dRUwS8lFlET6RXRRWCa
t95A2bMXqDoBJt0pSRRjanomKLwfiWA+8EAVg6x/yZgQXIBUuF294tnO3R22tVcO
4yzThlbcoKOV41ArQKPBBcHcnD5+zAYnEvn9nsm3rCoC1JoILeCxhyRzDHvAkCTP
TcH80oQh3IDdOU8RKRSyqCGGyMFqv5MNSRinQrS6jntvbdkEKc5UiYNMUes1BM9k
OKKxrIRZx2RT/e6ytXzV0zdwCycSf3dbk1ejWVUpzc2/A73y2XwEXQGBfj4SdXqa
oMwsJr/tYb7888o412aXh5mcehkvPcnhBBWnOPupFs9RmbzVjV0irg6Lq3Jz6q+K
TD/PuaoyPJ3fHPnCzInTb2VzUpf6xFNYMZQrvb+jl1w1Nsld5DxDyYeB35/l33px
+/+6hKDjoLuzQkCk8DDU9iL/uB1dgTP87V2EJ9boWDcKB1kwKfOajTXFLvka+4cY
GClEfESklvS52rrFF7PieBecw1ym8VpMbxjMs6N6TGDejC/mu0Q+pQMKMhXMEQEH
fF2jaQfgzTGwxewaF/fxc8c0mUCfPUqaodUJXO5A2i2b0ZjPrIYye3uabqYRWW4g
223E5hg+4jzPorNZR5OU5UsYXpD7cNnfmBYzFsldDyrAEa0xE5h3ApsGLZleyjj+
Z+J/8U6WKOCcFcGh1xUk7bizZb5rOdSHTwVaDvnzPkkNIhjlrrNrd2ZHc+vDK1bE
3WD3PfB4xWfXjEIu72Yn9EomB03wQgjH+viZfjdDFD/pDpy4o1HJspR61bDmddBW
ZmbKZ+pg6CQwdZElPWk90Hj7D53UmH91Kgoqhj4OLQlo/NXeI+kYDvC8G6K68LW5
6M/T5bJBxK/7REoLAQU1SOS8b0Pwr/KH/HABp5vrGXS4kEUukVUjZ7S55D06VyDV
PO/ihlvvQ9r2psiyKWv0EitePPib4LLHz4e9N5fD68hsK6DkCyIs4anVE0jgn0ut
tCRYFAQTWvD8yTU9btDrZj5LaDRJSAzE2Cy17pD+UBa6auAl35G9IFJ2S0grLaaq
5NQpcYoF8xYLJk8lNxWIIfOxbfvL7p9r4rirWJffMwyrWeIjltnoqTHlqC83tXUe
5H2Fni6Kj1zl1G/yelrVI6Pqj0fCKIFe/rSai3S1PYEqTV7gftWOugEiGuUVF71n
wFCY8LerKsj6QBb9VYRrQtjLufbWvqe/vFot8kTa3RdJ2A3qEH2I0926SeL6rHOl
st8tZcX/3NoPwQJvL/KqaIKe8MZAchhgEWRAHYcIEBP3TN/lQEDLdZPpGWaaZVbw
gq/eegrHHUUyJWu3H4tPAyceRvmaIxQc5mkIS1v3AwNS8EfCZGwdmuYrrXfFeEiC
Nszddilj+V9SEiuZZNTkHhRVpx4SlNOWpxmtcDoikY4iyAmztRiP604irgY1rmzR
UIPiplioukm+KGkvi8Xmf9J/RK/v2hzBRxWUTKSsdV4FaunKkzXnMQKsB0zMU3Oe
Z3DD+XxBqow6OsSo5bksTV4lKLEltUgGX2KL7X8BpzCRwMrPTiceWialCbJ2TkjR
faRtpgaXzPpIW+1wa2jTNERaxmp4ztcZ4BfVzeITB1gMrgKzqvCSPuIZpZ3OrLEi
PWCXFHHroJI1ziW1ilMBZXfdSbr9G/ZSaJhFMRMVR6+tDg1L6SFKhURvXryO2Ob9
/hiXiaLIejS7FGXDhr3z4BgUILEQU5qjHfH+UzPEG8Gz9ikEHCloD86ZCtiKXU84
uzjwEsZ4X13fuQ/XwB6eYtzN7/KYZuoMj4Ax9zMQh+HuHct331Tm/U60CwRGEEoH
kk4X0W63hAZ56yeA8/KWdA1yzI55rUbc93WnBd2zTVc+A821467R5PCjsoaKMfTL
lTxpmNVMJt8hlRbe7gh9z9JaduDKXo7PRt4voDwPSQkGtVc68qskKw10NuT2gS71
dBuD1Op9ahZ3NJ9t6HOjsGgXbVhiltJH7c/vsuxnbt7VhArByJs4b4ecX4xeYl9h
Z/VszTfLSnhB2NglNop9BZGH91zcX1e3XwC5W/AS/vZKexuNAz8tSsmVheB9jvGL
NSj0lCarr3/2jSb0mYF+3AoQhLoYEqBWMvV0Asolk93wLkNLYcI6RszlQ5W6NGSY
xd0UPt5pS674icdM0BvnK6QfQk/jkzaFznUSlrzmwfyf4NWzhfTozjN46x3kM1Iu
gvFOVnk47uKuXo+MxU1IrwzMTicpxK9G4cOCWFGuo+tIc0cI+S9GiobvJsHFghmM
zWJvEBcouqgaGvHizaPhkyi+DtG9l6QUz9aHVxUXgxmYt1FmQmUBsZdN5rGai62x
YL8j6dPSJCVY4kIiEkPbWvWX8tkKUWY6kmkmFmDWuFhQ08B7kl9PwgRJhlIvtYkr
93YOL3amfJHd8vFFDO7P8wU0sqQ7zyo0P4pPsbsWwNlL3Nt9MtyPBIp/3V49laiD
yZepkMSqW3IM/NyTG3cRqKY/OjBXhDrh/dSntc4dNewp2QcHYkPYEFu1DqAZBY2e
YygQMJcS4cgIpS2dVYXaS1HrTfHpQjoL6/+yAiqSbQkMHdF4QzR2T2ugjHiuezrJ
NSMEMG19G4UHGRB/k1ESYBhraPmJsLA7RirsGNZDVZSiXOUJ1rqSBdDUspQ9s3Pu
mkStJIARnWkLgS4f4jauvT81f53pizM7vTnidy/3UArSs9fhJiDiig6vuDV0iY14
Lc/kPmtv5cHZ/4GT5p19z0D7xRBkD7ZMQ1HYq9o8sB6wkhC9To9E5l5ab0a+ohXp
hqFjNWsMgtrXYx+pRI0vLe/1yeIq+wJJdKl0Etg4tCr7OQGzQqyV2W3WVYkudx1M
wm0lAEP5tR+Xrk26495i/mQqUJ6h+8JqHt00dvND/dCT+PZFtiRWPgHG+K0oa3NA
l0R9bo5Ulu4VJekfkn5T4wpWgfnvdcR8boXER7vXL1mF6Q+DTC9UOKuysm8i/lz6
7QvFqC3ciR80uUw05oHPXAZkT5bmsnm+Wma35TvxoBWhjzL9/XWZOkXx+/wzSs4O
S470z5OwYEFVSa4NJXxBEbtMjWMHaBV+hQMs8n9ArTRteye54994lzVvHSJyi72B
6QaO6+ePO6YwQUFz0/5lL4CJEQvw5FYc/hHhQ0xdo5Aupcx2et1dIP3y/k8NVV3n
m4Frrd1mU/2FHCKctq2g6M7Qn1TNmfcNqtoZDE+4D6nslrEuw5lhfrkGuXhX4PvZ
PG+d0uRlhYqgUg/u+mjURb14et+/Pc+nyKTawwPVwlyLkgP0sgi2r3yk4ALo76Dd
tvUHDOCwK1DFMhpxgEKWbyWNwe/TCTVWpWU1l44hs4PEWb9PYJxY6SCIcKle6pQR
+aK2R2nOYHPqQ6hvJHkSL9HoF4vyBJ2McZgWzFTB92LnNa8hvGfdcwEyabc5DAsB
gaOxZhGhP1EAziPDOzkUjvGcWp6p+pVUS8EjPaPL217Td6GwxNCtlr2mLQHHzQdf
lWMI7S//Cp2zRqC8wzztO6kfv7yoNT8JweOua5jGNpxsN2s5xl723p38jBWH3F+b
U0YJugbnz8d/5/d40orvsECQ6Tt5WC7IhWEeM5p9eYs0wwNLRxftRvGUCVcGcmx6
3+SzGQNULMibSerQkT3G5oUVKX2Wce8gicz2HmhK8OawJMKE+L2c0YB0yqCPip2Q
U928rtBJAFdDkmvnVuGtyl5KAjw+I7pdXfcDuFFRS5qjmNMlw9IE8pARVnGjdzs+
jSQHHcS96GKskm/5hM9/K0OuCbqOwv18VA1g004is3mMtoEfaELt4kClff5w7KZ/
k04Pj+P99HYBe4kOodK/ke72GF+KIyhaa1vqYuVxG6GFf6QeVE0kboXMb9c3nYzq
qug9AjTDChKKeZqZKo+LJ+tnd4g+51Y+o28TjSodG0Du6EvbzZ756b7XoUnu4nMc
XKtcWuFhjPyl4CuWScf+K5zl3esQv/axdR/AQ5llDyupldBsIvry+5R0dAwQcePW
vVydJ7PTW5ekUnE//n06YRg3nL9WreMpGFxaqLmcx/hndpL16EXBh9RFfblmtwqr
PffuFXZjzaq8jgM/Go1EwITuXBIURCZfLV6YY0ve+JvLHpDBm98/x42jG/lu0zE9
vXqcHg/rHatCrPErgwALu3ljZxspJ5N5uxi5apkaAyzPaJbuNyNMIVlw8CBMg4+D
/AugAby/d6aZSzvT4Wdj/x3pKnhikmqr2fqsWbIeALxWY3jhuHPLVIj1RZ1zqHaR
rFpUSG8ilvlri7hOgw0nkp9O7Oe0AXhvrOoB7YjGYFxvQdQSw933JOiHplOIFsa8
SWwi96gdrYdB4ptqn50wEnGYRoiIcLXaxD1nduZdq4bxEqQ1a6f+azcX3DejT/i5
BlZiNhgpdmK/0ENSuNsx2W86CCD+GOpAnt6sfHIA8h1nkrfIrnW1TCwk4tMveY1i
6s1gNVZ56RZKzpbTODE2ieJqOo2IGOsydMQnfYxVySNQWYYBNApT3ei/eD/wNj0p
Im1n2yA9cY+lr0CeZZH1YbUOalBKzJ2fcIy0SuPB+ulKnjyUfYkV09WkfjM83sP9
qoR6pFIMNxdR2jlV0VJZKECC9uO1ZezydSKUUJ68izS8pecVM2Fm1gbM/qXueqWT
GYTPjvNL/Hb7mr789OGVCY/8/qiY0rsedTmNV0Ho5+48Rs/00WvHo4U1Nu6gIY0F
8XIr8YlULxFlFdEDEr/zO+vRGJQM+/unEo5uC7FQjR1JF0rR329cql5tM0cLowQd
wkbmWLuf+0v+f7xyFkzVED7yyjQ69mvX9icZtBPc+bDoHVVhVx12Jb3QaO5GvJTS
hXaYDIkpLUkI5zuuxX2r0PGYYiv2jl5d8S+QOSS4/SpqlT7+YJH86BOjNdEd8Csh
uGVnxjjuqqN5hRNmR/snLBfqqJUrpyO3geN3BfiHR8l9jZdCOK4jYW04RHAosrgf
jHhgkaQpij1jdxXm1xnVn87eT/xr/fyFq/yTGubBAOujoDO4rtoZNCLsgXB5WoJ+
4mQVuyMyVWoUvtJCSajvoOoZdIP7wW8G9PzfZ4Ey0mznh/ukS4SKLl4pVsplOPFJ
qsYaa41BMB+O7US6NpzpP6cxF4u11AackuR8NgaluFiGbgGYc+GBi4AARqbiplOs
9uccyTx15LS3LMFyHKjZKbRVllA5xlOvCJRBo5Hgy1stxHsFGN8bDcFhcNQHQMc5
Wals6ZkOzIhpxRMEstCe1F9IV0FVXJSxJaccOiPX2APudcJJb8464OiHU1VbsNBe
OilfxJp4xEeTAM9M1Z+ayScBDXGhM3R/MhL2kUoxwZo/gRLyAC65fwn9dG1fYwuK
Zp15Iu+ONBjit9lnMF5pZO85lxAFCNkUHR8SvMP1Forb08L/hv8Uac3vetnMrvRl
w4v0A5nT1U5etybC1gaeDFPSnenKTdtWTTxvSXU4IJrYACeSR/vY4sU+qC56z3yu
nSkfxIw4grkzAHKciClXpJaVfvad2pma6j3TVIJ9ZwU8C+DztPa/fOiWHSSTI+U2
ONz7XcwJ2NR3CzDl2z/lJfkuTUhZZoPZx1hleJw7GpbRUJhG7swbJ5p5/VOevFSi
DSjvFIe1xfbUBA6+nL0DypQ9sK31QOLAbNkVbWdtyPxfCu4t6g9iTOkrmbRZv3xD
Uv1EroX+l9GrI0Jw8v6fnEaW4CX88NTi4oH1bb8YcNhjBu0+Rdw8qxPLxvoCqHo4
f7K+dJ/JkVX4AassagLUQTTsYvpfxY5/e5UiecM2BKw1JZOrjs3slYgaANtWtpB1
b8IBKe648K/ypv7lJQM4cVVu1+AHtH2aiMlV6xgx20PgnES6hkWRYn3k8valTq6I
N1yLIqZirQluFoyEqHLCJtw5ACslP5OT7g2gGJLvrHu201aJdQVDMVIFCmT5bGAc
KsImy6TP7lwShFAQJoY9GkY31hYnz7C6O6uXE1YUi3wjs73gc00bwqb36r0gln7T
SchW/7P9Uxh078N9DncOi8QXSqoyX8WYTcQOtWZMPC89g8g8/SVQMftswha9tZRq
a8pQ5apvlwCfV6WFYULVZ4Y8Bc896ri1VqCY8owx3llBVq9PICd2MTNkHx9vJgx2
vRwqKJfXdlcB4M4UwMVWHxhDB69jRJ5U2DhoHhcanooKxutZN+fHKX4d+NMqOnJ8
JVAE6znZNI1F27aVL9aOoG0t58GjbTfW35A0NAkfCWlruDiyHRP7CS5p2JyTVVeG
lbb5/SZ+dqzAfNZCccKbJUdFQgN55egbtipUS28FuCRC4fx9VTkVAltKC3a/J07e
4kELdcKYcaeE5zES+shvCjXQvrmTW7TEdyVCvcmpFxWRlWo+KiSxy0XWBlHC6Bcw
U3xP37Nv6TQHDPLDaA0Ya8cNBcyISdlPGQXB6kN0uyBcIGrYPgBMe9Gv1Ffi4WzN
ST8ugSNbstMrrEzSOULuiG9C8ly9ERcT/blDm+UUKrCroorHnRF9M19jQWrE8frn
CvEDchlD+PTvooS0Sn0kLWO77oYFfs5CPqL0fclY4lFKKsHeQ9tqMY+qN2KcZkeF
p+1mkxEd+B/agfF/MTben85SgMpT0vDK6k/5DWvqTsyRG9988aSMkBpnzoBwTgt7
ovgeyZy1IdTVvD1/wR/5mg/snx/ooKlnTbzlxFy7FCOIT3HjM2WMUzG4Rrlxqn8+
XdMf8Op+upByNoT/4X4hPHQXrgNHQVaghvH+AJJUkbx/CjpL66yLag/ZCJwNarom
OyL6MK6Wy50nvEOBT4uhdVoAwgy3hp+o3HkoUCWGRTbIjI4Jzy1sSP1kcz+mntgT
sx37Sd/Ks+1mBl5+Px6/EWEBrjetmxVYVtPreDQ/HX+0G8qrAl8KPMo31qKX16iJ
al9HW+lQWDpUIy2UIaCS+1vzh6svVueVegHBlwQbPzVlh4evwyfCiTiKcNtQ+o0f
SxJv0wOo4IVYG7fX8OIWhSl6u29OImJZAhk/2J8BA3rwvsiIlmDqXP8fn/RHjKhB
yo8PH9dh/zrd6uV2IKW6GML3yokORoRAaDXbkul367TaqO4pyM88gOwgOOTXvGVA
VfUh1Q3uExySe2yrF4xRt5MWlgOQEWDo+9qdoYr3aA4HZrDxLNQ1zBkzON87RgJR
W5gtsPB82LGKQheM5FyhoPHTEH94QjztCUHMncrCtKGYHV/y8jgpsdwXAwP/b5un
9sXzLDcXdtn8sOk/xkjEEfAfW98zj2is8rAj9JqT6UeeMsCohiSRxhrx94Fy3JU+
x2WiVC9H5h+5tgHt8khI5AH9/StWsZzYFckyWFk8SSgmQvX5LCGRA+jNOl6V+oH3
3HQRSsFqDY/SFuiLOO0g+8jas82g2fOjz4lONXxZPLL54SkdCDHoXmbwyxrQCiJr
mkZLGTOLQA+87FJI5mbyrALr2Gr7awIughbrg6obxzn80xeJ2xqsgnqYC16BbZNn
O8d+TqHBTX33hY2Ux02aQ654xVA1EhNPC8Pcfi7qqWoQ/l/vK3SbVGL8beeTUg1c
ZkYzE2Ak7EDy+HgISk/nEDJwKj44qvnAulcJC58QcMGEtq5uoUg+U1yIk6am6ahc
3c20gst3L96Px6Rkza0qcFiV3WXi8t0ptfvhxvc9nw1gAYAAhL6ZxNQnGMqkKKjy
kSN7PyB7I9ZMkQrSwkVxtWWHYYGeOr7WQr5FLq4ppsTHNfrnIRDnkn8+2hjFlKEF
8nd8zlUYGgJO6hNB3ni+4gyhHBvp9fcXMot0Rm3HN+IfPS2UmT+9z0MGQQWkq1h1
RospQCCAnxW2NNNI0USfBpLnqwpPV+VGXAh9cWNy/HTxLrUJ7KeS9e5PkH6UgtWQ
e1wAMASmXeQsL+D7r1pwLCWd987bpaj7L+U8LGaU240Q88Z070fJEMlSEkzpmR4g
w/4+ct0UJH+iXmLqaMp6KEl0DPwHYqtpLt1IXObY9dBs2yRWUAGwqs8puZBWSw+q
F358CTrS3g3PaxodV32Qu0NYPQwtfNzUMH2QaQtjZc7LkiM8ucIkna95VgCwAQTH
Tbkq4vgHDLp2c4ox8YZHPbA2EdWXJbcn3hYAc3jyF5EohqThzbf4Y/eET7kBX91s
58YHHqDt9azdh0Z5v2VFODvtfNODRMaPe81kPB1TTsMq4eVWSIwzyFh8D7uoZA4z
6iXQ8s89Oslqm/5KRhs+/veN7b31VmXeLRHEt2aj6uIa0KJKY2VHVk9Mh3hNimUn
xhQcmRwYtNdqP1OCZqXJiyiauJAgYkUfvp+GhmsYddDAFO7ASQA3WH9pvxZLioIb
0FdSVKJrQAdBNZBlnxwvgCsklbb1fFIJZ12pP+TT0LK4RwvV5rZKrOAvlsldNbaH
893xYIJawG6hGxChE83yqfZu/xhMskspcmngn+YCKRj75juyR7BizyRDctWwklG6
mCAYJZYJtULzi4DoTgE9pR5SfE5BKws2+cMfyj7TcDiNvIEYpOQiSZQXEa0OEek6
DRa/BThJF1ssjQ31+69wjlB6KFIxCWLVLx2AKBABlllcsv/mzI+HViCVPWoML7Y3
HW8bksAP+uuh7Gri7jVG6VcaLf3cN+qp2ToxPzUQitgjV2GSP0aDzyFXtiLH3i9p
fzFgLU2U23802Xoht53xHZsg4TDTaK5nTN/r1PB4eN1uf9u/4UAknho1eo0ZQuP0
mBfJ4Rzbps8pveajCAd1kOj5KvqwNzRF7qbS8AMkWTgdW0lxsafgSrxagP2RJ8bU
FUgHkbHOcdDgLV8XnvTLBOiyemhmWjuT9pvfTwOzBBF2r2gaJAMX/i0FAb5yX9Mh
tGrCBGVAtw/BFqxgOnwSRNcE5TB1QVPR3AbDNHVsRPyK326PRNMs/tjun7LKbht2
E0XqJ3ykZLqwV0z51NBNptv6jZHYshrCAmKgkXnbU8WphlkP1lATQ8XXNhmUElHV
y0CO2DGULzb+B4yqpWpCMkZ/OJ69hOdTCNkruxPNaoi4jax6PzBEyq/g6sxxzhOW
RTs8clDOHVVI17iy5HD07llRgrVGN/IYA3YpM352mwJE5DlRd3BuMjhS4S+edWby
/Nz+w7ZQnxY3Mc1LESobhnA2xriCMw1JktrPWOdjvt5zMt7p1QulbU3qyKGNXiCp
njvUpGKRCFkHPCEqYkawnGhwchY250zFQ4QkrL1Ti1vm8rbQL3c+jjkwIoLpmQYr
060NFpaOWtajyqrj0Z0UfFS4b18NKTCBUYL1P+xa/Cm10PYxBW+79gqgGoLDA+da
V9ON9BBBdXlLr650YPY53+xtyoD5dpIYLizrsDlSSPFu24yDtTLqYC1Ei7dV0h//
/JS3erSooOB1z/VN2su4vtoWDFDtNilQcIr5ZdPv1cIeNLCydVdGHgLGEJOOn5r2
WuHOsoZ0qn9LheYyF4/BKsUWgeQsBgoZSOsvpl/goQgZoKAgpxPilR1BtPutXDH/
MQb/IG7JnLguj119MN/PfoBQyuktJSfc88VetLxBLLxykIAhUYOY13bgSVtPg6D/
jMFl1IREzS/OCeQdryw7Rcayq/PBeWi6Kk+FdBt6KYwqYkTQghbdj9XF9/5x8AaR
SNRpGkissucJIMWNdz7Q+h5CbJyNk/nn4KN0Yo0oM9Ev7Px3jiDLEU88WhgbUj/J
C947/BzC851SLJ4WtZUbhvSMwAGubm1rI91IKmNBr+n3V2eTDxwPnI+BFfbMH6Da
oM6BlRQhHlV/7tzYQZoeA4GHvumqLGRY9Pz37BmgQ3SATjN/RlZGaXUcGiaSgJAG
boVIWWlAAX1c2zO7pzfhZWxTHOT6q/ypvAa9htLr5J5f+/8p9ec/akVaR7Ek+NTV
DYC7mUfkoJR+rIgW6qpU4TFzOD3doagGosRGeCGq/fnVUfbdUZon/2d5LyC0+dyZ
75TlQJfiIxQoyxDksruq8nKtZwU4Tym3dPF2VWCZvbUagarJ+WVWqAPf9t1Yuww5
GZd8Ceup4DEnw2s3fqUAeEHSlefOOsiUb4l/zI0c5XoQNQKpInyAwFsweFGx2SAj
EMNmG3P8ysvJtiUEoPxu/qgFjtyb0KI3NvpXLVPYKV5kclDenEt8z+AnuI30QJUF
CErKmaCz0iIJNDc2d/H8WIWwFySoad829eUcabaetSpR2Z35sWjSnlOpfLkXVb6j
pkyO9jOKWtlGIvJqYMK9lAv/S6Ybj3PiASf2VCIvl9SC7+t81GMHsd+wwU77lvhy
Db30p8gf4imIhqro3oUkf7mnUvo0Cp5qhXKeX2Av2NiGMTwndBNWUz++9Q/0z21J
1AO/iON/dQtr8FfJ96vcnAEpqxZbBcyXfpJrR9DCIr7PnqrmPIyLwOmKWYIqG52a
KC8xIrkyQyC3492nmsm90KDkamis7TDRmRPaOQTitNZnfqA14WhXb2E7bUgOSCQj
fY4pFLKl8FQ8hjkpa9i3wCZ84q0dei2Tjd+u4fvv0Syx2T8ms3BgEh0Pl6wBBN0o
lOvxu1eLeubwy30I8rWaNYr1tqXc6KAbOg+dj8/ZbTls6OcaI4csLV/lQdhUIH70
jsAop5l+9tGl7yTTQsj/FNYTVSxk2a1WZZExo8vqw44VwyyjEJqMqvmf/t0L10M2
0RLE/A9e6KU2WzjzmVcbkLWt2svA6+QzrDnyUiGWSKZCY9XpHAR9SiXR6xeVGx3S
81Cz9ieeDE3dhjfsSxbVC59tgBWTk0P7d2DQLVWw5ikeUeBtn6uDmBT/xzGABFPP
xAZjrIfFTZQ4ZJ8rZLUnEayau/kO8e3JMXyqOBavNlflcAbZ/0MZu4EvoQzbkXyV
fAGYgeFc+bwPHPlrJBe7MeLd5ocoxg08vg0dd3r/bCjQUZtWwGhzTQWkjUmgjtES
0UoJPIJ5bEZlRWJdt8vAtKK5BFpXcmQhtJU7a+DB4QETON9eZhnOEWY3WcMufPut
MWx2aEnpfFTLYN+cDxmJeCCXKesk8aAklZ1JNhI75NZSucYPQB+0z7mdw9/vO1je
SWUxWflnJmbPdynKMhKafRiVRzp68fpIBMUMZvn5wBbT2a/IjjnUcgNrIwpcJQNy
7nKgdCTuzaXZQLS8pqNM0W9VzOzLsQx6UVlQQhy4e9G5zJESzwI+1XZdrUd+nU4j
rEMixmDMcVH+ILY3xLhwcutjE5LXJe62UWub73E3b+djlEHRhbmBiLUmD0Swckhx
7lbELmvV0aXEam5PBj25r8sEy3FUwafEaaPCAqvUGU6XRwK37m5MqHKw5EpzGO+F
RRResJRch8KZbq3qKfk/F/KAXAVNNHifXNiASTQ3MoTp0w35wAHwCSNp+KhuXtMU
ZT7XpoAozkUvPcrndl4LxAjTQQlIGdDQSz/tkELYtaEyW4RxPFhGuM+bq16GUpPr
VZ0IRU+k7zLAB/DehN+y1zP9j/0tg0GgCTPyMK6T7XPhowya80Xh7Cs2CaM3vdce
xBnd/UzVCXpUpGWwFFb0qNblfD4t47Ohg0udUi4Tp4yE87iVnTV3EnmNj8bCTbMM
6NEMtvz75pWH/+VVOkxGg0oBUgsUE9FsSjNxYtrbRghr76A2Zu4JzcpglaMSkuDI
cQ6tpXRNWVbhQp2l7jijV9sf1ljUKwN6QKZSUJeu6vvuFFwlwjWvjyQcV8ipc3HS
sbyXpznrH6+E6uUXVSFi52rcEUHDt1xCOfdKg0LMQro1It6QR4cy8a3D47Y0LJUT
m9eIa4ggKJ6EqOfTi4K10HPLX7dpPRBeh7H/HoCM00ZcF7wHjwczSbC+IWbv/4uz
A6NZpl192ZfNy9flAZBZ0iI7FCeCkjYf4nV+HBfwqCUA/r9H3qN3A25dz5OvfLBO
XygQTS9pFwAwZ6vLZ75N9t1a/T9nuYQCbzyCpv8ksBj6rIDW8GiD4DNWb2M6uTVU
r/URKCExaPxH3vQ1Krj0mBvaJCIW7Cef5pFUczLSzyWgJvbvlUNAw1ZTMThATzBk
iYPgdIeK4PBCaTlAd/pMsCZaMoOMRVRjKha/3CEuXwaGnx+IoTfjgdVDhpJpOVOI
WOvCT+TOClzAclVeMTVu2JdqQGeqZ8t7N9/dfGHPvAKgwkZErOC6HFXEJkru1H1C
qHLB6jPukaTAF1NB97kVc3mq0PrNhtAaIvNC6yHXcxqrPAJtrIgA035cV4Hkd/wR
7nkOgc/sUKmuAhWcC0m2hgZruSu/08GsW/FiZyD1+BMAzDabHm6J0HDVxqN3TGmW
hdyAxUcwRjZ4Gi6qfeJagLLDsnrn8ygahUB0AQFR9ti8aUgUd0po+hWzv2YD0W9X
QQzNU/XWvCQLfrDlUSm5LQRN9R4IWi2S1lgIfH7jVn9DI1kI1mFIbXu9PMJw510s
CfQWAbMJqyl2Tf/DAHENfN2ODwGKjHdD6n6f/hTfG2EhZYgAyOEMfhvoNCc3iRwu
0GYdd+T3+CnsWRz8vXv/f5nccmICpqjU2R9xDCf0IUpUY55MTAYLjT3ppmbYFjok
7vIRBUXYiGu/a2zAOpD7bfgBCDVM0C1gcxW6GBqI9vAzRwv5RreHRysrJ1SsA1nS
7+cnPVLkWPwuWOIZc5szgSMQEzVhSRljRAop6vMTj6Mv39Vx1CHeX50zsHMRetcS
JDK+HA5BX8pifRcIURQ54HtcjjCfZFOASD23IePc8EUx1xTBih3r0ytGmkT1T88N
pJ2Mivv3Tc8f38LADEEkNMcT3hcbIWkFC3jI/RzqzicBZnXWZsr+fh0irxooRO/N
c2G0aXw1EMiC9FD3i5v93Yiv51rMi38sMneykeKJF7U5ic4XBfc5WZhNHmMS7TUr
bsdhCARcfhR3MWnFNdutAKnmyBalsZUgqHkNVuC7/PZo8Un6L77F/e5F8GoZRebO
pbXu1hBuOj3wODpa3BDMQ74zfeiYedRGSYHrxWmdwxUy3FgXYL5pYu/+ARlkFZhO
UuAdS74kkohYx2q3rxsZf5idg55PfYLQ1N0FitUCnYB+sVhmeya/lAZmKLduGj3Z
ISvBW0BtppGW+Eo9UhHOGGcQh+cxxHepsyk9IJlJU+tNF87IdzAl44pAk+4tmLXt
bL5I8dOFD4V36VbK8Cyc7c2bMn3/ubrQ54fsgWMulFuv4CU1YzBL7b0lAwNRatPj
6bhqz6hbsmEGlMO00yxWoL3gYEArG7opTbyFx4Eby4d3DqccMbcrAlBgV1g/2xrQ
rhz+Oqlk1uWY0KYl9SQWVCXc3+MUeP4vpBwFdB8N0AVcte0lIxkX4xZYkjF0MsVb
J/ODcWzFDIhSLfXOK1p9FZgeWvWF0HUpg1S45vFjR4+zsk5+dOgCEAqpEgHlMsPh
Ncv6APW48x+auw7ooizHk0SuqJ2T4is9SN1CTouCEsk1tfT65lbmE7mxFwm+v6WO
VYppGWXsvIGe+ohmBd9g/vIEOo2TA/L5jSvtaw9qn8XP3emqCzGCIv7Tg3XhCN7e
+nX+Q2dPlqj4zEC8zaVB5XdkOAfPoegirmQPogVSNL2TN9sIR+xjE6OX8/ReLWOx
ElcdZB2ZCFi+bA76ohBT93DoMsSK+aIeyB4v0ae/4B/7i5HzAr8/4L7I3TkamyEx
51mO0VFCjcfY0F7YxzJLWkNBgV3iHJOenqAcwQ1N3xsFrGaCqZVwogVXmveCTQjg
3cIUj82myf1dsdqVpMO228J0XjG3LmnDpEjKnO2OPLfL+pB+B9tsP0gutXmnPVP9
18stTY8p12jv6FF672ydsTH97rG8zJrUbsVP9Tq2/PlIGNB2n0Ijfg5/njinvtAk
xH18KzagZHqnrDcVQVfeBVGasGSRtnZH9sMKOVi+iH8GhUwEb3aeZZ7eJfhdQWUX
AaAHjM5cha+z+RIy/Df969jsmTSQhYIrTaQIHqZ1Esa4aL9OfibJe/48VBoj93ne
p1idz6arGYPT5Ni+bYjaqsZQYSl7wTYn3ccSvP0cwSLiCwSZXyHxYyfim3d7bJFc
dLOFD7uHVIWMNun3lrevvadgFQiaEEwpkcnlvfLJVkJ6od4YxsUoZgvWbsh398vu
DZVGtFKnHthNn4IvGbj3AMaCtx+g3R+/83CY3UNSM730hUzcLxSY4rHLpO4Cs2UZ
573yLSjAgs/ztVCxa/7lVyXiQqmPt7T5H9UEQ7eVptB60d81c7cw7H9NimG2JtKd
tTi5aHQ1OKJUPOVRxetxS5jsKxvZqmINDyOtsLl7SqqotdVIc13sK6nJPwg0rHGh
RX0p1LVoN1XRadDgzmnQc6YJb8xEgay5GQzkYgrYyBkehWg20TtpDguIk3dkyc04
0ad9B16U/N9WCx1Vl/E3kPbz5Ecmbb8wiDHfE9cutvhPdTR3Mat4WGgWQ/EWRvwo
nCP3tGvyx3TRFi7D4hL73nvexM4uoR4uSx07DXoNMex7fToKLefw96c0RdAxLrKG
K8D7uRdHwiTsKluW4sYLyeXq0nCwf8hftFf7vhdl9awYn43H+tduwhMIdbU9MyxP
lll13bNkC8V0IMvxz/a8ncX4zPO/36OOZAKDrDlSbKAfAZwSdnZSobdyPyKvciFv
Kd31ZJWk/nxq1shxClDwmKMGeFNb2Ox3e73QVIp4eqL9QWLDlk6im9CB3TKUjJJg
ws5LuzogNpJJhO06IfHMOP4zO30Qofgg3ru81AN79Y3r8seZNZOd1gZsCXmzbdBD
owR8WoHBsCFEHZEa31Jl/E2kGV4rqpuDSyuxMaJKWFYb4dOSBJN4ShOiR1Hqx4oa
lfOVgQgPG+ZG81nC0GIPcXJksYiGYc14/MWfUwx89EXYspgXsXkorDaySYw4ws1n
Kl89qkMrK1kgbSzRyspmj+zh4zV0EJJAwDYDmOBBuD2bqDAAQnz2S+uq3zADxPfY
X10RPL5mTUY19MF8GDaM3HM6DRfxInUskh/Il9IyV/j53K449qg4XCqZp6cI4Eim
qRZeRGmEZSo1yk0ta1ejPlSr0/M248eyEXfvulT6s9Mv8aQrTWAop58LdKmOVPei
VOL/UhF37nLInUQ31FRHe4DE+9vfPpXLMz8KU3gNgx/wWT8cHP53LsrIyyvWCSpy
vjfyXYe/rlYVqJZjPc8rJmrV6iiFqNSp6i0U5SZaGsXj8etxa0HKJjqaKEQMxsM/
tzfWNE2/gJgXm39WyPN6UN3D8M1qmQELdbTQbxN8i4Fi/BoAlet1wneOM1XVwpL6
oI8+HPmzZvB5liSSoyNTvt9Z61fu02tsO9ZIujEvATSsEOZSwn8mhAsKhU0cFRnr
/Zmj80xqk2yUCCxjci6ABxfFDsWX3amYVMWDzhVkVnwIviWNI4iEx3U+uu0Pp/S3
22/9xmmjOhMGhEI8Oy1BQB2J1B5Q+Iqvia3/0X2rc7JboGh3OboK/Q7eWdxM6x9D
Kp4/3n//saOOskYB3yg9ylGZ7JTsv2yEGa9JeRRXgftGnUvui9WGr//QBh50mv5B
pU1nHS7jX4EVZ3s7PnvYbardm05cOJE4aBiq+xDxF36vQtAV2ocADq/1uhRHbwWg
UepSlsEwigv9RqnYsuvff7fj/H755Y/7Sy0B6RiCtQ93FyqB64rm+GhvFUY21aXh
zikeMe6SY3YyC5ATaKeAPpP0VEY6za6Cd4dEM1jIL8irWiM8ugiZXgcF989kRuEP
4Vpazb4av/r2+D02vb5wYvvqox6X9Ryx+cZd+BBH9f4EEUQqoJdlp6GCpRM4wlBk
8/lufK5y8KHoZP7yfiAg1RT5ZhCg0pvDlOABGKFuASTqnxdNvasTG26ZxuQ991od
bKsU0AtAYQ3ingS7Y/sUTt0Nj14uZliSJ3sfqStca0SAAu9GY+A9e9zyUufR+5W7
po9oYa+r5ghpNH94pmLNp9Hw4Ex0KzyYLWcIxaSlFZNhv1GKsSeIxYmY7tTykxPi
QezqHhPS3fm8EZ+5ZMk5ejrCN33xJkLdPfhKn1QgZIl5dsyONYIKdoVIQCChEaiI
dGa8VXOjpt/8iE2W0hFIsAWyxPaUnwW0EyFaXmLCDtsS+ISAv6f6JVe2tOi6sw0i
rtT7R2ZErjfFyD5X9SO5d1HojNsNnneXXTejlCDQDmx2Jg23vHhYoo5HZqQvBTA5
pKtun51ACEHfvDqSXJ3enXDgt5RDShKsWypxYldiyqIBB5c2xv8CtZOTEKnp72RL
/3Ff+jb4571HgVnzNXB4+GLv/dZGWBNq5x4UebKIfXbbmBEfTqX0C6eg0Oxf9XBC
Bxx3y3Ku3MifcOf8VChevetyaovnMXSgygfoI3Q8SDv68kwieexnXXU44tJ8G+p0
sfwohS1HhjIwuyW5cksn1yE6t60SJbd4M5Y29NWVxfPn6pmaFOP7n7wVcOT2xqDW
RBulxoyDJTTyDrgtpiQaVYuCz+4FwfcJzqyJ0BeHypgcDzzDEWoVyVk1oIuVv1My
Kf1GnJIeizLOkKpsQKqQ1P0kUb9sLTVWmK60rBbZxRqiZYQ1a/gFeTqCpJxWxodL
bdej0PsnDx6COKi1eQlYwt4Og1hsy9bggk9h6NUgt7/C+VelKo1iNcW/amWcVt6I
yKUDFjUw4MAH9rxLaXh97T3xV3psVVE4h0QbaKXgruuJ2ZMmlwk39Alyj6oT6JpF
yX8reYMrFVji0/mY7Yca32DvzAyRJzcSw5i35S6F5J9xP2M9Bk3WPDsmMaMdA9Uk
AX7svTd3uDwHbaNranIbvBXP+bi7GPA10lctV0vIistSZVgkq8U0Y2O/U9JvLdOE
xqOns3EnhrDbm67p/JCOHw==
`protect end_protected