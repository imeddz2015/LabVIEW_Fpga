`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 63440 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/9huKRhRMtvnNqb3Z+UU7TahEoHV+T8U3P3ufru7l1O
3DlgtZzb9QxCbOjthp9+wDkjygH0eUfDrEl1ovhZG60O6SJepldZT5Lgi1x1hZE/
BpS64Ms3kqYnaOJs7bAArtzlc+zv7jYEWOrGKC0C/sBHzWD/cZzWQtDxpqmlZ6Jw
EeBhVMIjxmDIEo2rk6GoNnFrW0yvaeMeH3hOnkAOGUJU/lcsgP1HbePluInlWC3l
nyZFX2/FnNST4zuTDbTXAcXOBKaTQEa9n+EXdeXzbOVBX3g7uRSN0SveipDPTXu+
CZHzowg+P95v/mJQpM3ckRs8yj3nwcYkfzrVeUEv/12C911/GqRoTXt4KyOkJZRq
XC6aCWGBhb2sdnQIT72zeqKi84vFPbuZs8SHouhOx6zhQMfCcKS8LgrCj4Pvp6ul
BYVJ0M+ST/g4CSx4Sysulfm++NrVpxXgY2y4mRnRSBgMCED1YhOH72kRo4O2pGhV
V5CC3PsoCGG+/Ux7JAvb/M6MGVucAgdsJBCOnRtStbjFc64syILRAPwGjsisjb6Z
B6gpu7Pt2Mzzo/51c1kaqlpY330wQCLx0/bGzVjqsIpByVadxyAcM5tEEz1xR12m
MdCKk4nzonNtkPtyXrSUTKLfp7cttq6DTIePI88362OtgrqMyi+YffhXECpbDuhA
T3HcgjSSffsrI1JpjjAT3mo3oxGrWdZkehBc3XFaTsNLaKXqsClz+01y/WEcC9ME
FCt6J050A5OYgauQzHsboiTzZzTvPzxvtxp9Z1v8QvbCDbfAY8EZ5snsXtk9lszQ
DRlzKy9c2hsaFL/n6X3vIkSvK4zgWOVhK9XfIICvmpkKQeyXVshgtZTcnikp1+tW
HwfE/XhJH2ILSMymXehEEWXbZUxIn1lHIcj8Ap+Y0LHbns78KKrN01L7O+8uowBM
83Jhx42pecAWbT7kWgmwSLUAjuH8A+WAOZO6Rr7DSkYl4yO0m2vkn6IBOPu8igty
HNi+SrA37voDAiMpj2lJG+Pic9DpaLN+UfQpqzS3He45genqMeYbYvmQp8ftrm67
7YYVZwUwd0QFkU0D10P+sK+2HRP09uXN/ONxzNLst56rhQcC8EIuGtGk9GWK2MFy
bgWF+QlCzuB/HInVrMu5/M2Gz2Hs6MQdnLMooBYAcNfInfvki7uW6l8TGQomAJlQ
7iRFVYKKWVxUzx0en0gjKGIW7S0xUY5uB0l+rBfKXZpBbGyDMKn6iAXjpLkxjORk
9dA+lUU1ma9mqmuzMpw4vHGXaZ9eOu2fP0e8Vhmynvc58+LI87dsaDDz0iWuKmeE
gki2y6d4vN1IGNDg6+gg2NUgu/raauzDwVqwkDy+9+R9Zy4+Hd+wkizbm7Fr5CQv
ECJ7Of2ZcJ+BwA7YrR1oFbHCZvAIQWGFO783/QxnPOH70awyTQkzgAufZ0VyU9ak
CGBAxzIuUFdtCmcx4sVOZwSsQj0gHaUht1Hwb5y70Dw2W6USqiHZoVHk/zOzSMqp
mQNUjqErg8srzBvUhguq6iWg7vXbyDTiIEROStAzMDfiOTu0XnU6efY/SrUd4bIH
M31Iwe96qdp1z6d1myPF1KTobvqcDHj6bh/JDJahMYXfDHd9MRylk3JYEbOjp7nP
jr+M5m5AEjg4atE3wqWtNw6BNuxzwgZ60FBWTztkX1zmGtm145FJmP57dKAu7fkQ
I0YAKrce157LKV23JFYizqvJQElMVeyL0QqDZAMhcmYv2uc4n4il/IWv3E/8X4Eg
MMWYnmaBDyUSUFxESBGDePPx/KkT744+mJOcA80yNUKfAt0KuyXmb4MJpNRcQ4ht
3qVot+sgacgBDcbt3ZFKiC0gOMPgceX8o31+HISL31MyjYp/11giTGiByJR+L1Ek
6cH2QCkVj5gwD2GjfNH8xL6fzGgGABysFXMcY6T2TdKdaNLXf/eg106StFTQi63r
Vvj/bIh+SvanjlQImc28icjE9RcVSWhx0pWsSbGRZ3NBeJd8EAKf1srjacqPmU0J
CgSk+pH7FvQ/TUk48CS0uzkXYpmUmE5wgSgyjWZWFzhKwXo3AJTcmz8y7G8qQOm0
9oRkwV1rw5WVLr+3Glw77BPebl0G5izhIy+638+30jwK6gB67a0P6aQ6dZ69zXyA
feAhhbWrMBjDf9vY36T+OwCSZmzkkPp3h2AvVGltyMmZ5LvFUgv4dxclXhou8rAD
YtDZg1OYXhxLZKvjCndLI4QIPhYA4TyyFPZLI7G2hrBCGEAKqK3ut/XhNqdK4umv
7hF5+tKqc5yLPK5YHkCOlnhIU81isY7aCR4plQ70CeQ1544Ccuycy/Ru456+Sp8o
Hm/ijlD21HSFJnN7pC9Y+k64SA8xHWV+oSjNfkKieJJPTHh1hpKwajH+HouGYDPs
yKGnAB0EtEaN+Bg5Uqwnsk2lgWxjkRQ6R91tLeSoWok2Dn9JDwFAQ+bobgG7JRxj
ISCURsOcA3YQxUGMDh3zZ+siaBrCAzQi3qqmQk0EC0NrhVcmt2oc7ph81J86gPbr
dlq1G76kBjiePRE//4GqBFwnXU/ku7KUqc36wOxCsvs75acBzyG0G/GlpvAJC4uF
xBKf4EmK7SKjlODdq3dgPBPDC9lnTfJVzHB2x1i+Gxzrz2h5cjCG8l6PbMBCtQSE
ZHLOK2q80hbUaKsf5dk5zc7oSMGESaiHGEeK6b2aleZx27RUtvwBDSLFGuoZFfe4
cyaPUHbHG7F1DeRNZBcePsCGLh9vkyrCvQCbcq+7XTFKua4OpxsqKowthlds/nYT
8RlqXU/SfbojPtbEtNaUC2lty99f+eMC8ko+sDIiBsnGMu9hl7cPxgr+7tr1cu+s
nUU+3toMRsF2IGluWuw/KkI3lwaukqY8dR0kB8ONCmH0MORHk62nILYZm0y8F31R
5laxU/12TnQrtZO+rS8Fep3bpDM8jkfjqWSb7z/CyVoWHVV3GUSU8Q2niEptHuCy
+jfI4A+BCKNzHpNaQvs+P925FJIJwFJYwxCVEdBkBmkwMDrxGXqy7PzDoyH0QDcI
uA4sN09Sl8uxspH7gRQ/wUVT4GBbYekZJVE/IjOv+B33SBIIhZ6OSeVgGqoFMzdH
i2IFWt0svulYCK3q/gpYs/9P4KYxSQd3dEQKzGxumleiUt7YgkQm0UkFhFiIP3vw
r7asoUi48+4EPLUMzyaWl9+v96RHYzkJ3Q4QIrt/ejSY19NyNNLnlW+6KbExQN6X
00y9ug1ZR2MuZMgz3G1u06749Zp5aoH1ZJ0of2tDyNHydn1HKUPu5GsPWs1j2ADt
XRkdDPQ5pG5d7VS61b3hwINtImom3n2D/pRW4OY9roDDZQ+B1ToBNdXIbTYrmIWR
RLUUHMz1pYVx6fbFOypEDuJ1/jfHfXwzaV0duxBNHkv1vzsagBThZ48LnwaCoxe4
7D4XwyJU9TWr6IMPHuWBifOg/URYvvxKYyH90/WrFDgQQYs9nxDzh/3E1s4sq/7p
64P64LKiYrMtkI19xMxEcCfkCR+X56aqn+uFuIfDsqFCm3sBCG8EM4Zx95yhjx4V
t5H1t1qM0lpAhYMTyWPFvdGR6WI9YLAGFeUrirgKcQV8Um6Q0T24XBFFNsqs7f0Z
9mRBrDS5LzHK+aq8EVW/N5UhKvvmD7D2rV4191QpyXONJbzNlyUm5q9lJysSdOQa
v0liN1uRHIVxUAAwseWUmGWaC0s6KCm+Fw/Oc0EHadYPZzSptXs3EX4nDm4ts4R4
3JT2T1Lb+Zw94aqCc8BusaogOsmS7TuBUVxCow7W0WXZ2f979rcwiVWYys2hwdvp
J8a7QUzV1Y98vcyxCKFAHUdNS5T9iR8ZLbCnAfXmMkuuvYmkQft0/l8z0OfyomkS
cdkh5tH5GH2HjzR4EsFrm9G/OAXOnvB/zD/OH2EbpPcBPfql8+UXG8MpdGbT49XM
j42yCNk+MzVEqQpsyoP/OHvI5fJ8BXSg6EEqOWaakBPjsLVX0GAoMiDCDqTvqE2T
l1wFb7czCiQMH5/sjiJUrSloQZIaOgU2sJXckZof/YUJY786jp8dNn7+T4JFA+/u
pmeaM1p8h9KOLOjt6e4LUGvjyIjqcNbDdyccSffBXKRHVypckkqinRBgSdY5+8t6
WVcVwuV1ZX/zxj16gqSIfiAoSBj85+mv7iETjSX7nb+C3Drg9dEyXsBpRz3TH4xS
PVRYp2rk3OoAFA/Uj4M+KInbmCVy//U5ApngEPVNr6Wndo/sMBu3qqsS17nZlfMz
g1lkT2D0iD7GWmsm7YTFpZwlfjJ39BkXzkRgkhGMOFx/DX/098R66KSqJpTXljUg
HohmflWi4pqXIji/kdSX47N1gqo8HFoLr84mffZ1M9vMULI3Vsl6vEhi2Lc0zpW9
bVpTYWQSnSewTp/rXcUdjK9QlQjjzxzR6zxC2ly4juMlALDlfUsMpzZ9Qm6Av6wW
XzbCt0MCJ6RR010e4W01UkCSNvGwLjHAnhWivF7lVQKPelmMXDgxn+o0Ab8hpAJx
c2y3N1xCbM4M42uhKrtCuCRx+hZVXb/f8l4n4ZwR7ECyivlfdS7RWqm3fxJ26TT1
kR8wi01z+12wB1AQV4snsZWCjXujNcTXpG3K6EUkM1sEu89aaljPlmv/KTA/8/Sc
6+Mx5Zn5HViJf+LERtAUXbm0o8WXsKd8sVe6t0avdBreAtfscDekGBcImAtiOtyQ
lDwmuA0zpu0Ok+ytn5F/G6nabfd4L43L2VjRZHW59v3cIk7GzfE5dcORCQlBpn3Q
iH9gwF+M8HEVx6bWQr773IPNGjXsiSge9RRsjE7YbB9ujtrc5WS5WTVVbOVNqPa1
SOsC3dDw7wYc47+dgM+6FM/m+QQcacctKR9uxJ4jmk5hwtMeXFY6Jvplv5qw8B4J
gCQO9q5BIFo/2oOh2Umn7ruVLdVvsf2BMDEvcpPHL0NLA1hC0VI3FxMeBHmyG6g7
EFWg+4jRPD+WVwsGvTMyyZAy4EnwBS179ChxG/r19UWy+dtsOaCmDov80Gseu8mb
1x9wMrOz2xmSPSPhEhf287Udoyd5QEYpaO0m/jopc+IcwN8jnicnlQ17I2LY3b7Q
QiaaQV3Asl0hFnIJTQ17iF5QoDHTWHNYGZHPQ4QhG6m3+fJ+wBHDrqZXAs1+XyPy
jVLqAwRkf0OJaqEQA6vZws0MobLrX6e9G8LvTSs5enHSPBwefAb4zF4MMkafuDmq
Vvyd9Sh3YWvRl7/wLcmZkQO6+V7BbeDFoPgUncQyBTh0xpCR75NsS6SWAe1cGEs2
7vD3Hwbvb1SHSsuf+VIu72KOrR+aeTRGelpsmc3/+A+MS0VY2qcRcxrt9ga2sCgA
13dtptMrWm025elwYORMzynq94c0QAZewvbzLGbE+6dkEbk1vOc+WqYlXsBz58Y4
ZPZ0mIi2Fs7QkGeN5kCttspu3/kM89ZBEaNhwAL0TfaPiN5EBjWia4bP5xQNlJLa
U9jcUgSFgLA28zxYxx2SyxAOAUd/FkezoFSgVjisXzhLfOtvhP4lXb+7bsdHqEcy
iwf/X7OYdoHSuxkfWhiw1M/tX/nC8A6t8Vg9J7/PBfkpCydIJUF73ARBTrbiH0Ld
5DB5XsVK8k/2QufY3ohbXlJEmyBmOrngYbk59xdXnzttH9xJrG3Et9aK8GTMVa+u
4Z0QY5DqxfjVCxmzgM0nyx2GJRQPYf4SAGwgGHQRqpMSCWJRhRvwYmJYkJs1yw35
OQi8d0jpEdVHXUxA6/3OzI9Mz/Glg9+s7n1/nTJayFAwPMl+6B4iJhc9jKf6AZ27
JI5t7Si1B0fQYLbZ9oiRae2Hgp8FIyxJWPwzInbBUrVVZCdeaHQUguMCQkzJRiVz
gyvkPlKZERQJJ3zvE/bhelH6hLmv+YsOMEMJiWV7dbLo5vQjLy/PNevvYEUE29LA
1OY+dhMBo9ssLxW3DJEmRJtTBbdavMQSdWe1/mCwXQEjOv+P/VGCwoq6BUOGeMCI
p+X3WzTUVyLJuoLMJFDPWeUAqGdXIe5E1QlAc95YLpTG7gw9ZKdh5RkqSX46eXHS
CvblfLFN2mDMWFwsHoYDurL9q0tXyCcpLSNBZ0qPZrQVh4erZEC4LLKmnZxeki4r
kByO+UAMzWZhF5Q+VoyBox+geKxslovI+w+jaYlZ7f0LLaKT0rzMITV8+CNiT9J8
lyAXNm3bIB+kyg8X+b9qDKeK8X6DulIg+5MapCADhga8404nwEloKv81++IxnFQV
s41yUt45sDjv6O0ik/ziEpjDHg+HGchgnDV7iKJyNgur20zluqtII+tAngOJOrXn
W0+yooI7QZZDjrM2le1yIASql0HT1xeTBXvOsvoxoIvcC1Wgrb/kbOBEZmApkqJ+
eKSl+V5WuVpPIPWEbPLzaxLe8WsTBpZnaVSuLff/+RSlHrQJRGS6+CHnMXooQtmR
MDPVtPieSB7apOjXePR+lDjZ+e/nurcRooKvNSqXHA8wQBhj97vDyz0bCXAHTR1V
QXyl4O+9JyIIVHDERtoyFjkKpuqnINQ0Dg3YOQxe0IIHVmWbnYeDtT54wU+rgMiT
N1YWP9dkMw7DRq0TRHZR+kdoKyXOWuKXBaUfhoLQTPAP6b08t61uBX93fym52ZY8
jQHF7G8A4XKC7reT79V09M+nPsaMpdIm9WHti7U+R6uxSbqQIC8OTiBN+7J077zp
KkXG66EV4Eny8n3M+zUc6Y5KAdH5XtaGONCgflUQM0ivVh0dypCUHrcba4LhPAhR
q2BEhQ3fDVRyqZV6SceLRXY7F6IkV1IEmZeNZPVq5/BE2vlTQRjmWTedyYtWRTtS
9VxYBrD+SxDdoa8Nd8gXpj1wXzI5nrVNsd3ERzUIwYN7IlpNF3C0r73uye6jcylC
fMzblK0TySkgoVr7VeHVv18L3whBBrD6fhGrsNOx+4uDw641DqUNQST6lu3iVqfR
P8CtVsd6NX88q+rGNH0uFzf2svzEgo73bQzJU9727cL+uLgkZ9O2pVZypHsftuUC
6Ct4ALfKZuV2KpCAClYnvdO4dwIsuyNy4ilFJZgBDjxiBssK/4Ve2ky1O2id9Abf
/nmkLrhHh7cTY0mPwHTSNnid1Ul83eW7XgcfvpJ7AgIrVRfalhY+sxyhQRe7bHH5
6d7fSpX4N0a2HdyGIX3qDpswM2XtyGInOtg4ELa7LsJiYgyuzYWurzcGlV1TCyQD
Q5KflabDjqb/jO/c6ISznabSHSxcARTP1eECLmS6QFQ/MO09YzSZ8o/Yz/uQr4y0
PEP5cmGPhoDkt/zTqT1nXCBM19zaqPIEGCsqvu9AVMLCb4+AP9A+VP6GUfOW+dUR
21L705T1Ju0TUnjPhyq7dM1euL4qi2on28ZkvOizMwvOTn+h11Eax6ECZdxsfsVG
/KKkinc6DeqiwNPmG5TEWU5K4ytYYhxyD2i83hT+ofLAfPCjkFuVuf7/u5dmlTNW
JiHeIb3Xgdw5NLvAVaGoikt18+ZyVF/XXxbWGk4p2/QBipDVDRJHRZIKovpjWtP7
A/Cco7Vd9UaTcydvZ40mxbugi/Ebcpfr1nKTN9tcyowWt7KIjGvmVAzXjMtrAJ3B
HDUZvTmpCA2JuOYekZb1dw5tS5MgxPedpm/xo5djoOzwBkFJv9JhQ+vKWyekf01J
AunOOEXBVefJClYhq5kknMRhoHeQUhlbB0Ai+slD489T4x5RINkLL1VL/gJseeUm
tDlR5EBVcaR/B+/h+XB4MhY4oxMNPkDI6456TiA6D0wEPfXKm/vg0FUnFHEvfhC/
O3t7KSnjinGdFON5dLhE73V6fNKlgnjz9YOGkRaHN9SqeC2jl7d5vBm1zxyvEnzy
CENRJ7L6cFuwogpd8pO+yMwuI9LtD+7vcSyQIV+POW6GQ/s97oR5nfOsRpJ/1Igv
/Qhby0Oc2bzHaAmybF54x2fZ+ZXU0bnzH/ZNruKXyU1d3KIdtFgEzy4CeNtGFil1
8VxtkX0Inu86zzC6aRCq1vtpF508lzUht3TklymG+8cwHppqS00pgavESv0QXuXH
cHGE2l3bCEmlEyWy254vkKToVPTCWkbSQiuM9g9DTHYdK00AzHcWS/925faCItxJ
Nmz00RiivR9b3sQEYFZUq3le64LOE6OHLpm9zSQONRPF3N9lLV8chuPbZ8bsGMz9
o2Hprdr2xB7lDVrtw3x33wpEa+Qg49tQ7oL0Etgx6Pb5R+2TTQxKBowGYpdmKlIQ
JI1ccBKCPX5Ipu8D7puQCAioxznVJ4dAc6QlyYrlm9eCSIlQi0D3oVzserdmE4Jq
f4jQQCXo/mwVQVlB+9ijz28YFxGkx9jiASsJDwLEQhiwy89P0L1YtbAMK20hl6x/
O+W4dZdbdE2BDHnwU9ShxM/yOshhPrNb+Sma16XLRetcKbmZb5oP/HzbSfiMozkr
efVvHi/O6dFNeu3LNc57sx95nG2zALm44rsfNOyWVjyL9zWBxXYIkghueydIJNOH
nvi2aS3a/YbqUgn5piZDlVpmN0RiNgLTEUwixrw4OPuWFGCuM+3j+fB6n0nU1H6Q
WvJI9WVDXfT/HP4No3Fihid5QW+2mNQSxJfTrl5qKY2UcnefHSNgcZibL2BDarN0
52KLaWXVaLnJ5ZcgDhz7B0lVcC0giySPlepklY7g3ZKI8Ip7Ps7uP8DPOf6j0mBQ
G5kQqYOS0UQzott+WNJisIjacHNrl/4M6Am67/RilS4aSaVjh7smTtS30PvwL15A
ax6ZTjaD7HfCdmxm5PQ44NK+EyoQkj4CKur4AA6FJDylodZlqOtgGC8rUCczQqeK
ZZp4dnhWypf/d750QnVDP56D2AR9JzNtBparjQTzHEtT7GTp/uEmgEpvCtDfjlqy
vR+Jc0U2KYwsOk4pH2jMiMgBo9baDMKHtYcHeiIrR2efWrGr+/2nKM4pWmJ2Gu3U
9Q9xDClgXq9cBLjHdA4x2s+R2+SyTToCIlEYBxDASN90Nql/kcaHxVfR6lGor88Y
9ShqDZ9cc1MTOoPW+5qV5IBRUJpYgji9OabIcDDizuFRY7WwpIVnX9h8mcr7bXqX
HBvTgi1XkfUOhapGlnoW9kcm9cHbJzF9gFkrbhkpbI+Bf0Klp1YYvJaFoqwKOpNl
u/KIBhj/kc3oHn5cucx9LeVrRSL2nujPTrtw4Yaw9HnOQdvnO6JVA7T6m5gIdm32
veMp2FZZMEx/Kn1d/c3TU4uhffLvyM9vRbtwM/pdGXZQD0Ud9Ui65vs4B+H6fGBT
JvYzdfej0RVdCLEmZUCj972H3HVVVpNrRnIZkeQUoPaUx0GKjE1v0DwdyAVjRZ20
NDINALP+0onzg8axWWsMsq95HHLo0fR74rNFV0TOsazoLiIqpDv/kTNIJbOUAm+I
q9g46KueFSKhFuHr3Y06zEPSNgE7ri96Jl6y994gao3RJZI0xO5eVGPDBj9PsDH5
Y7pJ/lLLDRMiUUxUD6ZoudKUKK3mHhV3vSWuvLhSiK2lWhSL/hXk8Odhe/WIBrxH
IfzWAmaLppzWPJ4zEzEM27j7G7q26SbDsSq8A89PPnNdZJ8yJejeJLqWYclmDMEf
DHwA1bkgtGPK5gY0A6Tz9x06e6NrpOp0N5TG+ak2VPG+1MVWumzfsU0Zmo9s3Lub
do6v2LLiBtU2ZwLQIKxyoPY3EugeF0Ztgxm9+qK0FZaT8TaFsZHXfO3O/+AS0Sc3
KxRTHD6bA9DN5dNMGFfZvVEkwbCjl08xtRulOQc2+Du+ibPyY1d1D7vcjbRHVhNW
xO5pbt1cyRAjiq0BUD2wLQLzECTP+EvY8tQF8MydJqzFJIkR+2kpGnY6u0C7oGT3
bz/cmNjS+bRcIZ/m0oVJ+w1bpGHg1vzo1DZ9CdvTa9W9n5MtVFM5qiMaG0ZeBVc8
tC9yRpF2CD1Si/WYa341GZLu0F9mcZLfyevVc/7zou9Ib6GdMwzUrh/ZMyO1yvVG
Ics7TqI3jDJWgeXUa74BRlzYQdDalteFq1p1bkki3ufqagp5q7bTtmTk7Vgmw+c+
N9H/3jrI13H6EIDHJ3a6VtvAq/SdbBjdy1lkja5PN5CVaaBb8oq73ov09GwGMoOU
EBtZ/yNbyiE0NNlu9tm2CA7U5EnKgeObxj4tW6CEv+bOHty7Ga73RfZOZhGb8NdX
NPYdtpL3gs5TqmQV2RqRLNCR8EFmJ+KfU8YNPd5tM4Vp2l+0LKLwHSXkEdXrlmrm
mS5DOxH0C0zLr+qbahshlOgjUCmHHI9mIibT5UG1CY+Qdo2My0N4rUZY0XeB1n5V
mQB025+Wm2AqfToNVqV4w2gCjhORWrLx0ZLuk+C9Jto85qcrW4xrhRT2/vIeqj6Y
g1u7NGkvDl+B6j1tz9W8vQHp37zB4/oZWiW5greMovS0dgGoXACBJhIWpkjx3+VB
X849qBrm1Id2YOziJyZqqEJOiGtt+SKmOSpp/fYi8vwhJCDiiY/ML3fHCllGNs4w
ZdPeFj3Wf3kua3z43UZL4/f43yuKaLxGISWJHa+H6rNWX4rMX6AoVz7yif7VHv+u
hlgUtiuMvDXge+Es/NZFBzwizodAoHSBi9Uo599rtVML62AYV15+vhYrFaYcBKd+
+h8PQ/dFFIOi5WCx1vVqyoofg7R8mHqw6minmJHzsNkcLu1KqlbRes3pmFbMpAyi
DToEG53ibbTavamcSIW52hL8hZbub+i1d0bqzlRfnlosnW7DirLWERFlsgrfKeSm
xJOdxX9M/6sNnovQBzK5nLmooUxTO1yVQPW09esJMTmpcwElMm5iwKwOiGKGARhC
jox6LaSyx5Ejpcd8iNhowxYkuVhdsgLcpzTPASJrHuVh/obOrGfZlX9wEuobOszv
3yGYH/Rlct2yvAd1ViRmDaeTZsz7FjOXjhjkszI1v+B9EKZ9xWjm1LDDNv2uLpu2
DUbjhsV9+v1fuM/ToQc+ghswaIplN0UWH8Lt2RUt41GaA/BOLkaqciJMTjSnpOdI
ciLBmQmO6AULizlykit9oJ9gBwDIWIpaeUpFi+cvCalK/wOzqkbWQqdSXKGlBthN
qoYeqDd59clyvrZrT2ZQG75XJbHJIDNg6p7NkXg2pFn+IEyA4WFzRV55gHxACedI
aiSrBVRECp8B931xBN5Rq0EAUZx0gCHBrcyJUyCIkLFBxP2fGZnAK6z5ifHOuzHN
Gr8P3MKCKJmCFR87Og5DsN1jwWTTJF+L16ddY5H0F1TBrO5OSFm3EXO80EN9OJiy
jRKdV3zC3Ki/x3udrIvmt4+s/3oTOfC6ASP/RyEGiAmHWeHBhCw0K5RMDk0Bf8Ye
dkb6AkTXzbI2Gq2vXqXsi2TLjrTegQzYxj1lsOx+ejJiZRXFgX3c03Q3AOtlqeli
waCHltrd5tZCZWGIw33/5wqwjXjMVBaF7bULn/0TWYBH2FFe8L1z83WXfprpPFmd
F3Nxl/X9RVpdk12ERTAqOP0tJ1w1DJLOQgvJcECxbImIBsU20bFPuxSFX7AEomE+
quhOsZKM2V2RWX1MSY9mK3TRA3zOtlKGv8r92+jHJGjQ60eJ4mAc4oknYSEm8xOj
u+BYbI9vV8Rg4ADdDycpcHoKpNsdyMNBIiEY9n0Og8kWXGTs6gPjm+XaEgcfcKFU
jX7EBgPU0hSwzntFCE++OTk41rRZCN4eyuvCZwyyMkQVpV3VUP7mlSF4u5+5xLmt
x8pTYU5yXTwmoODW8bK5kwCiVnchIWAdIyb+dDm9UdyOpmD28sSUsC0Z7/3SOFHm
ZWmuxD6IBIg8JnSqlGneJmgjypVV27Mzy/i0HFeq+dsWvgHZ5Jn6w6pNDogqSUma
S2H8utH7ygsw4h1GY8sHzsk4Q1NGMJTUn5Z4QMIp4N1PBNxUiaGf22FL9mqIIuMo
Pj01m3Qby9gSAAi4Vdp7uUM5o3CupCi+RS71gZLaDAu39EJUdSYBggVxF+YaJVRM
JcU8la7O2S4H/MG26Nddy5pTnVuX+i4jj8wTgRXGrjCRQ/jRJ2YsgjpR300yjT14
qHlBzF9klOMrlt7m6j/hxV4Atl7HoBHRiJVgFlynWU8SfrmX6WDCvt9eI2+L+DWl
hZfHCYWoIqLLxXv3fgQnB8D7mL236+HQArQ1eNQN+2DsXvrQixOlDLk+K6M/qXV2
LqD3o454DE64xoACpM3A7S72Fe0Xhn3SkSFtZBCYvAbmcvlteZaAtWsgl7UjlioI
K/2ZsG1pqhlPKC9IcThyus4siWegSRWTYhW+fzOkBkrjwB2+3Fzyu6KSs2uUKNE3
MelgzMX9wznbfEMzPiWTnYO3I3nWHzV/JKQHaojuv9ZaWx6P5SFjb4w+OPACrebC
7sEzlNRWQcEb0pKvNxT4Hp72+FVJXMZkUQazIzgUkfC+DX5n1Md0CvDiycvwP/cQ
4P9ZnJeqDmlYmQmDP9EjbbqItk2Ew0BdyLK4PoQZGHZGwJ/ZX3J0sBLXoZM2+kRc
WqR59RlBixFN/i/dxziiMk1TR0Cgex1C+0bSrOJf0YhFgqPG4fiBrILWoyI+doGF
JSiPqvo4EJ6PB1YtXMzbDx7rbnuZ04XOn0w0CTcWhapQfNv8y1I4+v/boXshSgSQ
6NZqtCEfJeiSBw2lHtgI9DsM5VvYC/Pct50QCXfGrzEq+XYqITurs2Egv62jNT6a
WPX89qGtmSCtvv7lD3RdZdNqqSzch9fCSQdc8TnDTTdAHhhh5kMihOwVrB1FtbNV
9kmrCTxGLI9kTcUJGoiTmRoOYaCtUGXSvyVS9kCx3DCXqB1fJDgIMxqHKZ4ImTiv
7uGIUxvOJQlTVL65g2cUxveF/hs02G3XRkHpjVaidoB8pYftss2xSdxRQDlpDa5t
DLZQF7ZXqHlEBrEiCcRU2Ke2dGfPIm1SyXcNm8wFLoXS1aS17n08qcGf8KL+bhJs
J68BeuQgWI+KX7piSQJi6pxU0c+EBtYvRcjuBPrQZP86SROF/TAMAC2oimM/uUrI
7R9f9vQO3VFk+WSDJPyxyxeI8UI9zGxJzzfO/U4zpUYzwEd/fbOWnoCr7G2y0Hx/
t6jVOpf0Syb94wK7j4dYVIXsWhKiZxDO1RnqzgdumGWie7eqL9jFDdQqXVmt+Cj9
fOlqQxxNWttNQWtX5bbF1djnL6oaGtIoPPNqMw+b7fVA6rN7FzIX7o7JB0CoLitJ
ADKuYMZYQAQO1cxdlxaWTgrCYu9PgasD5ONe/U7lUfhdYU6uv0PwpRLefJBxB0af
eeDtEglPqVrZR3oHn27K6eRoB/MsGLC9CTK7Ov0x/EMqopBlkrj2X/yUDhsrcByw
o9UcB9x1EJh86Damp1rnGXYfH0MlCUW2+T8LPvmZlwC2k1ANyl4+HgP+3DxurRnU
cgKhhSafvjNM2HBA6N7F2e3FAeRWwNDp8h3atblxf2YIKqmVMBDe/tLXAAHzyoFi
pE59Hzc3q/ZHhs1IPNN08v+SFNb1Lq0o3/BjzcDQzE9kbrojYb1SGTaXrC8XFZF8
GxSe68clDKP1n6wtrIQh1R6XWun4gPjrhM78wyOm4ERIPwt04U5XYPU+ouEDiPVQ
Flnaip9A9OBp/SseUuUh1exlpYGCxCVH2FZvDFWcgGXCq4kv6TpTHacjYS2gWHXg
P6uTfG6JsE4Za0VjT/Iu7lcVvM4xxw1W6tC/5VDzSGjk7jImchjyJylt7c0u/gsq
oq3yiLitEgm77eSH2MNNgR+5XQ6HG7e0VjiXr1ZNjdwb75qU2zpYtviStmEXYCOl
16tn0Sd/vA4NOvcZ1RA7dTbGiD/UwLG6iDLrf2XEWLn94wcIn4qzncx//wD96Dvs
z0BfPgjidfhquRRX31OS1f4Oi3qg7L1Jk1D0w53sYpmQu+XtnUyf5Sykou7nNX1d
zmP/JDbSQ8sPD5PqM77nMkhJSpy4Q/4FGfU36AGDgva87UeAmMMLPfBOLnKPHCws
Z2wbYfjFdQsim6Q+sU22nxbOH55CwZLShrJzsJ3zt+eiK493dhXqhd5cK1S15vti
bW9KLI/zhPuecfPlCoxYo36E9RR4AXN0+1JFIUirbAmKUYS24r4pI+eelXphkMcU
5QQGsqiywL+hPot0mCzZPU+SWBXTJqjEAzTl73WSWnOeEvimj+bwJIASsNpdaXZD
rzvWMYeAF9dc1IBdRDFRHF3f4TqLwStsBpjlnfdyBGmxOhP72reLkkTpYK+EJYQg
mTOLcDQolo8CcfI/IzlmPkAQqHG8QK00c/7zw7P1m9YpIblyeWTnU5A4udEAxIwa
hLNtyP846oXO1ZMqMHB3EGpBNDrNs7CaXH1J32KXF/e6rIuliUog26SQFOA7pK77
ffUgsUaFkEAfqZR1efljvNYf/RPFQ7PTfQE2647KV2tT4RAo0doe3Zei/8+/pZLN
3QFwPcnk8JWbpPHflsxUroiEV0gnTcO7gdEGV4T/Or/oBbjCkexir5jJQ2A36Bg+
pBTilyXIA+srDMIhWK6BjSUsx4jb2vuuVOwJuWavjPeCsW8sGG49D0WArNNrLNXI
QC1fz3gyfsnVLKQutr+S6IXksFDQabbZ8RrErcxxaV1cns+EKXKgnYuftLh21Bq7
Xv0rmg84n/PY4VvVH9twKQiyiRsBBmAg4Thqc/nTz402NTVkafVoCwTTT42QndyY
8hRXktabkwzBx/gmqna/W54e+J2blyxy/hJuwSa/P3FlLq1FBMhAYvUKhflLZpDG
jerQBghhxi3aixULi8GdxS1P/rzTx7t0fRK7PFcuS/I9m/TNIpsCqA/+4lO/NZR0
tFqRPCTaY1IBWWZmm4z3qzH55/rxecqocmPJkwvfgWCdD3ky1EofSapoPINsGA4c
jQet1vIjy2xcPave8/VnLS+eUmG7gbxWS1tPqUzgkdpRfctuZhCzG4BOnZJuKN6/
lT3uE/vKvihFLrHTQI4L9iSKmO1C5bjYcUcbtQi/IZ89iTack6K+kjZeBd3NrJcu
TlgPZ0AvP+5ZZ9xCLYo2wxcM6sWaXMZ5QmpZ665euKLxuP9X5+rXWlfNIYkeSgGd
olQcQfsZ2QL54EWZKmZb/PwFtjlFT2JN+4HaW2wnFsHsu6tUFwcsAhhnatmj5nxV
iphnbaHtC0tmt4RSejcjf+ijJecSLIa6qSAJRTI4cebYpxYKdCkpTHz/42RsdzHI
Su4OPuAGpOIye2D34EUmP40iRcFp7VNp0BAuTmzdTM3e5kK8MJyEqq62/foO+E3o
i57TLki9lhe097MSy95O4H8UHVdcl+ckATmAa9tTkhg4HWJrcy/OIfTDejeEqQ3d
Abf8LiBZ1Kc3OQ/f236uaOC8XjHq7l7arsFl9Em1i83Pt0tdb/jQtEJ808d02DCa
cYAdLvy/fdQCbubEnfMbijcFya+4Kz40K7zET27lbLr4PPOjmnM1bxzCYOw9wCzY
QqyhoDQdeVJbLzrBFecsdHLEZGD7fnyDPM1YpM6IMjFCLk3Zay2CVuExTwqvPDwm
COpeeCmGXxKQKZuiRhkD2B9hfWHEhJIojCKs9aqHYkxyWyOf9ZMas4lHZNiWhHnL
YvWFe25GixoEmu7cZTfFW+GsVtl5jtaimZwW2zbtj9PwCrlipCkcezExGRj/NawB
a55RLPEO6VrEcTuDJpOIcbJtZv6ojoSs2wDz5HH9pMCkXF+/0JangVwu1NUemE9p
1CJJ/yOjVKBg+McfnBqNK7qs+9/GnITDyPXszFA1j5r0A7N/DPKJUh+XMe7rNm0E
1NfQMaqy2Yxlbq+Pw/BBffxVlFhVNkGtCsjuFlnnP4P6hSuYsdbRAmLB1uB6MZug
GdBFoqUa9F5sBtBBOiz5zrg50BUi6CmWyyYilT29JP/+2X5tgf5n5aA5tdozDqA3
KiB5I52WS8Tq1uvbN6KtwldMzuO3AFa2tOcCUOtrFJpYYAF3sCaib5FoYbW6WEM8
o9ABD/Zoc1RSuYw6O/RoTSmq03g/jtYGmcTuJSEKFg28i/kdc9pYoqQGdSSNHcXP
bJIfFtTph01XurF6aTiLXZfn9BChBMeBo5uyERg3eWD7vrZiUrNFrpBeIaSywC5L
NROFiJEv7weqYmjisFdTQOGu21xufmpRlAotw9fH4IGUVGyXmZHTGjND/a7/fAbJ
k0HrK0FXIGZOGDgVUCS9+gVCMdPI+gz7HHWZkX7oTuSY5rh1zfV+HLkhbqu0xCt9
VlR1sRjW7Vu7lQAZhRjdDUk+mXxo6Z4z3gj/E5afBetNb4E78F5TiqEPrBGz2+Hq
1iVpRlLEs6R/uP4kf+2f6KX0mdll4hSD1e9WKmQilLcjfSx6L8PY5tRFlRuqsygE
Q4BeGjyBzQEUWrpUVQCKrPQEv/IGD2YQlhvz6BFi862oeoc99fHj3V7OvJHCQso9
AL5XU6Vzx74snOdLoAJdGdoqnT1IdzHtYmBnrWZmXKaJwsawyjJ4jyxc0K4ONz5Q
bitdh5n+NEclybI+b1KfDIWOm6zQBKgGaoNuFFPwPo4KEdnSOG/S6k0MIF/je3qk
K0Y7paSYrulocvvVENM6UWroMNzZKc77VItrvBKsVTJKi2rrecUNEaVf6MJ0qWIk
tDgohLPeWXZhjP3sAJPUN3adecZptKwUx337mngEV1FAjU6YcQeJ0rWLN4mqrySr
1JyBZ+SD2DlvtfRPPWsR+KiazdugXWB2TRaVVu0XY7jwESpFsz3EMR9fur4VAnXf
THBOqodsDTg/RUhDPk0CV082PlaDYEb3F5/OLOnq/6dmbSu47Hf5cXgB+Nvf/7Ys
Pgl5WvpVMDcnk21OWDfl2iqC11ASGrjMycYrKivCnBFRkP9UYX1mI/Z+KYcu4Jy+
kg4MxIWldl6mUB4+Cjrf8VGnHbUycyk2ufwgEaQbhtsgYLMTAfz3mWa+dls/Z++N
SfFzNW/3iPYWF0OfPcrcKHxHq7RwoNoK6CmFLbJJmYEIWzNPeZoRidvVSRfPtUBd
0PeXZB3w+aSjy4sx2alVT98EU9zfEyfQheIwK7TUITmaf3snx5wxL260AXYaE4FI
vI/qZTWo3uahZtT59VladyUjVvU3kVIU2l54nyhpy8RjoGdFKcvH6VVgl7s3fYbX
H/Cq4vAt5guLYV0Aexz/QMaxVx51JDXY22hR9Dxy+YcZZqeTIALrKwCxA/gzA8rK
Drx9RidATEhVXZSsM0QR50WnZvOtx658uX2x56JMmxDDk1zV+xEq+pYitTy0kPmL
tHV3oGN4j/ofnYsuPD5vvGuW85GVaCwys6LEyvBAprv8rw4nFWNPh1777yAclRPa
acWng6yYedH/2FAXfEgVa1rm/QsRNWqvtIBZVqvPmA9Xd9N15xEJ9L0E1arSs3NN
EVUcXKvFA9S/9j8t7SIqXjkJbw+9rd1sBaUiVHt8CsbgI/VK3DSj1oNjxPYNxPiJ
1HDrx69fFpO3zq1fgNJSwVLGsKCXVhuK0pfgIN3sldHWpRUG7l0mgQnP8/9oH16D
4FEHU5zOs0QJsAMsdsE8qlRIIuLa994iN91xw8NOE97//JY94IXWJjxjE/eIsn6G
1KR/6DxdKyZ/z8ogjjQWUIztQFed93NX41YhsRh3NjYNJ/DzV9Q8olHODP5/0pRK
SFTRXqJQuiGOPGZ095c5IPcbbACZ5/KVkPrUvNJ3+A1AFYQyqCnGcgQZLmwCNznt
QXv15t2i1KBuQezJncyHrsE/mhbumtEoXYkMy4K72ORZmAwF/kDaRQ2vG2vpYf/+
sas9djB4tFLDvA6kJPlcj12qXwVQ/Y/10WNb81QDBnSwafpVDGcc2Vcdry4nCTeW
C8a5JAJg2OssUqi/dMhijnEI2yU8nLjz67W8OV+WzSVldBgrC8TxN1D+iR5BzrpY
ierERgj5qLJWqs9G5oCVSIBYsAjlehh+NyBrctTdf80BYNpmFbUBuzSMItRIakJR
vtWfCZY2qYxgeStgXDyTu2skUVgHkWQP7SmM4Oh63XH682ZTbyW6BXJnFzb3p3mC
b5DSGJlrlb/utDDJMc1++nx866INHL1XOF94hnHsiYK9PDLgkQbn4q5+ecPrHfWF
OO2j1ludkQWwel+zxrNEuSliGKUFx/UPl6RRPQUFgyQG6qDHzd989C7+ftd6VT32
0tJEZsJbu6yraCKeecakD4u4Yyw0G9fNR/WUTwiyJpjYB10o0yRj0mOkuD7w6gVk
GVbvCaz0nS5vlqgqx/pK+nq4QJwOpyrX96uPHpMTRRtPNqQviX2PLWF5YdBHO8ac
BOJ7Vw7VX3KwTHEaH1x11CWfd+tqz5LmhR7T+/FioHd2W6efpDmRtrahEuanC8sy
DLHwn1SR7m3OP2uQcay6cpVI6iqbSkOhX1MGlG0xbHyqYeXiZ00dtAyScEnAwDYK
bPDZkCXEWWj32rW5UmuILJzg8FMyXsCPIPf+lBFpIkiRvQm0X7+l6HwcuQ9ktnfn
UCZ+QVAPN1lBiISWyCKT3fK08oZ/UosxTaJ1Xbx0rmB9KSpUpVL2glkdlnZRgffT
VcPGJxPJyMpd3DCaRlHxa/A8XE1iEnbAl1hLEPNb4wNxueANAi+6NlkNrSCfjozT
EWq2uijhXm0gdOAJ6neh3XNpxqPFMMEjIB7+DnX4UPA43cfPAySztJe97S5BrHSd
/kkwJhIRZqvGfAN7G9azIv39pQvs5hEg1t/fdZ+HJ8jdrSdoVou5LIiaHx12KS1f
CGSheB2um4aW1JxjtWT/KrJ5o3YcCk2ddAuejhjYfjSuqXdXtF6+i5LV7ccqZcua
RBPTd0LUuGRtC2+xdom4bVcOR1nzvhvZG4eMx/1LF7BvjFvHrDAkAh0P2CGu1+oe
V1ZwD9aG6ivvTOQfLmyq5z0AE/TL/DokGZaA3/fTu07FBbscKEZB3AAOEA6ca6Eb
hdcNZ7jSHuR31a8aPnzd/bPWg12MQBh1x7txOO5cb7LG2dbQnA/OPw2ZKYnR+94p
bmX7PoBj8Y+q+YAEejpYXj43XBfIZP0Y4gLIfzwUwnV9hY7lEHmgz9Z/iy77pPxJ
u9ScrL5jkc0hz6EgDo4VkOorKEpjmAGZTD+q+XLFkT2AdYebSL8KHQXB91mxqoo4
nYAV6o3MYlFjngYRwtkkFgmH8O0XDdbrkm9lrLqRkfuxqIaVunyRfSdEiWI+foZ6
OS1jJhn/PSIQxVKPdqj1FpkzAu4ce5btVJPohpb4aeOUF/ueepMrxulVlqc5zaXg
Kza2NUYKPgYMo7qgoz9x16mJXv5+D/dz6TrYYv90eZTBkz6HByKCct+n4327fvv0
DC4jfL1tO9kCl9S5V1yXUIRQBfhq8pFWFZ0TsGyCUoU5jGEWiMw8jgx6nvL/EAj0
zXM8urvnX+I2WaIYi78MvJfHpkf49yKE2Fwqo/sp2tIlpdAZwNJfeMokgSur3tYM
tuJryKpthFrtnRoe3Q5Vh4Tlrbbm030FzbH0HLhsLCZaqHgo7t8+BptVWfKk8zCN
dAGxSDwUvTkwkLRtbrOuUI4fFB6ZPJIiBlZo/bdmpVR8dc902htLv5pXWthf5lHr
VIACxCqmMOy2RUcdM1LYCU3gjEdLB/QWZ143CEDfgCczboUyP1CZm+bKotnag7Dz
436oM5u1qlNJoJc5aWEcZ1I7wc3R1c1W31nCUT17rcAJPdEpURsWUeMg7zC8u8m9
nBqk9M3GeZMiY5jFnxMqgq1P46seqbSHaNUnQqmwECrwqCsO1MMTSDHBkQOxMD+/
lEzH6f1Gf1OMMrnKGqNmmZnIAl5SESidZxGzzOkamHMY36AXZZ4HdCx6QsmrOfPq
zovQG5h7Mby+UuMVeHe6FyHacJ7QI6ntPBng2pqcuXzopwQOnrmBRTbtO2wOgv0s
iWLkmuGeAkdks6Im3MMAl7svPcwkL9H8z2Ws98dC7VkNIZfw0pkD1BC2N4pdPxfO
TUDnO/9lBvGLzZzijZrYRN4stc/lxvt+0UuSzg9/qMKUPHiKFHIdTIq9a0SA3t1Z
gTytuhmda4VzzE98Lw7vSroJwhYx7lBXM2rIVqlld4oHYYbr8GsZ/eOPRNwOUajY
c5edFc26Bql2/i37lwMrCWD5UQdAMndSKmQX6RMdLjiAtfoXtyLlYVHgPcy2ak9Y
gaM9pAcwTbcZaCvOfQTGrAizTA7PHLXfPziNrh16B1oQYB8z2YWA0zw/iJayf7Qd
LiKtCsakFH+gZJlxiVIVse77BUMgfOiACJ5ruRgXTIyjVdLBSWut9YI6rhNiR2E/
JDHs1wEUsTc2bQ93JDOSKsluDCZSXZG+4oJMDlKqk4/TDjrOqymR4FLzP7dBJsnj
eYwoQa8SAGOpkBZFFQncTs9HAFfF5czzW8D0wt1B/QtBggZyoBhvcBdpcMAwHMJ9
ouYfcUoYzzbwCtvIQpba4l9SRHnIc7qXEVh5WQBzniWhk3G2pYjcN1hKI92Bi0X8
KOeGVHtSrBAYsrkGd22dtMr+C6+yxcDhFZ1RvnSV3fzX77O/ahTxjVlkzRjuAH7s
vzEpVdkBrnJDgdxtjyDNGTt9UsWHFGUpFjfp8qSA/W5aWB63+i2FZT3p/V5NmiNB
hMezFBMKmLZO+AoWowcxW0fosE2HvCl/mJf0uoz9x3HoCFbYK/7pXrSFgoeYYTrt
wjyRn9f4xSe50TNEoakNtuEZBZfOnwu7gIrBZhqYaNQTXdrveke2gjoYxTWE0+1n
NWRtj3H6dlVTebomuZfdqKX03rM0PUDmxyBZ9s6F/L3SbQBFKeHKxVil8rcChJSr
5UavJvMV2x0HsRf/zaYzc3Z+xTvLQ2HDNNyhwLA/0TQfYg+Nlk/WUa2yOfXxJQhf
SxoR/jsGLEyDM7OBroloIp1vI+KQUrm8OICTM+6tqUg43VPUQlzPXfFKoY6HnQQH
pfDdGk/Cfv+FmatAZ+YZee+VG6Ii5Mn1lKXWu4BSRHO8Xm3ybgGeWun/CEbV2dlm
lXxIFnFGoBfAfhdk9eAE0rlcP7YtJTzXC/KB4S5a5lOCH7Of6Px8/gleexzGnoIi
Sf7UYsZ5Tq6Z1BQ4OCt4XfvCiOWU/lEt3txcFPt/1AEkYz1NOAANIsK+d4v7lt0+
i0qWhFmV/LjDWClGBxW0ITWR7ftsQy6EcQVS1MqXsd3AB95QJPmhY/EGHJ1v76KN
ulcB7S3jxhWpAmYytpGCCAM7BW9aq6nTBrjLK/LG3nfQHMIOauNmtmM57Ica49oa
IJk8poG3yDPDq3QXSDIo8PwfuwgBkgpnoLDcy5DDg0tGq4m3qjBInZGzLmKlb9ZW
sJCV/JP58Z09G6FVAyL202HV2z49oV5f1MqOxm3yM8vBhMIJ7xb9eBAyC7NitiG6
QMCkHEfcUlPPR6u/1maN1LmJ/Ljp6s4Ajwx9eIe/GSs7XU71nVIyDznPyou5ZZCz
K0fDsSN77B/pvl+3vqDmo5EUpRhBhZTs5JhnEUmMwxIvom9LlbcjfJWVBmvur07R
4r9ZsO6XN3O4q5+ptgUI1NqyjaGJaZyx+f9xoTaaV/KooTvjbwu32LSppeKfeXNe
g+pd7TNzTtXIIKRcRTrOpLHDP+RaU899iSY3nu+SyVXm+kWkdrjaRIFPX+GE50Df
oFEj4goz10ZHKZvb31h3+RqG+wODOJYqOY9Ubgm5EltNJ2qOyZPxh+BIujal7Pdi
RLdkSulHUqC87SXsu5iwnFSJq+HeomVZmakira6fBqgac+vyEw+Im7hINSwvk0Ax
gLd8tHYHyTAVguLYaqyNx2osA+kHQgNY0zG79ZN6L0h7jUK8rYDoQhvfZyb78vg8
kni8O+Qh8x0AwmvCEtKPw51sqT+ouvoNcUDqFAYIXJOq6QWRHMbLzdlOLMb4DUnn
b5SGJGL6afvR6s7vujrn7aLn16Ug4zjK6jhFIu9raoJYUyr7aDYBaDl0w3WNSj+9
S4p+Ip9DUhVr91KWkYHuxowHP1QUKgOE1ND2xcX2sfcOvDOuiyJVr2+JpuREU4iA
SeC7GdTktwRDcf+Wpu4W8JWcq0jRi8o4r0n0uVExNCvD+qAyAWD8BZUK3X64U246
nJNhPZqQLHF3dgcPfUcIGI4WkCSuMu30qjhicIIZM0O4uyEOtVEhV5vEd5VXLOCb
1YlgACSOY74ESr2d7iMm3YQo/HGZuQiqGa3AljMD0/5puosGq5UoGtzsmFkW85ru
EXYnNbSjEYWUIKniSGb1et7javzTwrBPX3weU3tK96oHdZA5jspg/+jmE4RTSQ9G
zrJT+jhg0te+jVF1C7i51wQ7uqj+SUvesWrxeHGTOmBmT6XQCWb1HQ80P1OE+AX7
Wmawlyk/RVLA9BvMF+PdlcHNTwAniWn8ReUOrvpRP3Ip+Uv0sD2JiAbWRpGlhjAn
i94I1yoofpb4MJSxv+RUfrbn9/0BqjdvxmEQ2xdfgMHRtwhJmt/65czwIUgvPLCk
3nNCo5FJ/j5bBBdFsM+ScjfE7wRprWWhBeDXi8bgAu/v2WSebEzBaD86G4JcMxoH
fhqlkHDy52zW+7yHXdIbojuY5MiR0t5JJ7iJ5TJl4m75oBB07wu+dljJGpZRipaF
g8LNPNTPfUXOrNW8dVIwqu2aI13qMEMaR1xwCJsKTry20MMIcP0WRNPFZhODtX7j
DR5py4lybLRTbN+ON3JhqNCgI1zW+F/1vQS8VRdDZeSuObFa3Y0f6N9gc8cSnkVr
AqLZCv3oLyKi/malZSInpxkR6duP67QB9vabIcJAUL6QNujFtikxhJW7bfAhEgxq
g9VgCms45geQ4uGPvUyB/9O8O82lIQd1DcJIzhGsUGQ5uMgo0pmCWy22vx1MZaLJ
jQyo/uTHd7vtKotUhn0ppzsT5cy/QL30zYscTxoPFk25iCb2IAl+uUv6SQT7om/l
rTsbvG1fFyE4xlPTapIy63EN9xxo2pZcJKaDP299A/D8FFulfzZdJENTwqoQ9wnC
pq24xdKaDHxaGK+JPRLQZKe21TgaqGw/TuA8L+ddrinDI4xZcPeCnPZH/lL4r9Q/
S147VX5JIR4zr1eZ09JU5mLB63QFPog4F/ePHYz+oeR40rPauYqL8Ysi7huz/pqy
SLwWJszZW53g+S7uGJmxHzcy/a9ptLEA5eilr9MWRkV7o89DaSSbAzZCftXGiTfF
P46R5bRrNWds1eE5BD5/CEU0X9/nwVkwVPQqAYZ0InJ2IEXQTjxKL+rTccbBO5oe
96sdVvGeV7SeOlamS17tgpnwh2jHnMQAlswap4P0/fSMJeURQ3x6a3eTXYnlEDGW
xfzi1VZ+qgJwfHF8Q5iUzBwGKBNveNo1aRKY+RZdbo1uXnZ+SB0S3gCzXvj2guM/
y8osulw1xUwfpzrT4TlOSDXyfz2w6mV/LwI5eDADWTjuVGmaPb3YrKnHbZT2BAOD
YLJOygMHTJ/NF0NI1accBGuMdmdgmu+ryLZeYHRYVoqH/MPjKGj4KdfwYXBFzjMr
qkgQzWUau81swhbRO26FhuR0/1DvK9Gq8pTR4tt7pjozGGl5rLDshyqgzbdUxWyG
cPY9PSkCzO5g2IwoMo6iFV5Q4CzzyzRjFqYkGV9GafpeO4Zzpgp4uh7RP/jRvD/H
++5BI2sBaznkLBR3s6adqYF7Un3A2zOxBNTBmxi4NNtjLjBbqZWCQsN+5ENqTAoe
aNFc0HqhaFXnW9ZmmxDQzCOyrZTQRh2L+4AcwZ/u/SOMrxm8+sN7FYyT/OjFEbLh
+cFIdSdv4c9AAVvt6Nxxw+AahiEemfGu71ToPuXHC+oohq9MS+98P3Plo566v6I3
xEr6lGh6zmdechXNSpqi6oPpi8kFSEhGogCtulCpbjuHcGp9MiY3s7HqDZ1etNmP
X8Xs5016Y/MPZDz4wfXkeXC2rX3J6nvbINNmQ7RWyoSd6UND3p5v+E1vrekTAsnY
Ty7yoEp13VyIF5mmsoOY8Q9s5am6srmP7R6NocO6CgadRtYKZblzrEZwQE8un+i9
6j1pFB6zTMoojT6Rvo9kSgfcs2U3ugpLMKXR5cRRnP3/j/jVN/Q/4HCeA32HvgLb
OIINWDgv5mRdUpSFirTLkQJv72NckOTufMxglvReyp6GiLmp9ss/3xPfldFa6iPV
9U/Y749G6VheqOPKO5IodWY3ySGf3fayQKYCfPJAUXni6RARnyF0Bk/dehBkE8oz
/477HJg7k3e83AslFDAaY1lj5CRV1Wv9lxHKI9hid1S5k0vqFHdvNhYCNlR82bZ1
PJySXRvGxxNtbQ0XwWhsUoOkNlwFmS+6cSNn17AGpSiZdvJNFlD0CXRqv0hDbWwq
bkKoBQFH7HyyYx/pf80jTbiTzgt/zbOhEYqJlPJ+XrmFFwzl2jYimpVSAbVGPqUe
ywcXjS8n5DD9fXUsbAWW7K+xvcG+ZFQOQvgP282dTq0D3nSD8v8CKE+WcxsWPbKa
ZXv1wuC7AgY7RJxCXap6kCqkczmopBhqAaqPcN9/5KSaAXsPEvIBmiIemSOLJQTU
TazOJyHmdhwJcBWG1XCcVLDNYFwP7eqhEc0L5vDl1piqaaUIhjzlI42UZ1aRfbnF
ILmvJcHCNtr4iXfauVq36aXkkYCqnepXc9LV+G0fN6CpVbQPf9ut+fwB1qWx2Rvd
0WKaoLw2X3Q+/uJhtDmjB3F5Vbh2iEZWT5bClZFrj8wSrAS9px/YCYc1DfZf4oMI
Kh2ZDJvksgr919TlxdRlyrzeeiTxEBTpYH//PdxEWZjW3QG9/HoxlEjFrB7BIjwg
nFSt/3/Twong3RfsqxRogNjwH/N7+9yQFU6pMYTQbt0ZJNZGhsZ/y6ibiTdocJni
r7Yx6nRseuP//04vTsR36e/QU4n3bRAN0/0RNr2yZYD34iCE3WDUK9pgfFl3wdEX
hJkmJpDbUR5FLVUqC6JntCdcWC3MZRhSlzxSOx1GvW8E9TeuSnnLUGJacxDr7VNl
G4BWqv3ZtlwPZn0bBnAvlDCoMK6cUKpFXb6paoYlKDWmCmmlEMoCVCMBjpcpbSAs
3a1IG/NX5iGLs6FAiaJy+CF2BBEHSNZzPmV8jR8HcfdoYpGpZOIiArE/leoaf70y
NfyVc7kRXxuF7H9lbKLTD6g4BnW7mIj82ptigWouIcAixa/eyrzyUKEmXHKMf6dC
Qu0mYT7pmhFSpw/NcMkfQlup6KOuFnsswpz90sO72454ttwV9BVERHfFyDetUg0i
Ncxm3RYdSvT8LSCDGB+IWeBG0EHhGKeDvzHxokyALcbJE0+mU/Vk14eesQjXHoNp
x9NS4+Uo0yS56QCiyxNXWsxqbqEx+kmBdI8LUIQoxwETMoUg9BalN5GZSF1jkbM/
F86NeWAhImRc9tLqQr50aE1GyTgoL8z1cOILM55JVKAwDCcaPhjUJJcH+hwSo3gO
F+1bwfRZxP8nEVgonWzqhfqJcjK+gKA0tIDw57WMOOndibJA1LoPYKQz9mqxPCxk
ViXBHCDPIIEmWodtWmc4nFGC6rAHXiHPt8mv3JKSdXzkLXen6vLqsEQVvQ+c2RIl
740O0NXibNGfwe5L7sucLJfPFA80WSNxV0ej5+iPn512gYYFbBs88cgbCDSRKtk/
zvr0ZwHAl2pCEcDha8wN3mk351HW1n1Mw8GHfLXJa+b6ZQid06TZKbn0bOCBDhXi
cVR8jTXoorzTu8k5id2bf3T8rhHkS8FvIJVhn3nOmxT0jhaL09nRb9NaZvntioSM
TahXhF1U1GuzovEnHbBpkI0VvPa7RIzdED0A+6fiP6di/MMPp/jm7pr5w2rYP/Hx
gT6/VeXT5NwrF/rCOCK6GUvLBsB+7kvc7K3zWhbtijQreHf1QCRS8+2dEs1bIPdG
ozLrUarr5muiD30hmb9vix9ewLciiBoDyuKS9ePsN14Y7ssVDG42XJMNgtjfINT4
V0QwLP8mFsRKkNBA0kuOPfRAzdqhxBGX5L3pTBsnmA8CHDP/hbgWjgrpRpxU+AVW
FwAnTtyRK5s+EbdV/XY9cGmmDAgvAxbhO35lfmd4ElDOZ2uLP3Em3eh+i7mO88L4
iqG5k6mJ96q2ymnTUDigfYK5jJAQPLve2rSOS7pwfCT9+5VD8xqtqkc6A+pCohre
Dr0pwc/H4P2eXbzKn1SxG7SS5AiuunV5Hgrm1m4JlQw4H0Y9GqYGK6tn8gZ3cu4s
CX7Ok8hvVv3qm8vQma+sfl//+Zlo+5sFsbTJ6i4rfFsiZTxVyU3nSeMaFTG/+CAy
Ulq2DIjqLwX8HOat5HF8tiICk4y+Bbj9Sti/ML/LXRdfEr9TyrZCbboUW5xcHfnq
9MjZ5DlPuLzHLhHg8kH+kWlkSNZd3uLE+UboKOo4k1j5HNs4Ki3tKIW9UzNL+6+W
/z7VMI6RcGfmhnGetNPDB+rh3M1uq+CYQVZYfHY6YOmCRXP8H+cpAjx+F3rPDmi3
Xm7C+op+ENGXfsusDfIhFg30UK8faGuI3pJnZW5J+/nVz5mqp4Qb2Sv3GadidMkP
iVEHslhG04kVqkDzv31QZO/fDIy0ilMSa+eBR9v8XayPN7al0lMWFZ3PMfZTSorG
NEER51b//eCjWWriJ/Pljqn0XmrnWMaDzLLttdhn12lbYTddwPwZKg51FR1VtLW8
OguERHhEtiMMc+qQbhJo5opaF2qPFSvBZvDZDAlEQYqVzgWoiGsz8gvRk4y3F49v
CR3d/VLfiTD0Xx8dzIq+BK92azuZ+J6Jji9aFPetWpHchpdjXncSQ+r+SMhKKSuD
noJDimw1OQ802/nTn2i3lDikaaSTnK7l/FexNDoXK8RTpxPgp23tp8YdD3SoGSjr
4l2xAA+mWjbLt+8XaGNTVQbuzhEP3vEpLJqiyPqr2O717Bi9x5/Xb/J6cJCHz4Aq
UXEUTyCtIbiUQqZt9eBjxERJ7TBNeraufa8uswvMCS/ncU5Hr0Vh+jyhQznKu/SE
+e7nP4OF6RCHEG20dAJn/vQ1vL8FqinocQHYYiAjF+z8cH5SZ79DlpT8/CK8MJJr
wnO3uzczbKx/HvMsjVvQEY3+MhBmiHI6HSjtnG6RXcaYgIi7pmYSylNcNd4iqwAO
lFZxeWupwnTAtTfhtBpaEO2ydr21LFFLO7rR4BBcN75jN9BIbwaojg+OUhghY0AW
Ph3GFOzdd4B5v7hPQ/zU2vPfZAemVlrzlVSuSFy/GMxi3BuwoSnSmWEORod25s6B
PMlM16vkxKk98bcPBmL0anOVv4jWuoieUEDigYBRzGi7NZ3WJTx/zWrLYClOBuy4
Lp87yQfdBi5ut6gDijmdUgPlnhVQRwV9PhmIL/KvbVJ1gOGczOpL1cUWX7PoayM1
3pcHQ1He6xEU9J60g20XEQ9W+tM9/anavh5UxvSz8gUxsktdkLpyiAjni9/UkKUw
D+cWPYL4MMegk6SkxuvZBpJ4KWnPxHrr04U064ZJqhTU5xOBbgUD82Qf70VqnnQQ
Tb4/ivwHAHUDfcrXygXPZyzngnHVP63nlaeVLKh2OePHiQKZphO8C/j5rnUKww0z
VOZYH3kjWwTIN54qlneFhN9THWq1GP1ymdfy5a4T73rfDmlDUCGPNDryuFESv3dw
FV0ISKT8rtsWIiuX7itf58WbXHkdUtmuS40bZnV6fX14KDN3HBO2v6LnNwYSW6U4
mZDaJMNn+MmiRvFl3lutntOgJbOSJJew23gO5JhWyO7KgLwQ5RxblaO9FYr+B0sN
GBqvZPdOXIbIzeDovyiH079I4KWcS/xP2qm6BNzAsG/+DTEmlprJzYqkAk+n7NLZ
D2UZYYphXcTQL5m2EopJVKO0PTYgcmQoF2Qi9VYFHDeLPXPH3mfwsxk8oGVjxTS7
/yR41pNrm9dxkdvwzA6n2yXarcWwFwFog8yw0VB0oG9SepVOYlNET8MBCHSQXgzp
gqRUmA9Aw6x1NhzHCtLV1dgU1IE7TFMHQxHUD3G3ZUr1YLyBD/voVHqskUrRurZF
00Cf3M330cAsV+hzuiK8/zG/xCUr0tjojbgqLzkJZwbWmHOPjAqhkCr4o/2cVBIO
ZkwvoUC61TskuOEyZdjjwg/i52tAuNsR/2HHrDkJ/5eaH8ChnihOZ4mFD47VOVdf
+rsQozJEd0TOFh0zncePud46RF/Yuu0t/vOiQdZ2vJwMkvUkYZuVaY/Jo+RphTWu
Qa66WOIZOmYEmAfpUijJtsEfR3YZelzqtYU52AJUTB9KmuBs4x8BNPbAikZRXYRl
3nqtVwPm9TgunCrwNNLE+W75+10Afhy1mizwqLu8QPa37hF1sqfS+/6SF4F60ziJ
bH312x4ECO3I89p8xH74Hb9puMYjeiSNcX6Vt7NYYYrA2ymN9LtHS3BX5s+So9g3
FMvM+diwsldk3VMf669BGbFzmhlSpWgwIa9KFSmgc5BrIXaa+m7pM8soVlCeRHWl
nDW7tbphrXzxth8m1r7o1EndnJ9PbF+klcm0EnGMcFcjDRns+XJMF7Q2RcBkyTvO
T1qDweX4Yc8rqMuZRKclJchiMpjrL9kLQcGDXs0iy9fJer7GkSthHSJV12KDZyLO
fGFQw9Ym+1XNOBwcTgN5bnIxfcQoxQJUrVCky9XHXUG87Hc7vpetEire0JFrnsCh
ltrg9q7hzBaj7EsAhpYTpaD8kxSZf5rwHhycIUCcA1Q8kHBbal3WDqlZ3eNqeH1G
BQXzjOMrEnvrmwHjVXSSuMENkT2pbaEE7Cb+tVlKkAnwjdERxiLKw0z1FPVkYtyG
vRo9WFnvI7gqhF+fR01l5mt4ywfMmfaB6xcRPGsK+PG4FHc4kPQ9FSKwzLlyCGip
DPtPkspf9U0iqKjwCI06+VCn8YII7cAAQss/A1D35aSTACD+pEsCUN0wzT3R/5ou
WKowIhXkPR0EeMqIRoQKwWLGD6l3El8lsXw0EnU4na3ZBiuD6JYCF1rkqp9WPZxA
DKWNHpk86D48YJEtzXsNCNn6P61JDyQIo8nhchSFh6hX9vQY+UWXoKzHKGnsqQ4C
+4OUeXfOKowpzuyKDnpQVneVFC4Vp+QvE9dxXfqQCxU+slLBNnhIypF20vvL6B3v
53nQFh8ySvYyrTU5Kkai8nk6Ezy12Y4HW2xQn5WCy81s12jBvYE9IF+VsOBjoMys
iasSBUFd11P6gNmmXKCQZ2AQqQEH0XIMsKPYoG5CGbjFnwfX8RLXxaggPibLLRuD
GQgKI0072Cny764vVlbuQG9CRinIWowE+21C6puZTPiDWv6D820ryElURcrZ/TzA
1bGFcpQ43y1UpxKxINEV5ebHNPlHQN+u/xi/qQmt039Q7vGjX4vmdGnZ5suN+L8A
/eUOt8BPv/GxTh5qJoRVk5syz3tCyHqlnwCS1QMdytt5/tQCb2Rx8iqAM/HV81F0
uiHvQb4erhPO6PD08gMmSOnS310/wpbPpESpR/3XfcrODBI88dpTILo6yIne/L8N
UnedWbYls6IKjDk93ccL2wxa4GWrJtfiMwPTXe6He/wj/DVooXNKEvs5M6U6ngOi
+/gQyEFx2liQBZakPu82UAU0z5rCzH4bCDbsiVLd4/gBjpO/PCNV09UaabL2bAiZ
R6Tf5kPLrZVRDgSgLuKf9Tgk1rkwi9vm55/OYuIohfIxJvkZybxqgZ3FJlDBXoXc
MEhnnhqhT54De6qL2Ekbqeimu+jTUF+odI2WJRo2hR5i+x0d0iR4d8Jryya/kRV6
77+lQncrm6WIWPYT1u/7y+FJ8XdwSOpuKV21jgaCJYFrit19vFTpGcwoubH4eO63
8czufCQw0ABShR60xEdf5xvlkQ/N/SMI2hZpKT5aEhaKnbc5QHECR7toaeb6LFFE
z/vdltVXh+d/zWuK3UGrXnCqo6oBke6RfdZ/SjMwVpxAcwVhvXDW/PAbAIgLfb9P
4tFOdohG6xCoCtAg97GPEhkOeBPc5Qshdm1ecYGQtqgo5V08fwYQTJuFA6Mzt4As
D9VbpGHI7jjSMHMrTZ8UELUYgPvlT2MrdJAEh/NIzzhN9PuJ/DwK52j8OjZc19NX
zgguqHmGmCSfxlZJ1/zcGsN7sa/TWNUeuw70mnf2KKzAcArdOFdRrYaGVLO9mRoG
xBmbuVqDoGWKDEh6K5NZYJhh4ajofbggtqIHzZFbP+4sbSEZENxkVpZBmeGiR/H1
4DRklaq54Hv/P0L3WPfW4Q1dAljdlX3oAuPk21u+Fca/rc7DpiMVAQMR8agQ9mub
cM/XppsabsxYrerv6FoBTn7e4jbzl71nzO0ebDttHpVUtzDr2kmnrOuWwQwoiq3j
LeWnK47MwJ5qFbUgrfwVIPqHvqD7UdRtoatpVmHOeuVHviDFD10lx+xaVhThQusz
ZkeDJc/yMNGa0ORPuUSa2CmT3wGAOJwNxGDKWNkE/wb3Xl6LAWFW1ybrvogrNJRe
hLFr/QKwfou0Rfu83OdG7INmYSU6l2ar7ZoYarlDANggPPhDkTGlMF31SislAfBB
HheAKlOce3U15MaktyQHW4zaFovRPpSs0rvKxqAkBNOlgVzshv+juTVN499OIafo
jDXtj525RBQERRRm6mOh6TGN64Cr6DPfL0LGTVKbpKutXzisK4gR5gTDbJMjxLBU
w0RaL0mGOsD/uJdnwRzLy6UmW9Wtk9yxkgItNzHLj9Z8aOwBu7lynY8AfiiNv1N9
4Yx+XSMZPp/1x4uJUGVwyOzH/KKbs0OvpXFPsLy2OUApTLLeZ1DEMQyTt3zju9hk
0fBNAZ9f8J/zkSoFV5v+3IgUCPzKrM6X17rvm9A0VsshruTsGldCD0FYRioR8NYX
GbkMElWEpwIhHjjrMEnpMUCBxNx2GAWfDb+jc16u1Xc+U36xeS4ncsASyjSEh++b
RMFXbOiOBfayXIA/xYM2oWOHIpRIy0wngP3QYKszJpCqQOF4zjjNCz/AGB4rivgX
oAiRLcm/sPU54wUfgK9Dq+8x69sImyFzKTxQwlBTk8OX8aADTXuBnq6PlPQ+th/j
WMvKTBPMjHomhmbpREo6H+8GfrVuSdj6tohj8r7wDcJ2hCpRcMlf9KP002xPuLQS
F4r6hX1lEMmjLsZzePqLKyx4S+AgUXYb02CRn97kRLtuwnuDI4wWNZWAFEUbJtQU
9vWPBK4QVYr58vwuh6/qchfZ/5/x14XzmZ5bwxv2HYoBHChPUWIuX3IKOaxgWxZk
Tdc04nzWZX6SbTHUc0stowKkd9TVVeFVOtVdJ3G/HU2ssJejvt8fXKGiT3Umq9wC
0tf8J2+eGlHj7md+f7LnLVeFZCFMkBWvONz8F5WQ3iR63ZYtM8UJYY8d0Ms1gYMj
B8ccJHYD7Pa4xvAtY79BWcigdWLJGdSJCrWrc4LORXp+30fSE1ScjjYdBwu5BBnf
IaOfN/S59SY5SJd1cjfsNqCSGAyJEG8k3RgGSKQrVid9yFUewPruYUuFDMqgXsb2
gsfTDYrrg20atG8+ZtbRYw20CsiDenm8mYbRNO+6f9ZTOjc5hsWt/pvnwROz13aW
bvIx2V+dYtbe/Nu9BXhug0ZnEt1ai/gWxr1V0Z6ap9V44Q+hfY+n9R1NBdoRCkFw
8hHvZ0biiQ2K9d+M/32LujsDbHmrQy5JOOcH31Q4eByUZFxF9m7I0LAcDvAzUyzw
J6N1D9ugsCVeoN83XhkfkAILw2bUEUKseL4NvjTNQdh5NqPVpplwZSuediEqcr/7
UyHZEeZRB6vDPK1lffZT3OSLmMg5ovEE4miEbYGkbdQg6okzoXp6XYlq2Gk3LJoU
PNXhI7muhT0dEcmYikA2l9lW+AqhbXZJoJw9ncjuRSVyntACUnM46usCypGLsbQf
rtThhVribp4uBrA0Ye84O+g/WT6U4eSRrXnuZc6jepbDH6syZQP0ThiURWICF/UT
M5TaYnNN+bInIyOBeNJ2P1lAP7uXzcU6zW/edpXwA4fm4XUAXZ08qKXD+X8ZXHeF
EWKxL7qRiXG2kPs/36OHLL4nUEsyV78sPUhxL5KtNMSidqUosb/M2RYZOMQC7T4Z
8VQugK+BeaO2Gi03u8xlW4cV6xmYvMp1rC2dI/Oo1Xppr4KmJYmJ2+4LolpjOCI/
C8V3Yb1CjHwoED+w2eAWzlM9MZPbccKabwfS/Zj8QXYFCQf2hX1u93ImJp1mq7Yr
UDuCW1NwcPKzn9O92EXolgDOdeIq0aD4zBQBnQpSoCx+Qv0bQMNsaQREoC1ROG/m
HasjsvzFpoSlXgSv1cENdohPnC3e055cQhLQodyD22GufbCbdOesEU4eIkcGCj0v
sCEWLeKWOfByw9IRsQUgrZ9InvtUbFJNTnDqcAEFOpHfvFlvfmHlOcpqEHsuvNPv
hQ964L06l+XO48AZ0/o72Xy8nl92wLHhLEXZa/b2wyTOOofAeY+mYMxun1+jnGPL
Tu/YKVkckqDLBtMoPGdp7ZB5JUxLcvGEwDOro+goevOmYyR1uBgfZ6yFfJa7ROyj
uny4s67rpQiL3KWVhspAMA6gmq90/d6+f2eAJFJudI/kYXSpK8jqVoww0srXsfgp
cKzbCIcVNXKj46Zvlne5FbxD7qfakCCd3+6at6AV8Zc93rFd6LlfvNHpFqgZv/56
XQAIGRh6UOKqGSFItN/JKXYVZl+vakJWVzKxdflwt01JNEv5vNwHsfAX6ndfZbrV
uOXYBKv7xn9JaD7m09e40JDzB35XcpSr3cRcmj0QID+GUem02URp5agMidRsyWki
ju/59OjPqPjxj/pnfKA4GqJrhIe57R1pMM9tLCakxxpZ5SIdW+Cccj6fQCdeIyEA
+DD2JsmF5BwsZeFAfaQ5YMe7r/88MjNIpM8RtzPmoaq+KnPSrc6leBRYusejYNpe
9jGnY2qalvavVrHoeCMAuINtRjGrCzLZEQyNrkW0Obo43n+e+y/EOw/IUpkgp/7X
KK290QOL/C9J+zhJbWSY8CdYSGZ7VYYfuwXJO/12FZPu1UR4B/S5UNK15LX3AJlI
JaZnUxNGvMC/e9kXnawqeOhKQmvnW4hTkZQAK7S+c37Om2ASojd/a2nPGF5Clvf3
SeTV07XHt0fBUzn5bhbDg5S5qfGr0ts+GxU4TVYweR8arITe4sQCGjYQObfUOGyy
ji2WRj3As2OfKGZmCURgDT+U8NHr1GiZQE76uTmKqyZyf5197yWp7UQubUU81KFY
+TAwI/HbpaUAfOgOqYL5Ce8dC4sczmg83NPFkYHjy6ljCUeE47KM+RObhPNExP/w
idIzYpKuQwf2AFfb0Vh7nIByyPIBqiZLLbv2XBzzZbTNtkTo7fRU3+K040GF2tnl
E/N6miq88ayfOsvNcINMi5piLbWIHAV+MuFK/O/cT7S8zmXqG6IVFQDsmJYDCQvb
k28a4Tg+uD6YOVHmqwd1KyR0PNecqdLAlMl5vvLB43nHRQzdQKRLN8aQF1hvj3Nf
ExBI/aW7wJeWm8/grwYDX9uYgDkWXPtgSXXSyicckGFqmCUxD+IwMoxsEvbgMmIH
tXTx4kxf7M1DduoEkpzvYQyyf0xR605GzsSEzkibyLDV4TW0jQ8fzppF8fHlI9Yz
iOfxgAtO1z/WOm3DDDuQswLoG3hal8zbuFgjkyjtbKlTm7ULur9mcW/6Ki8cgMAx
FgRwnSorKXLvjsTZxOKXQO1sBtC4Tcr+yA8Nvcnr3N4MdhXcYacuoCR1RQVCE5ik
BHRj9ZjtNaWtp7w1XFoleZbeqSViin9ilWD0+pDVD81OLQrIARB99ZdoSrIZWxwy
0sqUVZThIajAFAeTIPR2MjQ+fUOzVWtKFKL51JDDWLdQ14pG6QW2hKl4aUKb13Jb
zeHFLpJPeqsAN68gfVBazdEY9RDt1b9IRmZN/ttrNFsJY0Iqacffu3LkXG7eBJEG
foitxpLwNTuJ/IX+GwKfYWmvZL/ktXldYmSnZc2RH+eqP76e8+mkWdmA1meXNEh5
5UrZZL+aiePan0q/GG4jgBqmdGg477FEac9FjCa3+ssZI7e9lUOb4IiyZYltVdjB
i4BX4wq703eB+Ejj9nWkobQQVLWCLRGwWU8FzX5DSmhLNK7jqXWOcUJjQ0XRi5oe
OypbK9jiAhwjQvymD30Zwm0DIoFaau/PdQdjQ4GsRHuHXAuA1qSQN3IRzQdq4FPc
7HDENog+b1Y8cGfe3MezgmEhjZIFJ6J7LGGBXv8IjAYGrEuvrvou7v15HUfeKCoA
Vizx+fwlFzGClBK4Y40IjpP7EZ512J0LXaNRtPCymS+SEqyv/0fQ0ouPTGdnLwPb
URyDH3kftjcGoQUKbsGz/mlHRg9voStKS5ALQQLYsRzAMeUc1+M2blyCnBy0z+DH
dNjUnUjc81GlaiTVaUntZJ/3h6YIyXnuL9oks6f01mLGNPhBwQJjmIWCMjaFff/y
HoK7Lzj5FEq9kYacDtsRPdYowiKM50wkitC591h349qHGTywducFsIRRjb7HM7jx
M+OPXDMgI9V+PJfrzMeoAWOp9PzOPYWvDFQT9yLbzlY+jKXxVwKaMztzrgORR1qr
gZg+lUqxUjkMwhM3BCEhvOIs7aMQZydhpepb6FuNWnSMNL2LmzUsZTDLAQFVSAk5
WeSog+8WZQqTVmmnusjticEs/yRgTHNxK/HUDeM+d+M7/d5EAPcRevzG1O4PhBRS
E4Shjp0mKzYjuDK4sKGbBr3/1GYBWJbA+e6B2rqAbV+uNZ4JEYT6OaLxbjj0FWGO
ubihxnzojXUitJiVMYUOohomkHWc/PSyRwsSMk4ohRFbAefgUqkWBpbvI8fSh4wv
Gjbkk3V54ce45q85wRHTPJu3wSIBtM7pcsBk1RswzN7Yv9Tga4eRvJglt/47UVel
jctWw5YnEnlHOds4pvl0lBApgSxHENrxWq/cQ6Bfz7Mmtnh9+cG+giXsz2F0ozAu
I35VejJFJUMrOGV0AMGTZDwABnoqU84rUhJGF86TNfnJZxTiXuP8keytE80kotF7
cvQiorOispBn9ii3XXBJzEy5ScknKdwPyTVs2vbM97GBgHVInk08wqRMzX/SSLpJ
YHlKGdiO8JCRZ9faHZniXrGS4BxKd0iPGeNKs330P0nIG+5Z8NoYOo31yY/m+O1V
pCATa6pZTNYlNRQT7qqTRrcyzFh8Dgw1QbXYYbOjZX/gJU7hGtRFbYB4Z8suhBZ1
Qq3l8xoudc9MymosLYa+klWlld3or49YH8UdbagB4catJHXFxEzHitj8Wmxg3ufe
deocyzG7sb/YyOpnktwWoAKY9tcBDMdpm4ZNIUc1PhEMuUWQEFQu79D2TiC8hrTx
zkYf4v45bwrQl80WSgHlmUJiBdHkC46znhId4h5uE2ftGz/DTFQOFk0LMi0nMH9u
a4BCPimrD4DeykBrS2j+VObSLA3BtpTxBHOHejO0vb66XuL7XvQJCzkacNWrh/83
bxTMJgT+5VeZF3fY9zZrLGG3sCEi2vLcs08uOS2tm40HqIYOXKsLv6pRImIdcbdf
40E0+/k/bKd+0WIeMibinhY7o2pvDQ9gxq8FfnuYo2uS8C9Q6HfZHD6MN+3cJOv4
lgncuk2VtlUFC1Fiy+sYfhn3Y0K9zrtpRqyAyer5CQwNoegR0rrwjz342//eqYP+
plNKQd1tb0V4XXY3Y+/R/11kYNAq3PrEY9iQrBtL67uM7hrMdfnk6Nl+I6HCRgmw
pvTJm08n/9Odii9Rtkh1Bxq6S7JAbAikYF3SVzF1BqFZ56492J6KaSuC6+/i3USW
wCywzaDpviP8PiVLcYhiSqJxOCO9K9ULbHmUQAmEq9RkrxUefF9fPESaNiE07AFw
OZw2DSAq4NahcE/JmbYZGyae5X/vBtWexWA0oU0ChURSFszIDH3Ij890+PrakUH1
utYmAmMTyiZiq+rlUjeRKUbslE+JthMMbui1zEU+EsByNhwQ8wTTHi+LefUjIyS8
3xUdmypfbCxjEcxxVMPB6OndOaoPnM+Nl+C2cExVLiLv17PT9MRImxRW7BaEyVnr
bZ/CVnmrnFPMOYlAwd0u9Od/qv1Wu1nQnZBb57ewdSfXyAOeziMKrw6DhBKgGdAc
RMtJMT/cBUt/jDYx3JIZ7/NLKJqpL5YwJ8btDq9zUq/L5BtlOJszdXE2Vlxz1HRP
1DmoE7emC2wANm/L1gVt6r+ISifF+cgOIJkGNxA8msNZKanNwa9opubVh76YdQcu
OwLFPRGp3uznY79iZ8jJHJVXHm1d15OB8wVnmFHiNEP/ZL0ZXsiLmCuHeebz34lZ
ujJTszvmi8DCagm69r/Wr7UcHoO3urk4H1qrLx8AQBZnjUUZag4vziX1WfqfL8OH
NWu9D9nxjsuci+gt/ySy069DbOVVSX/c5CXkazHsp2WinH1TvvAjXuykLyvvIvuG
5GkjOWtMZTNxG/DSCgTLnEGN1RHQ+5pAZOJFTqRJNx3/L6XXvGulqmzReUrcZ33S
uw5DURXJkJ1D2QV/wThaWG9lHJ0DswXsJrZvKucKZXih88Ok4E89vn1nyRSf49oP
ZUuSIEJfXq+NteoFArrCYfNYlwPaC6E2m6ZL90sqWuAEBni4Sw3FLHFdI5IevHjn
LrII7SZuvMomGr1mRJ3fQ3PjbrT8mK8DGOTk01ly/Ab0fdYaLpH6bYcoARcUgdzP
vIkEofrWjFPGEfr/wkb6zI1u1ZjJzPAgAgoGSYXaSBgT3scUkwAfN7+4A4i2tcVl
n6Cx4/7Q4AZ6pS/MaILi6DHbyLSmkiE76PP5ndJx2zlOT3JRtGZj4pLnyeCB31lo
fqhOF9JpVNnHKX4s8hnk12HoZgJp2Moc1xvrJq8j7e+dJ5Fmx5U7UnIQSo1uF5mi
XQ3xMHou6G2ntBy3tp1vsRzI83RWfHWVKKVPaClC/HIT3oAoRE84+CvD508acHyj
vFKuFvADs6ypKi1yQLHTPXD2mswMzquKwqLYCCOAShXV1blxUMSFE5DyZ2XqIu+h
jyr3YpmLJ+nTffHtHNovw3vxleMna01Fr2XHSvwBxyDN6WV2UFvr3/HoFG3/hqQm
CytBUGvCGQy0MQc/9gCYr/8mK43V8oxZCBRfe4r/jv7faQtqWZCN2hQ7NnzwgEsP
Ib5cMIX4hMOkBDRsG6s2iKqxbPLhRTgwC4GobgGLDu51i24aGlSitwcrHGsKZ+O9
uIHed3WDYxpGt6V72cbrB1N6PibIorFP300C5ulTOe/a93+9bi/HAt+Ty19RbwsT
SYPMY9WH/3YjiIhQyl8mjrING0q7D/8tzOHxggSyEKUyjx3y0Mq2DifN0XJ2t7VU
aJDDgr9WSuITAjH/HTSMXcZ/jviSHUAnppsUpfF6UWVwXxMGEup/yz4c3hHb6tGB
trdZrm3IPCVoHUkNxe6rJGAHrQRxXpXJSeW1OKfzJf5WDmRvgxNW9EBjUYulf7kG
7V4jA98YWqt8L56GJc5hpxjrm5CkIe3IvZpGGWu8HYGiRADlkiiUpCHYU+JdpF2Y
PHjN+v7VghZpAxa5rrMAurVJ64lWLolZigoKXVCSpNHGo/kWstQtuTleiW3Vqn3B
6+p23/NN3kzVw4GVuS1nsGNXqOsUuGH2OpbsxykjVgkJnj0ciJoetGy9wjNp02Bd
I9CK5LBfrYCTFCl+gezbx6eexs3+UVNItdeM/iLPSbtj0bUGCXiXCQm1FUUnISqY
dMYVgt5J4F68EoL9bJnT/EJ7+feBZI910qLw6ETp8T0wZhfxVsi3o2cr3D8pzGCE
+ron5B16PTQUnacFmdNwhWt8n+PGWSADbZ25TiWP6b6yGA/CuvluTNpBc27Jdpf3
v00E+jzrH6mQmsYoax3W+bdpT7Rli8x2AtPiEYrk3qm3MigNX0sbv+a1GwnpAo8u
UMYvXHxqwPXHhowPZwWrDlFAJnfo+qkSnrlC+O6tpkYURpFSw9TL1k+CJLnwQMw7
bfYKrLzkRjoh/WIeRdsfJBvNur3KAkupXnoHM5iuffmufw8JW3e1mBKraRf+Ukxd
YsnIR/6D6msv0sLxiAKeK33VTgNYhmNO1vfkAa7oiAK3aJGlWp5C/ZbZbG3gXLdn
qe0MtfNJ60txUN0NabDG630rG1zIbj2rgEYvbyCWmbJRxtwQVpLQ142Impbj+26D
c5OxxGSKpN0c1q1yN7tvFgZYBcZ+UKiAECR6z4sVGEZAIMnAiNtGX/aN8oBpFK4r
ZnIHkfSPaI/6zKZDTRCYBPRKPZ2EmR1STVao/C+vP3ps0QnR1HAz8B4/iKNegG9P
KBDsHuj0BOiMksipdQz/DyM4LDZayFSLdNk4w5VT28rcrMB0HFXju12vcadimVJ4
imRbcoNBbJV0ZCoVGTF2sv60rlZNQ3ni1/VGNJ55DuNBt+B37HzQlVbV/KL+3Sjv
VUqrG1OBTOO8urPfTFsNs8QMv4VblNf/Os7mVdjZfimqYxblNScSgxqpJN9dzyRI
N8Ej4VCWXpz//wUdGl7LQ/ZUdn9TqQtDjXhPhUTgxxJfbRBfMAzbb0LTEeBzjhqA
gV9UbqNVDoDn9vCxvHnQvz/Zv8NiuNcukA2s+NPl6O3aSYW+89+ptaXu1FKoplQn
2jBNfGAmdBilmD5Di5xCqRYheWrwCVSydaEIM1cyQomWhXOW1sZ9zlFzYtp5c1Ui
UZ9vpcGLarvEhegnmBFrKIW/Dsy5frYaFpJBnGbTkENfSi7FnrTv8yENXG4Hr6oU
6IWiPEKhrfpkiEe4IR0l8Aqvd8Li3AxMVBbn3Pm6+n117JAk7wI8wb9vPcF6VrnG
YxhwRsQ1FaqvXvcuIYHbxrQ6QVOhOZX0Q+/OBDKayD+Xd7GehZWzqoCe37o+XECQ
7QRTJ/RISRP/OaFd7LNruaNhC25i9tdZh2/o+nKNwymln7eevKk/cpCMv0U+r7NP
eIQUKT0YLyPT+5D766AWizm/BQ5xChBRcvfgN1dtKGiafHba36uQNWyxM3wfGMeS
dyNIdTTs1MyuV3t5JH7X5Ixzpr/UU/Zw4ANOXpwW5TwdDUlmDh7+d+vAPyf9kOG9
qXOaWI9cQhdXFeSIUBqPAgqtTryQytLADIaHY81ixOK0CbckR5njmLi7WgvNA7Ov
6yQMG4wq1QS5u6VUzH8Wemi2hei5xaLjls7NAQ2O1VIdrhdxFMuBZwSAOc5M72VQ
1iVkzCJxferByvfmtvU6WIX+WtqbyRJ0d/olv8W+QHwz4c+uHvRmVnKsSXiyxnFB
j+kNZ9GQIRJIk6WYryd1ziQDupAZl1fTvCWC0l0gV0k6uTYl1dJmi32CwMyztDZd
pcc60uO26MR0oeZ6em5sRxn2vurA3H/Sj9QhIKiR64Dh15wW7Cv58TVW2Cf4Ri34
aC3O+K14sskOv2N4HestQFLH6ue4D4YT1ltLYhrvOTeZn0E6g4GXwjVio4/cuIOe
EwGQ6bmX9NUjAr9e+NFoXTlmwevlmKJJnaIlTpaTTbek/Nl27HhUzlm8V6IZOe75
be8UJb9geimEsfV5gR2YaxNT/BfmRxJkU9tLk5AeGj3hhm469zr9/QkxsZMjYKYx
YKYbr7+gJ7I73nNkE27Tukjm8nDfg6ncsF35UzwodCucxsMRmr5hee+j8BPXc1Ze
TObOK3AQFqGhNgSXOI1bwc3dt+ccvuJA7us6y2QReMwvAOgclp25AdXCYZK2Qpvo
3/PaE8gwBgYmNxliCNQ7UCixT27qxM0QxLNGs7OCXJk92QL+HgFivJFkcK1R0kS2
WnJSdUKSBRStV6CoeFRp3x72+rShiTFkE/P3L8osBcXxUik7UrAvbswowPfL+O7u
KkNbmtWzyusZVsCSxmLFlhDvXYJsXkM9SPhj4lDdYWT5WAgfI3iJLfNtjM0J4IYG
SdeLTbl7MEIUX/J+WTqYfxjFmIJ4sfLAwUXkYByHXkbbnzMOI1YbyGFxwQJmotm2
bzcUTku5Yd7CBEPcEbgluS3hs1RAtgwg+XPgiTv5hl8k4R4T85/TcCLjFktcNlZk
kF8cvEjL3r5u7Jkyce6lvLix++7+yauZJp1xdl3zukYvBKH5UPtlAPI9W6wd9caI
ytBm7Ykaa8yt+hPq6Ww3g67PD6R1HsRqSpD+ZgmCp4DV3NN0HyNxs3kk1BLJyIV5
rieqejPVd1bUAMgX+sDmk+b4SNZtuZ2B/5gBjN97Tw7+RjkHsgBWrIUDEF6Wc3Ir
Jme4zc7/iwx14fgK9z7GgOW0BRp12LN3gsKXqxCaApJKeKPnN2LzkyL9Hhbj2Q/Q
kzm9tnvNvjZShvu9SxVboFLnwsyh+WGGX9zOHbK6ITzDCr5XQeNNlta1rFa4VMmN
Nl6jUk1fcv10i+Mbjyhrb1PPW40fm3qXv6/B9AsoPzg0CJZPscpAIBzz8V62CJTr
CczAQCUI/DEKC3H8fqe7uaVh1BDhEujOXW1yRQTtth+rg1AFiAnLm/JsFxUkK2xE
RiZL/jdCl+vCkhcUVACWHJgCr+MeKXzSgdNjuYclpHXlqY/OecSCHsWE7EiyDvWz
Ms2meOrR1f8cH9kjuUfygQKvAK1fQ9Ss70C4lt+fAERoQPyE1Q7A+G/iHo/V3Dr2
+9l4Sd6DJgw3vNlgYP/vRnASH1DSA48aUBB51NnoA/Ol89aJtigDJ7rx/Xo1sJhy
6gg7FwQhEkS+c0yXwn9iGU18IoU1SWZbq7z/OHgRK0x1AM0cqriakvyiI1/yppKx
9v5nsdx4ocq8qojjrDAK0fUDChGBzw2pfbcQVTYRKERs3ryg2vlJpee/sq3yoFiH
+wSoFHHscau3SwyhtHH5sC+3ik0jVLmL88ZYoWUBFku2MaWbvRfIqnDUiNUqtQDo
PS+uk34MojOM9YBTBEZdrVcs6wqEFRWP0POpGOQ0c9an2GoISx0I9fkfK/3Z7Eys
t9KGKjcO1t75lFR4FSTbp4/b7WxcsjH7M1rmtNYIrkY1+YrY4F1v360irc9ZME4L
QU1WJ8Clk7vaS1FvMdzC58v4iJguMEeHI7A4Op55CCCg50uuDjrybU0tJ9c6WGCs
ReKT8CnkHPM8tEzVmWQa5BVY7CIU6lFe62OUFZ4Ds7zlAPF7Mg1jUjZtvk1g5X/U
PcnjndOY6nEN/ZGwV03DY+8Fm4eCUPKxV0pXvPkxV8Np//zzzLorkuNn7rf23/zM
zfic+XCjOgJAhSP9FtiX/64byo4uyaTk1WTsaAfTSZWFNjZi3EJbsh9s6ItXx3ic
buinpkrhKi4piH0h7XbpQZv1OJugR/n1yZVdcEypE3A/03jIYv6gM3jgJQ92g4ku
uSJhDFwwqTROT70yJvXxoDMpIdToOIdQJy28tQ0N/XPnxJ2XfcGP2nWIkTerb3Sd
RjZpLd0tuDH2ZMQBBsOtj7lYFTKOcVgzF1YB2RdVSuUEnjO+BBf13/vquVi1GEmi
PalbRiA+Mf3Madn/K50wMAirlu/EK1KNoODLjZYYp0ZF63GBajMy75t55Lny6QQ4
OBGWD1uT7NbL5EWLVIqxXdMo3/gCSCL8Fyz5rNeWis9Oo1OgldZ5jT/QqRPX+Tvm
sDSYWstbWoza3F27DOwpdKuPr+3mAZFIyPVdZqTwQjfiMvn+r9FVuqn6PfkPjFk3
lRZn9UJKCKSyINE2OtkBQfw/3+omhv2DfOFaclfwsUlzBVmX91qQKfjTUDsHwn8l
FD4791z5+q1zx4btyTtDrsfrrZqMv62Ke+fTFbaqqIv9Q5INyzYydZgOoef/60OY
73fAu7H6NnR49VphhrROlQxcO93R1LNyU1uvGgUs130w8V9m1I7ALZix2rMlF5X5
+6QcHm/CkUJHS92R0FQargTuPnirDnRmaHhAKulA4YvK5hDKKvmsY11+01GOvi8c
LrLDc4sDI5moYkcrnb0YQUTGCEk/C4PcuIOpWsx/xUidEWhcxR+uz3TSlw/yYx7r
w3T1toPrb+X0EARol5Uzjno3OA5g4JYJdiitY75n3iQcLNdnkVNyWkV2w3RGEnRn
LVvzKOcGS5EB/As2g9G6XAnLC7OGf+SVpp/jkm4MOaNDY3RdSbam8wy5hi6OK+Rl
OTNr/NmUuZocEvQUzaPSWmfhwGx0nTEBdfp6Zrhts9FrwfhqRqcMHJpXt2HZdy2q
pst0cysBfk86SbwchsVWSAwLZKEzRLEvRbVHWVOW2J0l43MceFinGO/3NBCxfIuU
zuIs1g5HaDYnq7iLWmtiWaa9RHPyI3K3cCfZ0o630MJy0B0hVDEbGQEw5rZLsW6I
zplQHs0U4I8A13UUVYb6x8FN+oNQKFtP/Su9NNe5SeJ3giM+E8lyAdgYYs1FMDFV
iCjlmCs7Vyw8sF3wZ6wXaAAI2soaBkHix+WiyN39pFRI3TuF87EUoua92jQN1/LO
n085vbsiBYbLDzZqGcizGj0w63qMcsijmTZUErssefgoytzZSUme8FwIdDJQAygi
hIzj4KTV4TULj1T0TQ9ocVR0bXQYWHg5gGAk9emEvKUVuDNAI14uDO6aPme5mpXf
XKris8HecHN3S5GzDUUjTfOTweNmEtTOF5CBK1k9ZF5cdnJNfjkhMd3JhkOD9P1H
Tqn8egGLGFIxBIdT6aA9Tuc0DFWSmjZRUmwE83G17pDzXi/5LKPDYUsPGyE1eL8x
epywlYDC7KRrX+hiaBtjUzRpxaoXES5QHjoIjhxyLRnWvMW7+UY1umfX7EAnQvxO
VGcEwWGokJ3LOPljJoUqZM4fxCJNrw7s7TnAtE+wDWWqD9l54iTWydoEZ2AFBtiV
PsrAaZ+ObrbYKrD5/RK19QJixUhLLIDdzZYgADuxEnjGQdae3o+eJaoPKKSu6V0Y
1ZjSSBrlr5BGILxndr0RIz/RbCPUzZwBC06PiJldCDQXrU9sj3apXJfNzzuxdjpM
QVL9RLhlhJI8cJiwezRufCjsVyOQVI1iK7wtYIEnExGsqqgHeK3ulbjJhL/+eXua
da4hTu/PeltEnW3l3XFp7lmzm0sD0W3Gq4coNZ3NdKLiM0wAp32IfES3OQu4f+FS
RwHe/aP9v8omH2GRiXm6M41sAt4bWLvFI0TV+6CvonnqAy/wzQpoo/31scClLnX9
qRiUFN4va0I0vVIeCe5xIvmJ/cq8gXAUDo4zQ56J8iHA+/PNBtwyuKUu7eAn18bD
O3jNVdcVPnszX/3xDZSX+le6DcpnHacWShjFiKLLrpX2Zm7t3V8Y1qQVq3ciB/W4
YPU6tnsiRPT/Ve0ES4TRAtSy1CpD3E9bj9t6dLbzkYjcTSCm088vdlmn/USEsK1E
/ynRm2VvWs0B0W5ZxtWT5u2MoHQPhDZrGP87ak5snaO+vwWeYzahu+PIvyfPMNGO
qqnaS1AQzliuoRk0t59KV09uHMUgMVi/Rg7Gqc+hMw24og4aES1uIK9QAax67jUm
2bNdvaS2eEofidwO9tmpH1H4jYg0PauoPdR8iVWaqsxmykIP1cN78T35nol7NMl2
gFvlrA6KMbn6Ep58YOyr2gYBhxwHdaoHjH2kqSGBSHQcHki4nq1Ez5W2ZKm5/G/d
mHLCwpbPnMsT8fbrqQfJkzFnzvyJdRGvzS0sSVHWShuhQ4IpVNxzRI7Hxd1rbmyq
86UH1p/ilGzWr+yoEvM1KJb5XfF0PC+7A9akz5e+fla+jfz4eXLP/NVHriMC48Al
fJnz15Ti93IPOjxVdT2DMmlYCyDgPv7iO+i1JtnSj4BMnakNPZweDc2OBzsgHfVN
sXkKWivbNHJYb36XSEh5nL3cBhFKVx64tOBJUJx+ZVwmbK0A6lfzD0z8SC36SbYA
xFYRidaTRD4pRP28iT0w3dyR+nhp4b6LSQ6avIRSuqdNI1t3iR+Kde6CXzXq4TiS
v1EG/StdNhrhq0/41wdOCmN6zvrJMcC0Z9CkBwsWcj40rKJcZRDteiEr0/A5NT1Z
5AqNZhrC4l9vwda6ODxM/IB1D/53+x0xcsK7KRXzvkE7MgsmruWvRK8JMvuqZydW
lVhOnvEjBgu/7cKNSR41A/IL/dlywl3bbtxus0sJefa3jFPCuN4szL9qohYznFR6
kNDZXlIf0IQTsoDhdjvb0F4jLc4Nvi/bF6Vloo5q63M5F/R/fBAnx/M7EKnzJQzi
j8m/Xu4NvtNi52DIvrUotbBDkBdGjT84jb5QTI0JYZLz8jzlfeMNqEVtEfX8vBPF
JS9uG1ZKn5wcvhRhHFdmGeSO/0pGTGX2Ol6rB82oEbfOWzldwI7uxzXBTkGfVHLH
w/v5ubEThrRsCR8jpoQqdQ+ZzDxsRKgxjYvxjk8GRRuSc7FbkaJIzc4HbuZSnTDu
r/XHqivEvWjuwd51mvCC+QZwxUjKAQfZ50AJ0neG8NNmpHz76W4aoBgj4r58eXRB
1gCmxtyIEVqX9oxFxjzUI+Qqexrrn0zwUkefEufvOyyDSDTsCNpHB6HiGS9EQHid
H/XBxNiaqb42AfDUgC1VpIp4aHk4rOT6Zvh9xPj/t6TRf+L5GiU32OwdppcsVnkK
BIkUmagcAMvwi0CrUlV/qP3QFidW1S3gZGYjp0IHmjhFk0lWbeqc1468igZIbv3a
BCujYHqW6YQRu4J+1ZzFB1DpWlw9uEt7/ZJNHndRwn2PmKF6pMZUYp0Y7wzOgALW
8mkmqS/kv3bytZQ6T/yr47SYyTsL+NDb4mxWIVAUz2cyUymWoKTA7EAeIg5iC4ie
eXp4WKHY2KDE5kWbr1oWZc2mBqr7h1M7zJVDtA3YVyRxXo93W0il4HpCMlf6PfB/
JnYdVd936kXUlWkehZvR4pgYMBmNLJSKr6Bq78Ex12gnkGZiUE5O0OYWRJbEfp9r
LSMY4fixX9urUDmTwiuVJMkkOwtsZqshwAQZahE3cM7IdMMSYJCauIKvDUmBQqPw
EYOg09DjP5RZaej3D46cJni4WEpzOso4hZ48O8PAD0op+1Y//JfjFXr7gwoJ7/UV
eq+yx8zIz+q3c5JVF+YCLLnj+9cHB0AX+zIKskRp/LACqfuBj4ZUXUT+XXBXZRr+
SPF0XItFf46DfOXdxh9agzaA2kMK6oP0EzDnCy+VFNuKNncRvzgWEeJg3rgUgBwZ
Iw+PfU2TFSjU4c3LKSRI4K8TAf8NC/kZybC3PWtRRUpcRvYHcSIIl0GvVf7vc1LL
WnKD1D1E4pF4JgHvhKRDnEuzL6bQrgD3CvqI2TTeuxRDV2A36sqtpPhVXsUFIXEu
lNIVI8LfafS1sERwJUEh4HsRWeMkH1ErZkHgcJdL5yQwCaWcfxCubUc//JvUb/Kb
IxADwd3I1CeFhZ8AXwj73qPyWG4O+SxVPeXYhlT1EJoRjwHdiGwrB2h5FXDFOQ5W
HFCBGImSgs8u0sjEhnQymTE+KHgSfK60F4SbSYCYIqaJB14QLUG3TuCyDjsiMvUZ
jSfH2kXxXbnhGlIKGHFjA1MLNqmrhtq21W7VLSdHpq+J963PVbz/bSR+OeJx8JVi
+hBlJSj0GVXdOUT2XQFF93llWB8EuKWSCRJ1eTTJam165MPXXg/s9DR+q1TLgYi1
W6O9F0BMepI679nch5J9QXQ+7W9DpYdjgD4AE9iaWANml0AlZha3Nazv2VKFxQSa
xampWyN70T4YA+9fnzsz+Txvesq1RW4m3zgkHlVIRCzJd70Q7KUvKTr5hzm+jBYn
jXfIyPUtxThk5MZRsJxUrcD0NNhglLYWzCykTOudntjlaLbJCNPYV7ktNCkrfqSR
FhKsX05cNmfYEVLfmDjWz9OYHTT4jx7pO17wCzhhShHcFwWsuvvk1am07Vy/paXF
6CWcOW+Oq8uwYTkefiDjDynt182gdabWlBJMSwhIQc95Hmv+e5/qOIrRE6B9jsc2
eK57Ly2ojgUysbq8nyYTdh2y+wj9gvFaPBY1UZyiGiiEpms/cI5ThFcCzXTEUvPH
1BoW6h4HGAQ/2gc/65/Oicwux84jtrCCBUiLk0YRw5XIHwmDk0Xf55prkWFDysO5
qnwZHXm/k1W2izK3H5vPN8CS+XoD6XH1knirVfDlj3u+9MHO0M1wNiDbiFb74I0s
C25whKVHXl7gL20UnwVrt9X5xcCIU3J4PmLbzKtgv2k9kLKzypFgqp2P6p7MNDuc
ijnfzf5iVS6XS4m1W9Sv3W49udM7zmuwxZ4gDnE8qtncTOBB94oumxgUKyFao1mN
QJo0mRzkgiqvdspg6i+sh9Qn7kvMeIaB7NaD08Eaw5SH8Xa6bIn/sY2eDprnRoQS
vfuTC7VafupARwhVkdn6p+jdc/nowYfq/vw1Z+mmVH+JHvLDF6bmR1rEfhkhZ9S+
ls8fUQx3TlMnmsoZFTw45GsnuDhI8sJ9asisEl7hxED0KGqmtb7Geo6ps14M2Xx6
ufUiAAVz/bhX7u7618PrkobcBpivFeVY/YL3uOlNp/4Yuqt4whkez+YyWj87Mtr7
5IpM6CScv4l5Taw+9W5H0on+8LiCNvih8OhIxw3lN74bgidWh4xVZEWYVuZb9zZ4
kp1PCSpOQQ1lWREPpr4ANIC4veU0e/q82/oLqR5jD2AZtdPJlK+1FOquuzEC5HKV
T+NqKLzsvxvukQQMYASs9CRbmR87vENcxGrADvLr54bPwhmuTr8X2j839qMtBXku
4WvpdR8mQt6UhncTnh01lhNYHdYE9VyQJ6u1f8LXMtcbiMFzDtvvLFJ7H7F460NS
jppoLl32an/k+Wja5OT0MmcFNNFlHASp2aeb0VL9EtzAV/e6QEXrL1MB2InLwDFv
FL4Vf49+bjcOt9VqK4pNwAPaUZvPaXHCcSH3tFSFNg76rNTWNGKd6Ty+TlTTaPTK
I+CceuOfP7A+DBZPwqDv5cwsuvTPHx92Rs5S/rLKMXN3dUN5njFRdeSfL2K49Vjq
2LHqOVxK343qxVq4ViSirDmVMNFz206UEymXJSUDt5PQjBfmNRUf6aMRRhUK98Mq
zNC7O2tknrDRDxjosY1Q3/G6pU+JMMFO5PiaiERLDj2yoJwLd3WwPc6N0Gw42LGM
AbuBNrW7LHqXj36UKilpbAsSuqrsdg96d171XRkOpOyYyPdE3Tc2zMsLff+lebkZ
iSz8VhX636nVMWcAyPASyWr8Yyon8OtxjnHTeSxBKE58Iitxr+dPfN1LL677dLzb
75ShDhVwB8YIYoZSb9PPq9xU2k/2B5sHWxiNi4IyZ6NbJTLIX4ZkVvitVHD6XDiP
JaY16t6VlfdIDMFvy63LJqUReJEwYIE7O14T13veQ0BHk3iUaNzA8w2d1C5xw3iU
vVL6DRDWjOiI1cfPG+75jannUl8yJTHuNuVt1QfYDYxWtz0vhu7OXc+OyFRsjsnH
6xJx6CUVfVR06qtolGwI21Xh4bSHZRVbleZwT5BXx/xX9UQiAdnutlY4C+YgpSnY
by6Mo3kUmXuKG8uf+ajehuMfnrjtxUkldkJZY5q/ouH3S7joFe76Jd8lHo6FP97t
Dxre7Vy7xugXqVMBpNULzXwOVN3Ho1KzzrhdYyTFHKflhiLgTXjhbSSAeeBTQnZO
aciCMRKUV+XqQIvHhtKKrMUqEu11rnTGykTe75O1cFRlQxmjEAvWwAF2ssOPzyDY
f3ZK912BNnxbhOsIgIzUEzXljU309+JG67iuy4KX2c/Aeh6clyqjMMi1HD/PSQcf
BqJLHxB+ThvpcZTfvdT74TKYx1nqflUjpbhKIgx+TJwl2nq75Cfp1OoXkhW7ir9J
0c40M9jy+os0CSbn8RFaSS4QUOFPsuYgny4Wln4rc6z1SNeL3iMgzaGd15hwIs89
mry6ELB8pVJBa8QhMX/j/1e5f6gPjcXpJPmfddn44OnZgokbdaI2OAgPH4oHQuEd
qVxbutyDZmo3E64J6zVUWW4CsYxSeeTowCpRRZQbrYQ3xJgusluy9ZOXd1XldyLL
Go3FD/lYNeZPeyVTnz+8K+kfmZekVbbDIlSrjVv/IP9aDJrqYto8/0q6+ShsM3Gv
I5KvFeAfiGvKrKjRMeqau6U1+ivTL8AjAIxqJWylKeM1WWNOOGXywuTf8nWXKPcZ
H1cNBpL5pnjbLAluTND6fbJniIgvUdGsPxcA2Tpz7LnqIHSawd/hnC3L2ftm696x
g48HFGmN/61jnbBtPVmyJ/Rug2b+JKY6qGGVZd17XrC76W4rLDjWay9qQTBAfg4a
CLAwTx2hJRTs60y9K1hKo0D+3GGT35xhmhbL3mmhUcdequtWLd+5FaC/jcLQpVq/
fyBrUD+fu7cdjWSWBXxVQrjfvlj0dmAu7HXmvsPR+O+KIcFILhtuUphmBxx06q2J
v/FHv7n0I3rAbDyK0RElWZzrWPUaPXsW08cmo75KAumZh5rzGh4xo6t2vrfjV3jO
rfqN4XehtGGV4kvdTTNxn90uxI6gQzW29DbT5Cp+Kx5QHjQF+QKfk4ytXaKpgljZ
TvQzmI+EUcD+Wo+uDPp5bppFTwO/OlV96iKU4dkB41StmAVcoqaC3cVyINzpl5VD
4naSQKuUq7wjF0v9UWv5cLJpQ32+FXucvXxQmWKyebgR9uf8iD5KP0fbpXWnLE0x
Wh5slHStC+cFdGMOgHNPRff2vKqAyr8OxQpi7zCIsuZsdgATba2aIoBFNy93osry
SoSs5VchyhDqTPh3ejU3WApV6FXyRG7iZRc5sXlrh/mFDAvq2MIVV+4c2V7X3iEl
pcdTQKch/AUTDl6oKItfs5OUAAWnmQydUhmiyc+8+DjRfXk+d6ERn9xnvxZVWi7y
s2RUuvVsox4VLwhHojbAJlKVSCCDN/64X+iT0r+NcNbshMVOdQyRK787JjBR5Vmw
0mRSKuQa+06zl+t1o71d7mNg97RhZ7lui9leTZMmxQiTYwj3ZH3N41XCA41qH+xT
dysOltihfxDeVPoSpItWh2w1/qniXWEir3SFCLWhKEgCS3CJS4GZ5wDt6z8LAq/X
N0nGjt1I3wZ7BR53MfeBDJj6EfD4X3VKRs2od1EK6tKU6+oJstL2uWxjiVxCkq4m
pRPQ94wBWu0mpEjVBuJLXxUN2p3MyP5znDjUdY0XximF/q+mSy11OlRwcuGWvm60
0C3hj3SCjtcmW4m/7sqPXjeBB1mnXmXx0ARijD9NJA7/4Fy17H3ErzdoYKx555Hq
SDo/iznZbBuZcXEPBe3H82eJFRPMw2irRnCG9QW08uJ4SityT2E1EpOzTBHoxzZF
pQRY1LnSkM8Vd/ag5ZTAMu3WqdWkRviV2CS5m1WUtIgjKUG9Dn/oIQXa7ti8b9PT
rGKMmgCLU/6wbQzXMZL7kl7FK+fPOXwN0sfIH1GROTmLWITGrJ3XVrkgdmQR2C1i
COcc8dwlIf61Eci3RejAfwdpV2bJnZYpGgz4avR3ycBD2edDrjlvZmXgRR5LqOLX
DnrQhs4dcK9Yn4fSD16gbsirO+Yoq8xiGnyxTMDiggC5fMYMytcLlD72TIzuRVVt
kT73+4tCo+z2FuByJDDXSzR2BKSFqCaTnW4Xqy7gtKuduub82n2GvVoZz0j2kQiy
0rfNy5BSBn728XGKTxo/A6R9fOL46+j5o8+Qen3Irs35IFH4k0of+15NEL8wmEDd
f+DUpduHHp3pdojNgGm01Fq/SYZrEgI1mb+rlKrsH7bwgcKoN6QU5L6kfIazJWVe
X356n1kC7RnR9gDEfoV9tVdstsn8nV6VVU6IBct+K2pTGKScKsYrHsqQXXXklzSO
ACiq6KvfmhNdd7GAMn7/9JoP35bAzHHdBdwe4dFzEf4K9R/PRfL8BJ4K0SJ/u/6r
yzD1P3shlxE9F/8Dr8VRt1e1iR79zBWL8wskSsInlItsRBbeQmhzfWCq425w5z8F
4HmkrCHYn0MKti3Je/ARNRjHwAMhzsN7NUWyDekXSgyupx+aETb/NEAGMMZartO3
/dvzzS/E4umzfM8oF0uaStUgNcGN24qDVXDkYVtrjYjSLWfW47rtlvbFj6VI93VJ
TjFzfY+nUogoHHg4K+SG0RhAKs6KGHffY+T1ZEo2zoCp1ADF71SVHGiJMsmJ1B8W
R8qF+tuoRjkjP2RvaY0hygp7rBPV9vb7IcpkNNDb9Hwf0CifuPUDfK5ThmXPgIPD
etXTnXMnqOeKBthIjgUk2PlLgb3ql380P8TmEM6/Xd/1F4xTLscSuMVjiWMFqO90
Jge+r5aSmavIChD63SugZbGmAGxscRjNAJWJzNPHEu6KvUMe4/RMYzMY2eCNVvnU
NckKjaDkVAHIPYyISWfF/PZWauWnMmpNF3DP1g+DkD6USEdCI6v5+ZHbhm+/2CkQ
8gcEb9ITbJsW4fxn9prn8Zxu9jm5oFs9rbuub3fRxcucPL0KBo2AR/ss0ODXfvw7
G8QCYTb4oJZNJNFGOamxSG4A3PaCIVo6EsPPWSadkqw+DGh9m2ao8lAGSQYGpGXQ
5UNuocPTqaOKL6lp5urvj5pSaC6uGqkvsbhrje0C2jR7XfLCe9N4ckvB5M6uhLId
TuAdchTpWcreuBX5HsLDd4dlLrrDvBFtAnK7ssXzK2SLYbjvsUkM9plmcqz2741/
DpZVs7pdMuF+Q+iZVjxxev/CW4lZ6q499UDS2kN66L9Hww7CmM7ubFHS7dmE/Bp7
mbvP4ie6ndorO3EnwP9cE8+/gIBpI51nWHzFmwTm49iSsmS+KTPBNqXoHlWnMT4E
ASICbT7JRO8IpMGJBrNUzzMVcZ4S/EgK53Pv6SMMM+gYh0cpK1+BrUznGh9qcsi4
afOmm3xJEUu9xyTiC62Qc5sQ938OhhTMJwPypZGk3eOqFzp8aCXE7KBoR7HFu1JG
RntmV5JOnmwn7VJch1hW1vDOJzLmfq//acBn4WvTbY38wOFWB5DOAhdUL6WXRtuo
8HJLSRhVT92S82/hY35K63ikut/6vwH/mg4wYzCxFjWtg/lKZMb+TkcweuNRKM6J
c2pKYuG0Y9WqY652DJzpLgVola+bDOOjZRRw9g/1dXYD55SYSwOkq7Yi8uvx8V+g
CFqTlMdSDYMcmsUE537OR8NZKwwSYIfLl6mZSytXV4JizMjiz4evDH+VK+Cra/Rv
a9qjypLVSvpRe81/AKgWANu4dVz4P620Ycbs5XIawefT37eSi2hqjmgSFaWzMM2v
7zGlI6XvLsFfGYS3rNV2yR4XABZq1A4q4qg/OQfgcbczHLG/f5ttTXBA9Yhl6by4
dkPOjoam80hDHAwvyzcNmeVqosr8dv2u+9aJ83R6OXIZETb8SWKOKNy6cJNL8ZKN
RI12iOfNBsHjiqe8ixI2TUC32JkSQHr6312QEQBWQp+/ahXaQ4fGQObUjhXioXQe
2UD8qFtDXdiXob0x8BCYIPvByECwjCM0LsNuZPQQZvq8Lbp6CinOHkXlhnU+FH+1
uZR0VyVrQXWJAQLKu5htmq/tiL0xCWFDkT4oha2GXxYSVSgn4/iDrIduAGqq1UZ1
lZJ3yUbTqtUgNU5vOGWUAgXAMLxKGUTXTPJX3fEcLZEuFiMfRA0/biktx8tEmj3d
ISqoUu4eckX/GKDwV91HfwF2b3tgSskouLozXkUu/ktgxkCyXt5ML1KEAOgvVv9L
AxEDAKtAL9zKSXdJ60u6bAZomwGHbvlINtwBmOtPtrIV9EWxwb0UkP0SbGyf8o8G
io7HLhJxbsyeDzgL/RckUsZiANcXukNxRucEUiJXrmV/W25NwncYgcKvAc392QHl
oXmfLy/iMfZUnCEvW227P9vxNtC39VsDOHC6H13c4uV5TFj6UQjYE9agB+eWFsfV
fvvM8i4NgSImYFw6bHD+99ewtA0owtBebhCCwnqy8ZyGSdZm5HO6WFvms3n/OQjp
yCGU9RvnWrfNlTli190vBQYFtjgLGGASeApOHzBOlbX2bl0pQWL7Xe5bzpNKjW11
bmvoyK8xaibUN5Zc8Q60gQTQImf9D+OGVxl/gvhiDr7vfv0B+VT4qL125dGkqcdP
9r1JHQdrXVohVQN3dmj5s6BolBJ6BqXauIjdr1PaHY6X8RzDbaWMOrJ2mRLa3uAz
9VFgEGCoYR0J0BuCWoRNFppQYy8Da/oODiM6Y90Z/Vsz6kzJTh6NOzSLTolYqLKJ
U6NFAewKoGpfzvYS6DfhBh/MzATdpz84+M79AufCWySEMxfck1iLFkFTlI2vqx/B
CefhCvB6/NtN74C4sBUR6/xe+slE546OZHiyTC2/qdRPdSk+UH01y7ZHhroL396w
KITUfTt3ydFBxOHjGnjAko42l4ucd1I6C20msmIIFEFITZUPP51lKtpejWpGkgTI
OFtGMszTuUQ+8M5kmSRZir8tB8v4qZbRxrAnbJhjxUCAs4RbpO1iEvPENAgriNw6
gvSCny+l9SI8katQphq3bscE2VacPicgosDqg+aJrshKBeCeYvyiYL8O5VevrcFj
X1MT2/WHW5sm2diGhePAr87R8pw8LSLcRTIx89J9X6Pxa4lyoO07RZknZP0+91K6
082PFurSiRlNwD3cXCLuNWO9RiYBJ7svKGhXr905XgZdwoh3kzwmmvhUcHupP8QJ
6v1snoaNvt4obUFZKSf5Xa9x3XbZFlFSgneAkw4rlTVPo9DDCKuT9XWHU72yBhBQ
/K2XymQoHIjllxgBRD9riysVMuQ68Xb9A0E3v7ls64UROhwLteZwFlf8/PVTa0b6
x99f2PhTE5yoLgI0QWvN9YFDl6ZMxBf5+vm2ywcoocRWLXjvQFGEleuaoW+3hrQf
Z084mvIyLQBRLRM+sdFSyJ5LTeByZa/9Mx8FC0xFQoDjGEgCGIrGO4I7d6Zf5kMT
JnZyTyR4/Ykz8FMfoxym2/KR7lViy3tm46SFFElQPsmbeQRt/PWyxghApBBj0lr1
1YW/p4cOUgtJoxtOrVx3wy5nnOCYlf8FP/tn0hQluh6ttPsdyOogG1mYaMOlYR0V
SfJMU6rW0Ft/awRC+s4uqmUzarK7e27oMTNiDRIUR7cll24uyglyhHfZLIm+CxMa
yqmdyW0o1WN+Aab5PhA985AO7lfcqbUWOD1g1fkA/8p/HSOxTI24dMDUzP5ghtLg
Jgms0wj9jqDjVNXR+WrvOg1ryihJ/Tu2cS2uAoCUdnbhPvKHK7MQOCu9+GVGobkp
IsZVoR+kGf2NW+I/aGzsKIvqGE9F0aDne4mla4nGN271pkb4QdgRp9MgbtVRXQEn
bDxfrcfS188QBTd+V73dZI/XsMTve/N6HzAW9HgB30TcMWRWBw4z1jP5HVdjp2fj
ypY0FUWoUXONe3U7sfk32+3KhnizJ3RoxKMWNJIIayQ6Jx0r7SUeQ1yPSVPBx+mD
PyTdDaMJ6k4B+1BhOpTdw7nSB9La36ZsabL+V58WqzPHbdfr8s05tgddYopNTHJX
a3TJE5613poUYodVrZ1R1MNBJzwcWB5RSe0rEGcZlZ7d7QeZfXInvXec/DHSGwJm
hzZfjCgowiAt7IMSgka3OQwX9rQznav0NdBOqPZJpgE2bbDl9AxFBObeR/lkWCcJ
Z0qfMp1hH3MKs8Pq35GwDqvHVGz7dlhbgaQ5Y6+4xOIjBhdqYw1CoRxajx4npvpV
Uujx4Vh30sH9WZ2pC6NvT1NjY+A8/N6/gVc95ZhHDRDyYyMSvyizz2pVagMOIt5t
8lrsL3f/f2/S+xwsUqEKsJR8/1IK2+Q02Y9G0DOwao/TqFLnkVF8B2etae2SsGf2
DcXzE18zURYHGimEvbMqVS08d9pSWnmAVrZSDBjQNDloFRjNpy0nVAcU39/YrMTC
S7AHzCG5NMumC3HGVxzXVdTw/Ih3OgJQpowwdCzKOB3du+wgD4AcaUXubMmVLVq4
IlVj4Y+kWcB9liFKrem8ltHOPt9ZTq/SK/OvmnCY+CJew9bwKVeVddKWTFrk66mA
dLoW2gppKd03nRZ4Y/DNoHDfEnPnDOgDf7OmmhFQU8acqaJxWhwkfDjU08sYg3Tl
T0cgUTKswd6GaT6lFKI1HEKOqe+ShLU3psE94CWxr/y8/0F2lhd0dGaRaOly6BOB
EuXvFGrLsBZjZG7tsxZ2BAsCGHREZeU0iXbpCfsqWfHSQQD997CdiXqEnonhyUut
wFHozLSYJ4W/hvqaGYReltS3iuSZHAuYINVXkxiTSUGgDvVJy+UYdZAPNn5Fd9SM
UDQkkrUkmk5L/V6utQN0G6o5K4BLYnSuaHioCaAIJ2NaGKjVb8H4qxTFO4JdaugC
8rhqtWTPAZwnTfL8NOeIItf5vddYBG9ZSB3ZR9VmPSn2tCSK9W39Sa3x8+tDgHv+
NfKHKPu+fGGyFPZyrIYG45b59hx2bJpe1Pxie65bvhU0/eDF295w7JiMm/vVHpHq
06ZTRBjoH3MFgSNYyd1+Y3Hgii6IgcZ0n3BX93GFpNyFy17Dnp9Mue7NHFae4u7z
vkAijXTDs0N9neTD0W6WN2JJU3sCxvGHfPgmJDvCAPlGAgLI9O7gKxe8UzO5k+lx
eK2NiUxjdRhsMm+reo5sLW8rQdqFybVkKsM3CoVDzKOph+LeMSaM6qdqw6YSvgWP
E19IigspfWs+p0y4Z4Onk1t7eGgdeZ2GTgOLSHXi0Z9TfDkJV7auaGzPoMtAJvLU
hZKor0li0DtpRCmJllAp/qSF1NbiFI2fOZYSZYckbPqOtYqZqY8DSUjUHLCmPGts
hGv9QER2Veja0BKWxPdJp9f1RFD399QoR6d5/qzAWflgsIiRBV3IKsygsvD13ejR
UrpxpIhGLADr+0fTlAtuDR3FkOckxauEZspAV4wCq5lxRVs+7tSGvZClKwYHtiy5
nGDBngYV2juevyEUpfxpDHMSBRjjSPvBOmpDEoxIb6ReM4tH6uxpx1FoMbMzWI/v
iLPLB3ytHzbR9NiJnXZohxPhrwmuKosyX+IFnTh9pmWuK+6eQmhvESXf/0GTyqW8
rc3nS0jAruPqALDQ0F9ynpDI7dWkfDRC3cto4No3UPiF7l72DPtoqxODgj9G1u+V
H5wYjY+RGBJknIFrRRunCqSYbZNndeA1uNhmXM4thu876WqyugWOG95E5V+jUYoc
iSH4DxDgEdQ1C7qR7LzwVMPJ0Y95bP8F8dhYR8xaydc3gUtvuu4b8DASIjtEmkWd
DzINdcVn2rSXYPUc7xVbFRINq/kWeScK+//MVO5ax0p4OdKsQnT2QoVyDpvXMGCj
Fxp1RmjgzuH+gQB/rMaY3Qak8YgTLr74RPNC4oQ8poUSdFoOpETf8h5hScnzH0yY
rjj8FYJPGSCfYiY8idBISrqnsRbgpCWEm2qzROCjyStsHLCirL79NKAGiPUPzutO
R+UPQqrD6B1Yia1IipIBKIjok27fAn5We+kpUl9NqFhcw4cJFKknw46ACxBIVHdK
J+rsDXG3KzO/L83dlENQs3X1SRcQkzRnmcEoysbjy5EyNU1VVh4ItX8mWAo4ZQ8w
+WTzHSiVIeWQArVxG5/Nyb3I8tzdKDmcEk0yz7ys0aabTxa/HvX9LsvTcrODTEu5
aa+PnWNdcmlYYaqVH0Ja76MAKqtLnbQhJzm92lJsW7ErMM3764AjBbya9O96ivVP
4wagyzh2Q+asR5L0C9ist5/K87fKLln8lkWbEvSG4h1HytuEY6cTSWJpFAWq4hGY
wXjd+UXm+87RkxSRPCHb87XOuSaeZMUKt60ZIckKosEg+FVFaIp23TbTwYxfNM91
3OfkkUS2kGQDfREFmArSsRbw41ej3+uXfOsQKY0fpdOE2sNob0a6Obs0GJjRyk8k
HfqrY+1IjW/2kA9ToRjaCfM7cuBlNy9guOV4mM6qo923vWfmIwb57zrpr916mi3B
d7HFZEhm/TJI6lHJKrAa8+OfMcqso1xK+ol6ISLciRCwoPDMvJNH5EBzDT7xmeHc
Pk1IQOSVtB2eLEo1HIJVSEvsHBI7zcoCuFTmVg2FcUf6d1t+3MxKhmVVJthV1WBr
w4iF9HgfydS/s76rMePjKM3055sX8odb4KEoOz4chTE3E6LauZxGjRTu+eAHDi9k
UYoC4mDrZRkvsKVSTQiOepIFUggz8Xh7XSQvjgWS0X9U+qsakzklDSHKojaXDh/J
YtrgE4phoivGNFIDyqF6bzVeZbIGNSnqaTSffR/2Z/WYNVB5JPQ5Xhxpiz3mqoFG
azIPQQSJhPpEM84bkwOgzsts3cNObRGoW+weJ/oqc2eB/pcDE1ehwwkZa0+nvL6E
87sieT9PUCZVGk5lwycNbfFNgg+B7rVrtGvDKITNsywVtgyD+3H4B5SJY19dEaDE
C92P0b0RPRnYnRWUHjCHWC0jOzHafzzZqZ2/ZI46CF/EUNqYrBCvil7DPgpX1ZUh
CxcB4suLBHyREM8vSgdQoNOYYGRRaG0JCfr+Ic7TcgknU7hgCvRNdGClsnyrZTCN
XBg7VkOHbbfZD+GH1qRT1VdNlgtco5iFmb1yk3f9sHn+goRKEtO2eJxyYgZlZPw3
6zbwvXaSqlehSqNokay2kzzUIwx3JK0VoDe0l/BFUOONcf6aDWEpNzsPXrT5Q62a
odL1PHXsJoYxk/k9S9ARnjGxUVmh44Wu1hSJJxcrEI3ePpU1FqwNQwvMQARBIbiO
iO1fnz2KjrB7Rzj0AbneZAgLb5EFgJcJq0mTiQpY3YYoLOCDYJYDpHV5DjM2fBTW
BEuPIwKbl1cSNp4MVrzcUswKk0Zoed4nhZQvnbqEyq1ar/Q12y0MSb2SK9Sx+9UD
C1Y/fOOCCSV0CQ+k5DsVfAqw3wRbnQ/PszgJI2xz/fEsJnIbxvWYLXzE6SJqrLJs
NGOLh7IpixQiWQicO0AWfZRhtJTkzE7c2AL5RCu72CJ+JYgRgCOxPFfSXyUdYN0/
gkoDH8gZzYKrpgDu6ao0sEz5mWR0eoQmDyWFo6zJjGCmNX9rv4JZx82rP2Hnk757
reNXGPD1JqVmWCjd43p2Q/TtZYM78m4aE0cDVAwKx4MpOYbbFOAccH7D+3kpeTD3
eo9nwX+st6z8o6Ysf4cSKAxHF/V6iSygKKw8oYZgdcof8KxF4X1RAK7Tw2PaxqrK
6P9pBCun7bZjHDphpEw7Z6hFDbZmPEzvTGDjOECfKrNTEHcK40eFRhPrG30jFl/P
YgmZn7LPd1jQNotqHetqb5yOG+DzJFIriF4da9qdFytPD3c50r5iy0BZNkQKAGPe
4yJ19vmLXhrF7Uo2g4nDsEeXzYwT0DpAHWjMq+MvEUvrHBzCvYdrRvmalEieDTwa
GMew+W/bKKL8BeJ6S/rQ4Qpgnv7QIGSUHWG9kd66SbTscoNeb5VSsXawMxur5Tir
KWPYiK58QgGCrBCnOtEFFtvZjKCTCELYfTyXd2k2ZFRu6XRYk63V5A/GXX6Msep2
26hHwwpxNVOKltH2x5beYwrbY18V3/lAnpWLQaBsc4Q+MEmDa50jANs6jUOLbE2p
u48mnnxmiLrF1ZVGbZgmiKK71KX+iTNz7EwLpvQQegayethE0QV1TbDZsHd0lnvY
PrQHf9ERCSehx3y9rRI/rf/pC4F/h9Ds2Dr7NTZ5/8DlyIqYdvqkSD/nUJp+QRhs
WjeD4Q5Fw4cDS8SL4NRMkWU/+w6On/Ogi78Di3qL2BdBmF3hO+aaSN4pxQSOD5F7
3CAQ18qmJIQRh3xrbNG57/EkXrMUHnV6RM/JOwUNFnwX+1cO6W/pb7/3rtGEye0i
dDYwgJ6uSw8ughNfixwHg6UIieGU+mCyumODq4oCwwBEk+bJtxQK9YF7HPuJovp5
cJwvhYgmYFKhoV/+iRw1IQcCUN9vA8MgjEqGfrwLyjXOyWhZdka4RohUlSTvwhzE
I1RVvD1oH/WYv6NHEk7RGkreEVmMREukaTZaYdADHxbjW+VITSLXchy3HHQ2UNzN
+H7/qJBZ3NWveMiV1+Zavjko8cEd85dE+D7K7CMfHvxUUcNDlivfuBp+T0Ez/K/L
BDsfhGqSIbdj6ZcVGz3imqIWqy02XKyWuV3omrgGZ/RC+a2qqqNGrm0qxJK6wHP3
9rb/xc6xQXnL8Q04LJpzgOftcOQ10b59yqIExI947SXAaua0kz4CxUVDHh6KJrzb
9H57prFkb9Kn05ZVtK8wUYP+I5lcd/u3MJuXTQ1A/s905j7CL6Eysd1p+Pdq/3fD
7r7PdpBaCAz0M6ronqFnmLMAZAM/ZlCwtMV2QTj4QzTx/OC79P8rrg3VgsEYVW4L
0zcmeuDRJBF95MxX9tlZ6EtpigObUBrbXCsrzubekpjbBGz1pv8GS99x6ymNtekr
jdiCPMQZHnwN8qQoI+9iQXQX+R4Smp7dkJ2QK4fj1uocMTVTxFRUDqKGYqCsA0Kl
B9PtuxB91a4UBwQ2hLIWhAbt3xzx+O+PioELCKMA3PaQCnVGJtSPK7U/mtarZFs2
pXqgXfrcqaIB/jqyypdYGv2cKEnzr5BgfEhgPEDFY5pkGQPythapkmcxDNnYH2bs
kFaEU4WM47Bj4xSHDX4+zhEfQ1a8AvDyelzxxkUewdwmZNS3a/GB2MRUfX6ZD7EY
8kIp6mNWPmruiWU9WnKofv063MvJ6SMaehtuENQP73vQo46N4jIW/YD/NyrvYq7Q
dwAceO8NKLrzAZXM8A3qJR8wq3FrSEhpAdb1MjOSzJ87DDo9d8SRZEMQ6YdvhG0d
aSozJNj1UpFt1U3zkEWYSNhZTR7PV7o57sf0LBO5ryLHNfNcBkoRbqbiryWOYRC+
ckuErG2al35bnfci+wTaGDO19M8okgetEAlFPDf2FdhE8ee22d6pLUYSEE/WLgKa
hiPTAQCQBEYJiVB7YvhbAZN0Ac4y7uMu+gO30IOtBpCN0f/uTGeE7XUNMKBm+aoN
OyPFC7mCrH/1RugF28vh/DJMUT5P81VRlpTxRorJtF8jYdJCEEaYK7+y29bdFdlK
6HyjwtYVtsncnt5ae70zPmYS6HyK3z+TQ+6IHf7Vp2co2b+KgiyXcFf3/wO/ccMj
A0QzL8YQvCpwFoL2qP4weA6cbi+p592a10/brxd91ox4JwWp5a4DY4KqF9sUwPml
qDWTc4E3DkXSSx+82vCv5ZRMYxpf0HTX40xTdxdipDSNwWUWwmg7mDaszRXWVH+E
4goaijMJigYguBTenW9NGW/gl4RU7zTx23/LtAyL1Zc4g+JyRTplXiUC4PwcP3uW
gBfEmCPse5Zm2AWLekJhNXaDzNe5FYNYc6QQd/L7xo/c9byij/q4ViLNsS3vqXHw
QjeQtalJmfi39KimuwhuTSgtMQJ4hvgu7Kz0isV+ohy93TT+x8edCruoTPwCfPrr
Rj+QVdLolM/RxONvvs6aRosGNkXsZetsq6V/1hsKZrgKNZo5iuB+3pHdlunALcPj
smmQodvAarQL5tocEklBL/3cWeeXMod3y2ksxXebXOtGWPfclGqY9HZgxGBE1VQ6
nA2zd7htQ3E2ilQGELti6AhRHmdiYjfpUdBF9ojKsPZ+DBsVwPxOq+JkJ2suQVRs
QZOu4HB7ISoWYrLMHF25AKfjrxun1TtztMRXvQT9VRD6UwyIsn02xM0tLkem/Axi
EIp9hvAZoM2crWo7E7mQrE3pQQE0++UVrbbclTdf2/TvKEjGnxGttW0xS0iJykEg
TzN0D8QezoPRsOSpucRz+leIxkIA7JFoIXBjvXXDxMBUHtIVpdr/P0E9/2smVCa3
YDjIIU4wJn9vObF25G6mnSm+aw976oW4VAVWNEiTkQUtijGTiAgMPpx7kkSOyNs4
gH/SNQxBaloVzIGfMJ6Cp+FKSYyO+fucy7cHleXiOE4pfAcSYSl8MZWljFYJSCYO
0xdSExrM8rOylzdbsMvxk0B4i7ov6bg4nMAFfHouEaNTfNapBxUS1O6alo8gqtC2
Ai/L6YehW+MfAXhZt8FIjaAy9p6P8YOk1bmLB0uybDsLld/HMkmZel9k5AisoMZ4
ARZbE569ZszGq46m0fw7/RKd6Chj4RrdzXzQ/Apuxe/L6zVRUCgnDtfhAfmg5gao
dlbogZOEUWR8qrKuZT2hntGaOiLhp3OuN+iFyfrRmXDexyrGB5vdiWAQoOWOm+iN
DDTGooutwfWuqf2VFu+xcFRlg5GeEjDmi6YcC2BUFdGQ0sTtWBl8V/XXRXJYRPvO
asJxsVcmgVwB2IhRft6lzKIFmJhH5Q7PQhnkFXUcRk1foezc5SpZAzDK/m8iH/3r
4u/1LFSi8C2YmZ/Hon0V3k8CT596wX4D1ZgQ2xjZMBzkCoYJfVCJIx8TKZa+hbk8
jNt+Vuqc8qvUxQsCZasJNYKmkMLpCwxTsX0QH2PehZJ0iC7z9HALUYtmYXx8E1xv
M3jX/y1PO7gVhX57eC06orzTo2F2DWCmniGbcCVHC+hajP6V4Z5LmDqT7HYjKVo6
JAhPl9wyio5ofM7G8gUMbfK1RebQJlcg5RFfqlSyE67H63nXFzONcjDhOXzxtc0p
SEIz+2URbD0hOCrEzCSPjRAusBrbeTrnShzzYzpZFW5PXD8f2ObvhAsmETVZ6pu/
4jve45xy/msWQ+9mAYTXcYeeYn2t69cME3tm9vemEaWWMPBcb+3kitwKrl5dwjf0
V25g2xLqfhjZEobW0O6jSt6NyKzPyGm987uOsEJiQG/yewHEvCLwEi63aiAEDp34
WjNTx2cNBfMuuWdF2dNFKh/0nTmrtxC0nPqheFu+FCoppvIrYjThAKOFsETStZg8
8i1MauHX31Ob3Zq8+SJyLB7yzNTN9NvzAu5do2xHhL4zL7ei92YD3Ou/dYagJRob
uVo/rp1DGbcCHaPMzHDJXwlDecHJk0oohU87hIBz/iuTgHW7xFfM6lKrd7W3bXTU
BE2be5aAfLxCTMUnPa16+7oO/qedojLAFIxvDqderi+oHzusBK7JPE3tXmdG7PmJ
Jkm5fZ/UNB6/aXeKLNAK+VciCn3BjI3w/7ZFIUZhBuFQpsNajB3KGRlCRvM042QT
h156VMMyQFxA3SZeF47hGCgUFcMKeKKsaQi5iTAbNOanvPv3A+cmsiI3c+OauV1q
yGkM04YT2dPt8sMvltlUWaXDcPnRA/o8mQzz55rz7Vq/qrwC77Itgyhq5bHNgcwW
oPczUdYZ1991VsgUzc8KSgh3CJKfs00UCzMHj1gBGnrkbqGcxD8kFIma8pSLg1wR
Jzfsh5gFIGtgDjtsIQcz2dIZfb8pixrnrMJr1qNQBvMg0bjbjcn/hjHRNz6D8ThW
UTkppjFJHUs0HyTjMU/FgA9I/uKemlGmUHNczG3LjcIEUGhKPekoG3ManyOv8Kmk
QnEOqyH63CB9eP6YV8s75y4tSAPBp74+CWmqK0R+9w43nDMRY2syEmFmXGo6+9GY
78dCwNMPhQH5nk+SdsgF6iNaAgSYYRtDX4hbwejgJNTvlnd+Pc645hRCxpwPBVyb
Fxj/OQctISyn8zB3BiDLD+VER2i5jGyQwy4hMu3fiwRln2SBN1mBtebcpSSGgo4C
e3IeylgHw6DsrC5c8LRzdc5Z/3JbbPPiqdquBC//AMZ0r3xeW/tLDSZ1hP4CTAsl
T+KTyXGr26z1toKx4cJPR6O3H/ddo/SEQFYIEOreceh754xsCuyZL09vbwrEWrzG
a51XSc8keWJd9gUn8RqEb0psqcSbq+KXGQ44Adhi/ziupO/oilVqGVUGH7gVU2K5
zT9i9Je3LReZ8GAiK9I2P0pDw9QSnW8EXoNlrVRJDlNaIm0OW9gj6aK2/gd/6Dyn
utAhs5MgS6wYk2G04EX/gQ+wryHPx4IwQzwrYqYgnZUV7np7qo4vaC01P8RVFoJ5
svYOyVpfnuhWV8NFY1TmslGIphCk00YmAsFdV/rpi/pfwvHfYG/eoav+HwK7hUtk
4gzdMaa38MR9nWvqXbqBEAk4ajanCOxPKYhDBEZZIrnbEfQuH2PCxb51zcNJIaHz
55lpcZXuDVsY9QJLFxk2pJ9DDctLmYUSkgBVR+i6pccWRHyuglC7Cgdx32sJzHVS
B5Dh2ghldvwa6+oORgIttPdpK9UhRwPNzg0RFBlfDltCHyJ9PBF1/tuLujWkyVWO
S/lFBhicNC3VZimFjViMcH+bdLTMSHNtfXaP1dEsxo8D3pTeuDHzKcmk7m+pXp42
p9tUsJqYNovOmpLUCXcDdiKXXHX5z+bmuHFt6MVwel5Y8/JcnGLKQQwzyJq3lg6Y
Jp/jrAugi7h9oRSp0I29xy/Z4ykh0NNBacIJvErNOsjpfA8eH81XAB96SBYmDF/7
euF8UoPkbLSepLcU9BdbPqZ9G45b3oUPSIEo1NvO6Iz8UAutfUfpMyd7weuvV5pc
1+hHy8jVzeb6Z9fn13t1fCpPPwi96Ok3hKtON6K1F271HFzavoygM9T8ehP9GFoI
N4K8q+Y7d6DnlLAd90tIY6jtvqnPcRErCTwJ79+kcGxrRYmj9FMklqwu9/zCRVjz
Mh6oqWDK8Hh9CtuE53Pi71AK/egla/L8zWYDMauWa1bkn/qHHD/nRfUgISbj/FOc
watXOjfN62Jbh4HjW2HFnlAKEOts2FENOwvszDMHIKkofFsbiIca0wnSi27Sfyk3
vjFdqh19Gcegqs1Vuf2LSceEvpmfO48nozEXTSEIv7xKz8tEDVsDqdB0yfP74uwv
RI9yCbyfdDO0is7nnKgKdxNRDzb+2UORBsIDeqLoiICtrkHXWoeM01mWYlGncADZ
JC9WsQa2euOA9pxIKhhNAqbGsY4W9CU9HcyN1nzQbZ8k6CSbsC0ycYUHyGf1y0mm
SStD3qess/bpAJiUAlLLlVIeptgRNzEZjf6P2jl+fcG190kMqtXfIH/DuPlUupvH
fIbOc7P3p4c9lgsb/5UIwk1lCgcX1pHS3W+V1kx+4/MhFpqIHgvorsJ4cFgyqcjS
rhH+v2KEGlYdhZi16Xq/3TsNXyJyEvKt6ANO2CvRRMgCg3D6me4ax/HyYuYm8J76
BRmU8xog8QLWXpQ12BUOiz86BrVXYUU8BU6ihayFWioFB1u1nl8wVJDzOIkyw1Ov
7pz5p17IVJ910SPpUhWbqcmCRpNnKbScpJ8gfBiSovHEcQQyLiPtAyQN6+6U9BwL
YzGmzQpJlBJmZKYgxKNpt7krhwoL7ijYEFOFWQGlQOYLnDPDGWMzNadlBk+FuBrl
URB/XFb7p8aYMylgas5ubE9k1atdxb1q7W2ocKwVntl5tK6MBIijfDZFQ2Y3ByFB
ky9ktnMxZcfpIVHOfYcFBM7zht5Lv3wg+S5j+3EmjDQGJB0DviPcsdRT0SHq81P9
CSkYaiiC+Q/kuwvyX4IZbGs0k1RQIs0of4iId4eMvpaF4kuGupYDof+Qojpu9ziz
nQYf9PNGC055QuUphWGZJNFjpXqVYeedGk2CJ2nelrrHnUr9O9mRgeJCDaHEeq41
daX3OzV/1/2D4WxjE0FhTPz/cf1RTgerXIdPluOB4coeATy+jXP2hZhfy8P85SNC
ijugPazdX0SJO/aCDVx27OLFEFZRV8GxY4ipc0r1dIr3oDUoM6MyWCajFeZR5rU3
Q/jZirsiyfCVylByfPKgA1uJdQSVnzfFaZbXMg/Mu37k0P9w1qDckAQsQFpRbrML
FluYkziCVsnzV3YuQnwkJO0BBpVln8td+eEd3Z0yXJ0VBy12IUg6XAtnPkRmOquy
gEUNqszWcCQDEBAkqOF8LMtSjggSLLV+UBiUFqBr8E9dSf40o0lCDfMllktpjzTo
1qIuENmiTiF+X0lpThLG4oMaGtahTyA37DdwVEdF7KfYwfLNl6Rae5iTN4ilYpql
kK+vO4Ogb+2/a1LUFnO9BGBQi8AEjvt4wpKr0tYK+f33hIlbQiRwEzGDQ7S3gjFs
T4E1oEoPm5ybJIEQlUKzvzSuxFMryHJ6UX9oXvZLUgq8IgICKMGRKUMOlcnwVbMB
KvYvRvelwKy5ksve2WuuwiYgYRfAjy9PiQJ3eTzf9K7XVDfYVgzKPPydYVFnZk5c
JgaSGLIDh5OPyi84X8W9/9/4BRYBAQ10JM6rOvvJH7YkSx4FR9zd1WOKf/H1khWk
Rp/LsSzM53fgIZgMNagyzcRKfwBw/O70CyH1FvhSA8v1jKT/T84mFfG8etaqgibG
odgkpXwJCVmiY8h8b286rdOszwU644r7ofiT3mYiMFdzdMawXbPuQ90H7mZkSfSS
MbC/dIFQdkIgowS56gOiL2OEaTLz/mAUa5pEQucjeM1byaMdaoWkWLQXqzFKcqu8
aiLdJ0PfGGE6F+IVQhLxRSnu8onQCXIfiA23RgPHneE4v+LxJ5QdH3frJfH2mlgs
8a/NAQDhh1PJMxd7xS1wpiG6naokjzMVxJk+qOYaPe/8jua1yVFPAVg5e9KzXb/5
wRAjhD5t8cvJOx7+VqLqKZTZ4f8PGhHTtsrkpWaACNy/atjmn50qikddAcTnCRXa
Ww/MaHRuuLsocT9soAdFI9QjDhdvWYfB5sWVSSVquo0SzXTfyEwjT1MHHSq1sgQH
6eIQ9yflLQa1iUgm4AytnqPbK8Ved/ENo/wx7uxM+SXlIMK2vO+jDsxA6GOQL4bq
+J2/MQjK6sJu6d3Tt34UAFP/0hDoeRg2NBhmQ3WtP8SR1P0nUZtiwi/RU02Es1WH
Ox6SJbYY9WR+TIgzYXKzL6L8Jd+J/6rwA6jQiB2TMNUvaIpxZslCABzt3ylDJaii
HM5H17SSGAPjuRVhfHvEYbGj3tt9FMhFlLPFU6sThHs84Bw36giU4zZy65X8rsdo
Pi8szggsXb3keD31R7NL/4Bqw7vIwmImkBBe0r0IuJHC0rFEGwT+CjxftnWIgW+p
qmopbp6VOuLMX+9clkucmPhZbiKNTsRlpAK1rtkKha65uhOvvKwSUre8OZxfadai
w75reY0VF2l7A/y4sbgNWBWLYKfGzoYEz4FjuXQC1XdzQ2XwYn1tsYc35pkhWEZ7
p1YhFtaa8jThAgGjGAH5z+AwpT2TXKC2tjuXeW2gAQ6WYzO0RV60oLYpi7kPbg2S
Q+Ju4x9R+txUUfWd1TT0xgC/iGBgHjPYSFtKFaepZcs0SqBcloNZLGEcbQfKAdMI
QvVBykeYmCY8bOKpTSmGbWKH/MTE2BvN+tQawra+Jx2XKI866iLXokOG3LeRK4ug
bp28Nz+9VtgRA9v+rtu/+zhPdnvzVX/mz2F4LfNHQE3FahO0uVjIJPo8l94CMs/9
WKM6+Mi8Frl6Mye0fvjyq9FyhRBqzL4zdc6lTJYDUhvxt/VxPDMLioUHaYruMhUD
uI6q98m8D2tKE5uU/YWLzG8W5+8KM37kLRF8BuVNu7MyfLP5WYsm6w2O19aj/y4Z
L8EwebNZeLMPPpBvJQZBMYgm9C40PhcNzoLT5SiCXh9pefV5p/4tCm/7QA59zZhM
jYo+ymFis3ILtOF5S77BjNTf+z6oVxP/W2wYNhMzBaBbJOThzsBKuHbnE5qvKl0R
yVFqD0SAo69tYX/3tWPIfCNyUXHve5uooC3yzVJKu6YLha6lkZY90Luk0xoQLqio
WCMSgjjg0dBGHrajxh6vX/ewnQnTxm3OzmDVOr2BGfZgapp/s9MhJcLP+/nbmx42
s0UI8WcWiiexc1AMleKj+AlVJc9sXvnGG6Rcq4lmkbhRqxwE+dUJlGBG9MJAxiCC
ctWzUoTeFN+F2jk8IzG+f0cQDWoec0WGAjeZ0glRLSiqkuVUZHCW/XwNX1m0Uc0H
jzR2dkhqiEQ57pVXjrIY2xb0JBSisW9uDVMXSv2S25sOuSQThxw04XfxDjtWXBLS
8p6TlwyFs6eoH5eUvONFRFKz8gAYgtFgdktZCXWbSq/jCRJ2w8MKnvK6FWB6tF+B
VypiLNOu6fj4TJlaqEIWboyUnWSBpAwaDRIfGOTvKzeRxn748sJY7f73riAX1pdn
MUJFokJtuBqMOCuuTJCKclqpC2zhOVMuEnzBTOeAxuTfZ3LZ4QkzVhUBI2Ri4ksV
BrvhsQwNSL5xMGo6vJRaF+4YbrJDEr7njHHccP1ZgqCQWJNjx3G+AZ8I02qb5lHd
ZMPqn2u2X5rboTHd14A8w6PKbQ4JMA54NwkjVvHTmjVS3LWTF+5tcbs2luOiDSk6
imaIWwGeWAkTpnIOZ7Z05izTwB6XsP0WAqpevtIUU3Y2UC8FiMwSZaHffx4+6reZ
JT7w+pCASCpJqFUGkWGifcfNurjvGQn6J2+LXPQyaAjPiJVixWYJQF5UQSGzLO9k
sUrlipvE2Fz/ZKR5ujKoph8FlAar6gOEIM/jt4rWn6Pn5AUMpEYthGpDL5yvia2a
jYxib39CwL3wmCkUrh+yyo3hF5F4Exbgy/1E6hJnIA8B9xbbFBEMKwDoovQY/BLD
/1OCTvclC628UdAjETCIcI2etMUzMaBO+LdKeOrLuZtWkprW5kqW/sZEvoddv14N
cxV8VPlc8sJ1CTeDTISnCejj6QXJlwAkH5ubvVRC7V/XtCx52Ypt5JHI3zGoi101
Xp1B2koPyqcwBdbHiGnRs+Q1BWyiNeN6E1Y0Wo/L4kOcJ/Ioe2QAOZPSyY3oDSLX
qzG/dPe4V2zwe3+yZlO0zEdb5AfyBw7MECQ/KAYSj3h7QNLqocXL28I7hE/ICNED
JHyVPFOTlJYDO1Uw1O9UaOH0vY2VB6JqJtVHS5zE2NCKmgvBsQAtP5vJ7MxGno1/
qReJTUxllPD39UycQKr/fsjNlpSnvCS58JXpZfFFKIfwx70zbMxdvBx9EeJe4Nv6
wfXchkgnHNPRcE6+zI0gVmg85ME2d8CwWxAQTSZn42Dyy6AqyGqJo2Vs9tBn8LyR
woVAcbH1r0TCU7HXCp+ODB5VcCTfIkRDSpLSRNGybrwDEi6nYrpusbfARyX+YPKV
MyRMmBIFaI7cUyUlHqtzoJ5qgZLZFXxkV23LBVdHA/lzl9rSMTFGdbIq3vHe034Z
UOg1zZJlxWQgbDusgEzMyE4c8ofJhEPitXP1Nod0gIh5haiVP/h/TbQNWUTTKYJf
desGEKpOSMgu8rEYxOtJDu2i7KseYsKgXJW9jRzhob4gEc8C/ZErbmHOixQ+9B50
Bx79XuqKnhkqJWAGOGmGHDQf0Kk8+GAiZANXjJuiTdXnP1ZCTt0MuRcwe1z3x4PU
FRSjtQwl63ZsBTIm97MZo1Iy4CBLQ6UZUGiMB3E4tVPjBnGunz6pz/53Zzr9YyjE
30MFzbhrmed+YljqrevDgPw7ycnr990kpvjMibcJ9l5+4I79gg4KdaKPP1SabqTx
XtiCfNYLAXIcY+gO6GzUMA+lxkDw/NDUlHPQeWI/HIq+pQKtq9qUSeTMrMEjWuXx
+KGj4k2FLaU9WhgRlhLsGqwH0y4zqCXtA5br7Ahd23ymxQkImSAFahZiKCGY0IOd
ipz9dNdkxsm+7X3SbBBfmYn78uD9qd6Wko8L1TAeuLieyv0u+AMDE8M/uqcoic15
jfznN7/H9WOXfzkpodGJ5b1F7Os4dW3fiG45Eu5SLmqvhC9I84pACi8dZFWq7Ca1
QB1RbrCR8gRPFVmSuo3wWxIMbtV601kxNK4801krvTl+7uKOgDb62cAaCJ1sx+2b
8XE1ErKj+QdhZbXhUHn1Cvamh9d7xhpPDccCFVGmyzMOpJq3aTtWZGPK7/rv98LA
VyDQj9C0odty7Ux9tnYgcXeCx/JMZH2QYkNpxfk7vs/ka29MbNbWIgR+nPr3qvcp
6YllRa/k2Glc22UPahi7iFsAtb0Yr3Su9mK9WmTB5v1nItAwTSZF4+VYSUDubirs
GgBVeBiBjW3lKxNW6jep2gR7wbTMJWlpmuos2qmu5dl2G9ok7zkl4hgvPY/yqKBT
Re6hQE7wXK99Syd5m03Ml2BcJaya8OibGyfPZ7iIAnLq+u7V98JKfjn+R6WvRyI3
op2wiByDmPxTiJ3ORrpLOZNpiZGr+4/o0mozWn9MDPUII+7WadSI3g/6otnutSy9
18i9jpY5+2999y/Q+BfKDjF8kca/pRKMpRZabnwhnHAQdj8lH26ZuWhPwcVQ2D9t
kTZWo0vvv2rZtPHd2XI4sE7BGcFL1ru4AP6H6r0jmOgKQBdPZyl7Q3C8yiY7GmVl
um/MTV9ePav71PE1fO/aRdvqkEvKA99d55D0NLmexoo3VaM/6EWnNssLnqkL1BsM
GCUVvO2V82ETrxFZpI6CyPOc3qS9tIuVCF6FV4u0+MWJY0q8H+iuicrFrhiQD3IE
gQG/sivYzMEEsoXzn9nXCquo2BKq6hwZJLF4Hcww4wYYEJkVEts6KbQZnDX7Vr6F
/xoR1fc8inB432FjDJ0pft7wTOOwFPM9IuvC+2q/0tNRUacmVkoP39XM/mwGh/ys
bM7lYAFlEal/NZ6+3/Kn+RgCZSDSQ5k8L/2ZF+r6OfipVyayBKHIXvx5aI6z9gsO
uYylg1h2DHfyWx/J3qcT44YUnrZybHa4PFUoByNffB0rseR9gNjx9ttdqvNixiRz
/dcqpATULelgUZqamZCxeNPNwHQPaPw7zVp5IPFm47KjGTf/cAkxhSAiTBJ46HDE
BUY6UDpijL3mST6VJQVkISBRzSasX28owOt4evzG6sIMzR3pllRkPGLyaHLEjGqJ
sVD/it8ru6frnpBlxShix70TcyldrK4h58E2XpNItRVvwbDgapUExM2t2FBH3Rk/
ZMYRgtwklcBgObfzJ5CZ24eOVOGTERZKjh99fab5m8yJzJKjpEZsfBesoh9qv8X4
Rjes9eKjYle5jaF1+rUs7Btpnn8bFpvTeuNZuTuhhaxFMgc1tHxeHJAXNNvQ2Zp9
yAQGf2Ef7ilL1D9GWPUcHF9scnLKg3L+Vouy02l1uMzdEnQSsoL3WtKAM93jBevl
kCRRxB0wFJ7J+N7pWsWZmdeg7O6E0osDAZXw9FlkltX0LEesUArrlGm4bAgszLhX
XZff3ai1H46wVYTKtGDXwguLthYb7QAh9U0yFI5sFLtzDrMNuznzOdoZzcB1Hadq
g1jfswUy5Y/THkSR4ocxTYrmdQIoZM1pILC6YELLurWJ0t7+nahRVQjV2g/bYTQU
Ma7IckemMqhJ4JgUSyU9QTIf2tC6jge3vaFYHJoFh0U1kEsOlkRumSutDMkwMY7I
UBWM4CF8rF4dX1GMSKEfmhsMdNPl0azmvjYPGhCNS+8uRwOdfuTf9u5Q8saspbkV
7qMuCJntUbCYbYgJBvr4SeH8QRslIsXhipV3ODhEjrooslnIQVph/fvALYKH6e7A
3nTLvL8+MUQEzn8dkpa5xvaVq0n0N9QSnjAM6Z+SEN69Eb/5A9hDscbB4rU9bsor
eFafyXTEwVfkFZg9PPmHVHq+ioAzSVumjsDBBRMnMGwl1BaC8B4EhbpRwoapfYzf
6m9F+8swyxeZrub+HRRv24CoJYLS1aKbb+Gg57OuTfs4z8FKm9F0PavuUtOY155b
RWDXImRFtgWko+qir04eaomtpa86yDt3ljn7w8oCwv08iVVRLPksXfEj0HcfG0xq
fQdS6++1sPb1RnPM4Q8JAISf5HrBDUfNX6VR/Be9Js8E9htTxPQOOqjUpOYvFK3x
/txVSu5d6L04IeuZjrGiLQFMfIRZumX9uFoGVy9Ne++5VsldlyUlfAknRrn0uddP
T8ObPK3I/GvCdOgXpNyGKE/ibrNGO+0/M0yPbWhAehJ1668nDHvXJm6uDvlyrJ3h
+Z243hd4cQVuYU1pGWNTgKsHtUdYmngjyDZEAFnecKoTMyjwoKOZaQllEHKn0pNf
rOHaWlG+SpaVncBDRrK1llKRdEPGsqVzGDH2E8dMRIdTAC2NPg2SyDU2X8Om2+Km
XY17cjpZNWZ73OCGw+M4yjafyFx0YmKRlrvG2YXJyD7viPhI1VWtzDbbasYm7gSC
RyOKbO962eMDKTSuZzaSzbjYCyNku7qlPnZszeJvr5vjce2p+k+KVzSqsWj3cxL3
UU4FYTgQSrS3a2smkCM/HnGuyXNQ+HUckOLxy/FTCl8FfWbz2WbWxeTbOMj4cYbk
kVYZoo+hVIuzRP/9j5wwPRBdqf+tpC/zUbu9gY3jAjAFo1ypIlZNwSvIBnbtSTEt
jJKrneOubG8pDLcK22AEqLG/KfTmzCihF5WoFxHWgvl43LlEKKeR0QqW6+6j2VBy
oUA9EReMJ8IvxX5RaFIWcbJlgUCst0Zpge3f/VNYXdOVwcAlAQDPz38b7ZOTYRzw
uiK+HCok+ZDQ9GSkReERlMOoKcEPwOHCRqEJDi2uqPFJeRoD49Vilhe4seN3Y6Ze
O99L5mm/SoZw2oJ0RcmQ4y7Q7zNlEQoXlIedBpJVSr3eXzi6dPuMrEyktRa+st7S
02jqt+1k44c/2vTbfIiWy+nZgdt5aCxT91cTfAAl64w1fjusUkRjVTQYE++zZpLU
Zwh8XsTeIhLrBlJ3cS+kSOOGY5haI2Q2y/WfXpPbN7+8Hqqli26mIu3scsQ5JmJX
Bzg2gjAybKLwFocWykh0eoTxUIGjJst7xzqXVk5ZovJQuQeGdetgw17SKKo4KJon
/TnPBL1QG4ihy02uFbUqhw9ZaRA5P9rZIbi/Mphz3MaLFbfgtT4xtVmE5tKF8L+L
U1VgudcgBwqdYShC1KwcuMQc+MPVzE1n19/Z7DxF5EYzS4xrRRmA9h0TBLfxzmUK
g7vaO1F3u9SMQD45RlgTI0fo/4Yl+NSoWZJ0oTRL9Np2xtnCbQ6zHmEmfw9HnaLm
Iykd0XxwlXw1YnVm21W9MvKaSBlFnCUXh974jv2XN1Hd6lJMs0h5jfCzqXlSXXsD
pBoLoAwRDC7P0d5qXkxR237quECEpdRfwrBJ0bV5Nfl1PEFjEpWoCvd4eCNhCWss
n2HhTI009ZOBFXSpPcj2KKSMY9QK2/lzjIx7HhmwQY3MetZpZFv1tT3jWCX5NZZM
MncdtukGHWYxkkW0NNrslcu+QphWcsGh4gWKAYpQ5QT+LSSenPYj+9a2xFyl8hUZ
iFbJeChxclVyeHhvrFyQBX/0HPQk8k+uwXRmPQjDnNs+ia6RYjJ8ACTuiMCU0WD9
xbRLVC9XXRBBMUWyBZuT4AvEBjZcLPTSxUkGyjlFjBoX5CAGKwS2zqYEetoru40T
xyBvvrhwoioe2fyQKU2w79sSEfUurxJpuEsKO29dRXnLD2f+XmA9RK/Rp2Z5p1Bl
bYPJq1cJb7JIxoO1oFFsi1l9FV09A9NdyxolQuz5WIfuQBL5XA3t2IJtArps69z0
PkBfHvhaSf8gCRLH5Vx/F9NyMwvwaAlGso+YnyX/lQnnF2G+iQJf22idGWm+F1pb
yM+kRDHsBaBWJUeUZMjBFYuf6enHgsVUPyuhaTa645lhUtUrFRp6v4ZbJZmRDi+O
PqXKRzlxY8nbdWWrXkUbHfCSJqEbpivamXS5cJtPU4rYVAE+fr4Z/VB7xJO918Ag
JRSBSepVO7fwNxLbOhHmdcTphzLAs/q6kpwXynqzGfvg+aoi6c2msr+L2Qs3BS+9
PN8SNbLodF4dH9kdUtODjeoUicCksWM9JgHGUBpLY8GRcyYuto1ngxJONsgZG9vy
Ad9emGYmsNCvXVu+noVx5LgwEh+up73vQvV11W2/dqU2wfGB9xAegNuaH/HKgv5l
6HfR+5DgNYSl9wFB7ePOw16Ix0fbqBx4X8eChmhKgV8ldxdBxUwVV2G6xwNCSAu7
lBxnFzDRBFleDCxKdfpf/dB6lqompfPxZNq4c0BUR/YzaOqxFeYbqSfcMdswRrU8
qO6gINkh0lJtaDT1Wh6qz98X+bJ1viUFRE4g0MXh6MSqRBfdrCFw5JVUS0qPQVZx
2p9IVoFO7qume6ps765z9ycG/ONOMYfTeim7gBVzSBkbO+7e9wJ9fjyn/gEjFTdL
H0EKRXQZo1ITaGXIzolkmOOve6He0DaIHu3neALR0yx1eFV7mGo1ebR2EaQmKNex
06+L7kMUQnwb31QHwUjvcHwfDHm4C9cKPYf++VaUHq8RDShS3pBICb/skmVXnOUK
enzyMwIZNUa9vZvKxG73IbESBOpcUNz4eOebxSunPB+pmwY7cROMogfInv3YQxfH
ZnDHjKKlSoocpx6G/G50vkr1T3vBd8fOwIDiPayrvhd79GCmNr5ixQ5llXE/nMAD
2lCbCUIbpKlwbCOg+hCwdYzAdomUQRFUZPtBu91m1JemekPpddG3rhl25SC1xj0g
ud/zP4Ri2KhLDFnPzHaJSj+5JSljBCTxtqcC/r8iuqgA7W9mWtp1h/QelmOdrFQo
YIZtH8nD5wPc7mLn4UiIMSUK27IwmxsraV3Dtd8+xUXjpId6H/lUc5P9pjZ3d/If
JmJ6Tm/v+nURnnl2+JoEjKG1SVYqKNIQjx4sUzm5GFquIRlwoC0WDwgSeResFdDh
13dpXQ1lh55c4IuwbuFPoLOkmGbduxpa7yRrP6MuRkduXCIR1gXoygDvCR1KAKiF
0mJKz88v4s87bZ5ggW0K3VnfZn1qujeXXkzCHmrcGtr/yubFYS1fV88iT9W5K3i0
JnkJ9z8w0F8Xz3E2zbxoQqLBcDz8JORAtmALAEaHPkwxKJqvbRcRyAFRE03IJ5N6
JtqI1hgPqpzpzsLZfvowXBZUKQ2y8czxZruH74vC5KEhd+e8HB9Yk70PA40xFoa5
tFeCnRgHypyyMj6OsuK9frsMVGBNOYhJbHU0kQm1hYI30lzwya6uljIno4ltp3ed
C+2M4hv75II30IVML/4kdzAnTxvm7KhNJPMcNQj3S84o7OXDWl1PCsjTdU79Mmf2
YNhcnPo3ywrITbWH7Bfhwe58H5wz3B4d8t23Zr96ZNZjoNNm89kD3AvmKLM07+2F
1J4dzWDTaX9lNFYw1spMbJAmGJWWH/z8h0Zmiui37hbw2WeRHB8z/D9CpcSBnn9B
bLCzfFLvumpuH68PJ1naCxODn0DpezYt9qNZx9roQZfuZpnb7O+ts1smtQlaKMv6
MEUHnndAQQxDtnZ433th/TmENuJynmLWt0l9Wxm9auvOeLhElvZB3HMUbXsLCjRy
2J5Om2jWZxnUrO5T6MZUdo/KITDyUgHIpHq41zY9aYhfy1kmRNF74dF3Ad7NvJcM
loUT6107Qzi691I/2o6LYBlEoVL/Rl+h/LLGL0BKRLzu+KxB6m/qQCOKKxOSR5n/
Pv822yXHkWrlUHic+jiao27rNpKc6ZOkJUnIpmbJZMPg44npszxycnDdZpZGatIT
faZLhLQBvk4/VLny52vblBRmMbbDYfxDji2frlvOhPjqdSV5XF1+XYAWzHYzEA8f
V3DUJ3MI0qpIi55Nfw2yr53HGJMaVc0OSgDGrNWidYt2hSplm71lHDd5pcxSg5sJ
0lENCs387ocDwdRemjfWP6xyedebWLn+9ErMriEIaAYFtkS9Sg8mwCUSsK7uNayL
Wvb8pYjjXzQpHlNxJCgq99KQlCrPQnaj4iufC7x96v8mPt95wHi1I8qDp1bNMmE5
+XMhUZcb2ZZm8phqA9qVv0qY2cvs4z2tw8paAKZG3t/iPxPiqT72DhF2rHj+K2fv
4A63EhNAb558Eb/XYBc3XZFCu4IeF8FtjvPBwHI3Ko0r4fmZ16GNgwN7nq4gTi3+
8bGUj3G3cgF73PIvek5uxMXzBKRUeegpTxOdPDWbNjtYrLGHOZpqZwcfoPs5ikHv
DaKrz5eL+e71hLPYaN/k3RwIqogJnYYhZJVob/x3xKhvGRnO7chNi9khGw61Nnc+
tIlVS7Dy8J5vSEU4hSV8v/w3uwCLu/7z2u2Nu3+pvQpvOLnR2GfwASOOkSZIEVh4
B2rHMNhf1rYiWreU34vUrWXa4R5mEhtOEBnufp8QUdYmWdWjY+zpexc4EWlNnFLf
qjAsL4sLRhnsH2Ip1GxmuiK0+CrYd0xy9bIEaEpNJsJ98UWjonzk/mpY8FZvK6Ou
qjzhitYgOcTTfFJhOXn/LNMcQIOJ5LFBL+gqOcr4Gj2wkuwKqBWsIw7IKej2ZExM
Nm62y9QJydodG3v7luZh/isWxOZqaxYVH951f4/+SVGfPL+094DQqyEngnyBwOjT
pZEwZlHDQwqi2vgxommEOFld7zjiiCDywApgRrP+5Y2Mj9eZE7AutRezHgj6kzVr
WF6Z3Yh7BJa4TKCyolUDdTxy8cI1U4ytZEmDztKx9X1YkgfMiDLOAtpWkDA+ZOCR
SMMihk3Bqxx610eebvdAi/LhP2FQN7vZBAPt7DSBus1oGlWJrfhALQ5KFPNZ1MoF
qTPB8P88wR+nxbqtlKupFVhWQiWA4zqtjitS/+6wH1dFdy9+aRb3ZbijADO85M51
1heDMNkXqkHowmJ7RqAYMoemgOdHsHzRqx9kldn4O0jdhDdnRU7eD9iG1iN586wj
xbKkWf1rpbhdyaG23HIpouv9fpH3VSgVNVuEC+7JHWXuLbWRa7M2A3SIw6vkD4Lg
vTcfVj4WNRIsvyHmFcH3KqXwvaxjG45nEchfYzglKzuJTbUs5YSN27UDPYFRgDXn
ZssO/2NZoGyqBbKi4T8ymUIDtH6873EdO1NhRTfhVN2KCS4Tc9DyOTzU7/ZHxL4G
iOD+2fbCV0j2x7CXG4gwOMv7k3KYl+71eUTwNxwODSB3jv6D8laVJt1TPylD/b/V
53wYuj4zie8NJpZUwSKy2KSXsBo/zgMAYlk7YNrebEnunMK1P8YlHyCa3x6AVzrU
OMw7TChYXNtw0XlmkiyadpADIQ0zSkI/SVUUDmH0tUFa6KRStIqgKZ217C3KbFoL
NAQiuhL7sj4peo8h9uJhGayqooDXXIrd0f9lM+NuJftkq++SmonFscCjPNF3uT3r
R7oXvH+BbZ2T/6QROMN43EEf6pAKwA99lT5X9j9PSqfV3J35U/cwLrKncDlgZXbt
qg1Gj5qPU0LcRhO58yJBrfcnW3tuhtoIcwwOUv6YCCAsnFH94ZQkrdeohHpL15Hd
k/fwWAoITrDR01PyXxDczSIQO1fX+XFCLCOTbN0R2jQxrWp2QYBcBLv7c8UIOZCS
Fso4qfnq/XyW7iofDHNCc+rK0onSby0xMu/Prx/XZ4x1Bja3UWB6zF0i/77Egc51
oa+14cxdNAhYbL01iluRox1MxSQKZnKj9C1UfSnKKknmnxAqRVCqGwSge/tfAH0U
ljo8WIABuTyDTZsoBbhkZt7GQb5jufk3rCRNnGrkXWuGjwJCguxd2eDHOhA0AFzi
wNQCh1CSoZOU1XoOYqZliyjlJolK0z8ajfZ8xNlLYO1sMX5fHC5QrKeMzoUjL5Sh
JRfepQSs0heggPPCYjBP8wMmK5XJ6pIceOjhN7GvVjiddFopOr18/A8J0pVs+GCz
PogaTdeiJ+jLmR98w2pbcUgV6e8lcUz05Ek1PQznYwvZMbDaMZwKFoVwZjNsZQYo
D2BeZwFIL1WA9in0fQm+1GD2YnC+TbN5en0C0EUH5iamVkfSlFtL0aVz1BU+8kCj
QyyQN/dSYkFogN/JCUh3+kHdGSsY35ixGcLCaMzFC/GRwNuc6o4Xy7xXzOLjohrT
IoOxpR68PP30PgWN9ogrHDDozdchrCqTuRi6C2XQPSMFoiahE1yrn+BjZkhGtxZz
Ifb+FGQ90f9XtLt/rW6EgRvCNQzPjiFfL+aPuzgj4iSY60vNcPRyNds7Od49GuDU
2VhiK90bLZFDtH0iZp7ty4xDmdQJv+blc7Yd2bCFDGZ9AdH1Rer/E53OIaxznE/2
mZ1RvogPlcYk5BuD/yVTYk56k+nm2EnprKQCxGlggZN/wACmPLhfCuXzYtNdVIcr
33PlQxIHERzSLVv+MpXaTS/vr09bIiR0CGxN7R4vKn/epv9TSqzXT/xn/w2oeBGt
K9+n2+KVX13mOC8e75xkb2e8xHDfKWzqU6njp9vfUSiC5vsr7T3kLcaB/5Hx9c0i
IyXSANvdejoMDZ0jRUjVzZ5glAUhSyOVWUcq3iRpZr23I4M2tRea7b9pxfrAQKKR
4ZwZTNPN56WX87U9M7VczOwkNf0AfoP5uoj+2ZPrEQvbPwfGFWZh6MQ3IRU/a9EE
UnA8J3MKtv6iWWwwsTYj2MHfIobUi3S1IEGzKMAx2qV5T/beMohK85yUKfbSKyqF
7z04bGzq+50h21t7o2vrsVwb9lmzoLN0Fq3JcbBbJpkWyWvEIj2l0l47i45lyf1i
+NLN5M0q2MIhWP3E/h/+x6Zrp/E+M3TozyVYskBKz6r8ubWb+CCy1BmjZAGFMcpi
kT9mDBBQc7YYvrJzto5R4zM0ea/DhjVg/fcl2Sf/EN/7myAbO2PnunzPfq0rk0jX
HEMFswjVYDoRsIg+NsVDorLWmbQSTFBhxRtpSwHN9gA7J/gxXVlFz4/IOFwootsI
/d5wPtZ5KaxSsuXH2eSPlE7ivmAQRhvLdbo3uGmtsCjrCp3qFB4SKDwazaZcNbMQ
GUyEU6sxrq6thsZq2W83ux4TvWoB1HV3joGz0TwCBoVHPx8hrqbS5wTaN6rDyPjK
1yg1o3JOFRJq7ZpaifwsyKGN44aLYwcfLBo0WR8rq1Se3YQO0tkxjdm0h/6UVJ04
Jv7OmArggPLEBSt242/So1xmhND1OTUjf8kla97baZmIwsupkzElEl9YQW/y6Rkt
BMYJ0ojvYHrVdBn8HcHOF7HeWa16fR+4hGC8Pwrv2djpd1LkKcYb8XQtVxnKg7QV
wlGesYa/0vXtIEq0okVnA0AGRTFpSpnrmrjq0JlnESNm3RSdlwSXPU0a/f+eJ05m
Fo+2nG+aFq4xUz/6oGGywdbgmT6dQDzIJ9peZIWzqaVpKe03xUTCthpbmuk7BDkU
85vxPssnW+fNxKZ3S3SzMa01CRTZZk9JHq7o/Tqa5+6OeHGUiZx3dFgD71Q1lOtr
asnBgBWctdlt2PPVZib95GWEwMusO+hi7sBnXrOm1z8JoKDleQYb7S0NlVc1N4pt
VxURD7VlKsRfm5t7NumvSJvhaimHK0VHQlUNDTVoqVTBKLVbd30tw5YJI5CL/ByS
EnVnOIWG2a+My1wshyk/jNWnYF3ATtu6IqDCDrxD8bqsu8OK6paogQ1u2w6BSBkn
DA9uuJnWhvSb7lpwJ3UXREU0NxXfuhmGJDeAvBmYb/zFLG3XcCs3D26fxbigClyd
6VdySY9byv2C2e3stWOxM/g/KsmcGsVaa01dn67gPZwPvYDFJgN81tzQK3fQ6nJp
baMLokiPzu1QgF5rnqlSIbHE9ywyDRiXIfQMMVx+Q9D1jXR8RjEKICPJPqc/XKBm
3sM6PE6Fxr/K1WmZOeiauws2JNOodAS77acEA55J0pjuWyXA/RO9W+Yzu30szSpN
iLhXm8wnC1QrWqDgQoKYEvdeHyDxme+1TtKU2Etl2nFTNV+5/+YU+yo7Oq9FQUoq
G5xRBO3q3M141RKdvYnIOuDjjUAMkrWll1hxVJBr9qNNGCqM3hqzDCeLWpvGrwvG
oXYPo5cfhDpxjvpek1HQPTO+rnapyvH1LDuCAKAxzM0VaqGOkX60tbTSoWlW5KWg
d/g0295vNjlRH+zCq0pazBE6NKZ+5Z1TNN0cgX6fAald2LA5ffsDx0Wf/UKVCX3p
+UEkGI8+fQHpfmw+nf0FTuJd955nV2E9+aql0A6TOP0bxv3aAjph9LDAAm3qN9f5
wN7REV6N308hJo7a+8ChS8Oq0YmciEoa0FPMQ7r6Rf0/hiT0gqdQRdybHLTttzjH
qs7RCw2wJgdtbQYnz+HTuZev6dtddbaGEZy1WLLpYdNtXh6nafLHd7teYo0e+dh7
lr7ErW0b8MIIqje8L7Mu1CDtbxaU0W4cP73CWvgxo2hho1MtHpynEOZ0+ytfCexj
qzEfsxajb/ifCg8QL1HrGofHQi+D/b2hLVLOpWP+IX+xZnA3UGecmhcaZAjZxUjs
3ybew29hitexQusybxjr3YtQelbITlhnfWCvY3hmZKx4lhx7yHKF668zWGroIIVv
9DEwX1QGHAmLwaOnyuo7HC4g/z8nA2o8zBY6aSGrcBE8dHJF5UsIWvNWY3Mg9Noe
+Su722Dup84fPl2k8UFoz5/BnUq3sIoTyY11H3nm5S984vyZ6QEH8iaaKdT5Dfgn
H3fpMxH2kW9QL6GJJwewHL+XRcfRUJW+7ijPcLIGTY+wOiCIgxFECOmPd5xHi3d/
Z0EMepz8Tj0ybCd+L/IQOCGrYSs0S8jImV3z/x4r5n1SCEp0uFYzWhXHg+ZKkeaR
3LVAkFHd2jhXAbuYMITzZaRpETeZmkOZ708Y+Mp9F/k0BJHFXkwGl5iXv7y/k8Fc
DV8xwNxqNhisD/XgdX0D91NTIgzZlxpiSIkvmQHSqiM30Ze8y4w//w0OpFOQ8nn1
sXoflXjh7QcgLaHSK5ZIFeWTy6ss4uGbJ4TXFyNqstjTe7gtgCMB1wdg1DsFaRkd
dtBY4DA59mDJoU89kj9TulrQWd4070+Pd9XgwU/x4q70/bu7M6mejCE61oFjpWax
6MT1L4K0ABqNjrkExnBfAr2F8ntb+1o+dM+RRPk7qihOP6v92SPW5xvfvUy2xGK9
rOuwDRIaaCsdJ4rxCp6OdavD6om6TqSFv4fnbIlVXNgS/znBjwejSZQMip6Ae6Nq
PX8YKkpFEJ7BrD3AnSZF8P+BPTqTLzJdVeSrUdGpr5jEfgTaDWHRHaRzrXVo7p/Z
KdWngVcvJtCH3/xfVIkEh74Mk+0qkTkzpf/6tIfzGNcpPObdLbktqnO+1q9lrpKf
4mxkLk5JwsFbHE09AZQqLjBBwnIg6R+9NsB/OUiRGjtda1coXTrIaKdMEYHsCHEe
7dgRZ4KXRcfVtQgGwzyLkXI4uWYuIwfRPG0gzB8ZeU98cqm0jiTkF91w+aIIuxmu
b0UbOZF6ypg12lXm/ZkWP+xLVvXBozahP176gypTPjPEgi+632qJwzW7yRhVnqoi
Iyy/Dav+gL85Z90U+u2LPkJMxQxibXu3HvjfiKDBsp4RrqM6Erp871BezmP4TVeG
Ujt63m48vkO+LN8nx3/vMR66lcEPpv7B6JK6a3Jal9ZfHdjmu7m/FSq5F0r6NhUg
h9KcPOhOA/z8PQgD1JfDOFs0Yqa0NPip9GdOcwm7gmGy4SI/HrU3yndVRMlOPnXQ
erVlNq2S0VRkko5sv0GXrhgCbseXCPke1iXTJ66QxbGHqLjlsTz0anFzOeYcs/Ep
haBLXo3l14cwSP8aujyMNebObfeIPKOy/WdUqsRWIfYwjq7GKCrW/e6mAaLPGItN
mBYSQ1qvY9LhFUnw2A/nuewDUxcI+hhRgdcWBYnE484czBEn4XVobW7vx67evCcw
2pWcPfoI6FF9johNx1+km+jCkgb6vscXVhnT+HrQtPkdt/9N77IzDGuNVgSl7aae
65xQ4KrTS1CK/JnCDDu2bn/pKXzvTTgrG0gtFHSgq5UCC6rfVnxgmaNW09JJgLJo
dZ737qDsa0boEzTegObtx77bTDn/dTluTi1xuXCArNwOi8Tk3++uyMO1EjDOHoZd
ADNjfQDFLxaw+CXXMrylgrLy3cwtjAvRdzS3qEnsHPw3AKv9eCJvzGaJr3CFT4tk
8nF4/4sxxBILxTgYEhIA4eibA5pA39QyiMU4pGQV+QFCixo7Dr0JEQQEegCdU1Jq
OqAUdZp8FxxM/C8Cjt2At2xOUikZXf7LUEyffyVWNGivBqKJIL+QHQq4EzpCUHsK
HTmyFVKeJEhR2fKfDLi9nB6uxZCPr6onyPYXlF2ys0fz1q5+Yt7lPUss79U9DgIA
ibAjBybiFFLQo0Omt3nOi44FroeClbK8FsJpeaAIsoRZMuUXv5ZzYphCy8Qs++nD
xfU07c+fvRvXDuMEoClb1tO3vMZuX5SMwg5dsN5LzSuVahIg4Z48TAlqd2Ufxm31
M6hCi/cTfp8xSl5eNZpVKVFsUDS7D2uZete9Fl95ujYFhDlQ5svT4muiN6+cEYGI
+ZVdjKbnlASL7zGtsich92H5/pCOZBKO6sYkGO1CFQMDH/eBZFUyckYblCRsPII7
NjysrKAnf07EwcLi+08h3DGRII2yPmXR3M8RetvWGkELA2FjCMydbui/jNMfcDW7
5tCflhrBF0SM75zK+5yJVLSQWG5nCK6duEhOlWVr9BVTsLYnQBaAjbZlOXFaKWys
Y2c7AclzqhI/GIcG9Z8/a5ldidBZeU6+w9Haif3Cg1nhFPiFQmzTioPwoo8zd4Ks
MieufWLNDkn3FVWOtMku7TWYk0UIlVj/vbDxp2JGG8z0RNqJDPq4syA43yTMAo8R
AV9z+E6cSiBCoSWj3bl6sofmZNMUEj2waOgucpOwnIgI3FerASZ9d/yHB7Iniv/h
buVPUebizkw5w9Dgo5Cx4PkVT5Jn3xdMYgmpcNOSHmLRbv0fPkTXY1k1MjFVUUKF
s/zGCsSWBXX3+s2Dwe7/00mNCNN7UwvSbCAXnVd1/UkJQT95rbyAnlGMuuTKHNQb
Tuta2ZKAdETa1bC06tO7Z82/WgElq80F77b6qmNllmdGw+NaubYjMP7tjnde+B85
EU1LtUPCqdm7T1vAW/n45+uDpM2GPqwShxK1VSz8jt9JJkSy4LEwLUXEkplUVmpu
DNqPEdPEJ0xR8kHLoIwTcjG9RsSJOCqqaYS9Btyc96RKuNK+oKWedSbjYKBIYgUr
CZ/ZWrMsqKptXqDxwT+45+XknfrKSD6dZChOgn0emH1jJ+4Dr5Rv0PI4xdxYpZ0O
qQ5KreDenNdcyDG3S2Q7zDRsHAGqqO3azgApbzNnZ9QOLRJCLcSmdSDcfRlTtl5Q
u2Xcwhszxh5pMweaVXfoSynAADwj4K0hUGBeh++xuAWx9Yv9N8ySVhyX/Al/ve1k
K7Z7nsCrsorJ40Iqfxlw5x+LxJHZ1rNiVCrb2urDmk/C2TO7LRXNWEa9MKv1EwfK
ofAL5VIpdoCBuFUcPMrNAFXzk3WEcd1D0v0tXIr5gHm0RZJq0ggVV3ySl+cT4NeT
Jly5p2d34RTrW+irU6Jp02SO9mWWWI/CAZWf/2ROe/WDjzuRCQY0gdALnNS2Dxh8
kgBAo3GS7DDUjLV5hT08kI4YMhsytS5NBaJMWkcWOnC5cIFa/Y0M/z+PTJthe5rL
42A/HHOCptlvb4bNqOnbT+yQAglRmQA5iBTPxgJvS9go4EdOlnYkjSTp+B32ewzk
1Z1dO5Bvqm+bJtwYULLAUn/prV+UOLDhLA1kfADQjaM0j/Oudc4+yZwPcUQ4ifE+
aHvzUcLd4YALVGKQ838heE5g062aPcioVqIXH0K4Fn1ulWMn8XaOYgLdvv7UR59K
5y48RpyuXs5t2H5hV8/U4r9gaT3FmFRWEn8WRjD4XA0KQYfzlYCmSgOrxjGJn7Rb
iBjbhuB8XoTPesDbc0lKtZr0vNsVCDsydCAoPxVYHjauwn8SRjckW3qPhUTMPz/A
U0QGqM2YwV3mfs6ziUpOTFuMvmNKeqj9klq/FaOHG5l1kt+SeM2hTEN5KCuFmtGn
/OkDMj5KXRcjsi2c40CCkLvAvaJgvJOUZSUzHis0GgQ7axI1FBhSwL3dk5f/cT2d
xDRsGNy0tLIwV6cHkNu4CQ7mqEnvxYYxxHTXJ0kmAwitjCdrPY1dTZGx6+zVZLJg
GHnJzPS/KzSfZfaf6IGOeNYerzwK3bH9o548tv/cp14HZDkAm+NlB2VJ7+cgupEW
e34sD5M+yQbHgRwIEgimVnPxq5oyk2zTX13xPD2LGvLxEf4mXLsZbaVdY9LLVIL0
vjc8FHhIWHOQYTq6UT8C+aF3nUVbyOv98HyFOuOinAeoTS7iUE+BFZbSxzhuyKbD
ovPF3OrFj20umCIwGntiy5a3ZLXpFo+QQG90+xN9a4MVMpUa7Dri6r0lcQbXisRP
tAGTXWjH71E0Jsi0j7IORxvZFEKKMcVWSnfuL6el5uXf57RcxnAMJvQ/iFomnl/I
zru/Q6kkeO5gxWDUngTbfYpQi23+Rz3vh/uAbzMdCXitbC11bZxn227Sh/ZYSL1d
G/cp5f5QeEJQnMT4hMTzWAuozXAMMZ6S+Iq9vz03xfE1xmh5BgW3dQSXbPw5TFIl
u/qkzVVJHMwoWBFOWmqmBu51cbTxDSkIwUcV3BslPQFVofoocrugDajVSGht2eZQ
/MTrOMnbU+oH+IVXo9TQiCnvqwwhFwsBE/yIt3bWJq9ZghzUGivqf1pu5Tq4BFym
qinikDerySr8rZrvIxL5xeLFSN3UTPb+tQb0TeGCj2qJsFuN0ZddojN/Dz2GHYD0
jNsU0nrlnb/VyHZkAsevXSFX9Zwp8RemXpPvEfLyPlV27k0Cl8mdrVDvSMLJxEyE
ILIGke+p5QRhDrqPOEY69m6oq3ydeWDYkdkVIIHMfrPDZBPa1ArEYWveCwu2v1cZ
OKLWAZ12HiIBEco+ExK3EYCZP7s6thoGzsRmXpsWuraX4dZyHmmmcDHm+7FZMWyG
zjgvS2jdm/R2VHuiiBrHqYJ0iIlCJ0U5vPuIYmdYXR3JEzf3TYKoCYLhQu1hq2D/
6SxYQP1x8VGHQFzvhjD3cPgmBQxMhjXYieGy+iR0/sgrzMRaEgUAudEURHb/mO+Y
6GR7A55RwH55TEyty8aXjQpEVss1J4/X98lfIMWcKMG38/FTJefAQUZ4UbImtsZO
ylc/uNqA6LeMer1TwJqBIbNtDnerXcYmHlgwrV9ALqccYdcHjTCwIH8xMc2WQy/P
fe605QN4lvZZ6o7FOmROth5SSmAk/GyP6MMWWh1jWJWQMGVa/FoC/RN/d5s9uEmY
7PAfHc9iKauCdNBe9JPu5M7lBI1sF0Y83RXcin+160zS4jgK8k9sfHSaZMVGP/Hd
YaMxY318OYBTqO1DjW1e8PQCaNgEvl7xpBKEyy7uVoAZnCIauQbuptfeSZGOm/1k
0+g5aqLCLiYEUEbalw91Z7nxRqm7J9H5Fk+dL86XRZTMVAUH9mHoJmECSE6w3id1
Id1xH8lvm2P6dXOfiX+PmVh32YNEYVXZTpaeht/OdIJsR9u8QpqfgCsnafrWwsrV
p5rdAtmdy1KWVr9yTtUwqG2Okkl11Nati78D3jePDFypogfGKEmAovtyE+/RPE51
2B0U4y4MM9IPUzOBdW+2YX4CadB3+XlEPdjqOt0NQwjFQXRoq3gGlupq8j3vEprk
F4Pv+gXRbEGR38BMAuIt1hiu8y0fDgnusyBnGZ8Wwnk6+AFty77dfw1EkzCQEZdL
mhxRZXDQ+Xg0Mqb7aHRk0Lxt3YdIaS4xP0A6cs0lKIDF06g44Qyq6Uv2H2/Jo7oz
FDSZ4DyHSECdwXQPIqOb2DbGIqEjYNwyioke4XaFoVWNHpYBdZWQMTgZ2KhVen+7
j74ryOZDC9HGaYl2so3uISX2Fjx2TMVB9o4tMZsQPNY3S07KX2RNx/k3F2Yi6k+o
TW0tNJSg7Z5KAUXoRW5ucr3E27yuwsfcwTCRPNkIkqns+JtxtpniXSIGtdwp2TW1
MIvUGD2ksaZFJxufXz5Nq0DIpDp94NDR0X7rECjjIl1MNBO8058/hSL5E1ofu0EI
A65s7HK6P6vMqkcsVrSYrXwXt8y4JFa+RNNYyQH+pptEMHnI9pY+GyhEzYtZgtYs
iMnARSdOOYJLk3r2G90gz6QZR3lmB9bYpFjrHR/uf10zHvWFX14abauNGMKc5JX2
O43oZrtMpkeHYNyYlMxzg3j0Asohv1eSYx3z6WT1gaIHrzEGgMLAvYAAFb0ptx9j
+fc+f3kvz+EFhzBbsQIYvXx56J5hNCdBTUBDqodElOn02wN8NDZL8cjLBThEk3V/
gHOF5KezbxWuvHeFaPnUqxafLEMZ/iVPG9tkKmCVh9P13X6WaC9zd+RngzpFvfi/
MjMeltC9ABZRFeq6h5kuPRq7OA4Tz/VVPyUrWhn8cM6iFwNOi8Dy+p9czRUPCel9
Xg3RBZO6d4ckCexJSayDju6LTw0A5WAQkVQ+HoxPR3GmThbss/u69L+DML4xX1IP
8dkXwyT7efaqPZ5YdVYcQ4Hx8t3NQq3APJP3RZxd//RifuV1wbb6VlTNzXd68xzs
Dz8KfCbW+LCHOHOh9eNLI0tBxHbGVYA12OfTR/4Pmkyj2MV3xMqmKGPHznw61+BR
ZHG7Pzb7UetgOpDaBX9O85RYwU0PaqbJqaAQ7fenVO/5S+ZaKDIzFY9cFHjbmm3v
4/O1+rHys5QSW7rebcN8SmmAuSpiwHkxtB1XayEf5jgRj+Lyu3eQ9DvghFQ0l8cd
y+TdIMwRadwrNIrOSwM2ldHKycX3vQ1owk6agUKS6LRDJ9rY0l02vyM56Ab8JzUy
ek37hkrqF8znSnd97lp0brP6lL6wcuRN2K9BfRVoq5GqWt0kfSMsExTf34Wp+/6h
JqU3NBMFArJLiUpxyiso2Myy0fFEUm4wxz1jpSkXzS9c0rVgx2lcXY/AE7o/VtDB
GltAhkrbRilSr42DykqdUUvhBekpDxZiwHIH+rJjs6z0jQtkvnXGt46fnofIqbFu
jnIWU+/nqOFhEqnWFgdgibN9YueLgbIzp0kq+ESiqqUUiU0ocEGTtcpEaEWpL7QJ
7qDbjHV8cmSUR9KSekcCNAPFpBHzVmWD7X2lpFsLVij74Y8v21JDbfi/n+bEkwOe
aWlJUUOkkKCk41Ecnk1K8CSbRlVFyaI96OpWH/ZoJQYCFYFqzQl5/KFyY3C8irUO
KW1M9yvULtcbhyvOly8xHw8l19eeUPvxYODhj7boBg/PMwPsJ2ZCM3EKXYyv4upW
y+8JFkrzse3GBE1/eXdBMTIWFjTHTpqL5LNaXIShp9PDUBxMyEuY3n6QaF2vc2Ny
rMZswCFAyNLY4Qe314TJLdUO1XP3vDk+8AqjOfC5Lb0=
`protect end_protected