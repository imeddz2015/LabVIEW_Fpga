`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 3792 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/9huKRhRMtvnNqb3Z+UU7TahEoHV+T8U3P3ufru7l1O
3DlgtZzb9QxCbOjthp9+wDkjygH0eUfDrEl1ovhZG60I98lfhEZH3JbnarXOIuXw
vdfQQq18+wILjpw4Ebi1+AHfO+CjmV9Zf2UEGAJp/8NCu7j2y45yhIib3/RTznKR
Xe8FbAjxZnJr70l8n3AHq1AANeS+mE0sQdEYMx60n53mx/oFbw8ONQkRItKAG4GL
P7RCR92SzWM6Ca4C3f/AjZgnl4+SyEXv1+QtCz+Z45APhg1/TRtHVZofvjwZXWd6
Ml66dBHba+UegVMqBI3KLVip1F7Yns3XzNrzVcU42A1EJdh5tOufxYXVF7kIEsPz
xJ6G8gk1uoNUyhI4Fh6Jfs2ND2TkDSPoKqyNjiCPemqbtpDw33vG75bu5JVehPLw
pBNh7IOOEKFfMHqdHSVlVx1c5nVvVUwAly0xt8LjJHx/dLRxVUzUwsNeRLUG1U0h
9Yl/1SzsBkVcZXi5vmzvk0dFBAMlxwCPK9vNfW7b5TiP8YlJsSLLwYgABPPUDor+
PT/FAJWBPbJIdMIe6t7y8k3nDOmrQqjc0VEN9F9GOoM3dpWc2tRnxPt/H9oHXrsn
/mSIDyrokMrFkasV1lxgRE0qrvml5UZGQwHsZakcl8PZ/5Vldq79AQ6tdgENir1j
ESLz/pJojEpHyYS5WhEh1UGZjB3R3QpQX4za/A1xiyq+B6zNN7Q4uFCRUxuZ6HsR
6Mr24/I1iWzFGTJMUjAGD8BirhmYQCsbLesyDD2v7zaSU+wp0RFYvjprtntMbtq3
kJ6VuvNqqpoKCbSz1kHfaH1Q5e/sAbs6Tzu4Mo4fsbFXKsd6x8ielhbTqPCtJvwT
pqkIyXHvYe0Qm3r5oTReVFOE597+BkPvtMMXrSIwx/H+Us5KWU3yp7p/bGALzySu
CzQWRDdyT0IJkQT9RbzGFaR+Ca7RekPvptlOSz/BSPeBq8pSO5B+5tVtfecdU/t0
Ftw5E99zld5hAP6ldJ/M3uWqhQYQwmbI5XkOqSoGjde5/bqf+JTzW8uybi/8Ubto
ilj7gE7ktXh3bPwDSzhXnqRqh/QaL1lu1eD6raJzLqR1lPcWTWoLofarnPhlia5Q
XfHwqo49VTjABdYulE2FKZdpSkVqhTd240DuqceVYo3qjspkQziuYNNbdtdFA/B3
Nplg0S2ISBExnch7LBUar8zuJr4LfjSXVcHCidXoPDyGXcJUg6djO3+w4/4C/1X5
CVKouQ2GkLO3adagh3xbYxTyFr8W0FE08tKiM1Hk8nGvsOb9EaBkBbxXuZkeKn23
TCz1M+njnszm5FbqJK+KJhghNJAJhT4WJVGcM/zJrCTUgC3M9+6HwUkFbGq0mUKq
7+TRKQZBxd4jUrYW6Us1qIGr9T1zeIdWLGYll2euInJMzOjaPjnaJ9LMfAxckRRg
ZnZNgNrQ69uJIbzMXSx6yqOwzz11LJsB8PkncPQwrS4PM6sI94LOL3vrARvJl6NM
HHR0cg1jmsBEseI0fZKdMzcDeZktK9SgH73jqe+/zUrAdBACQDSL2oYPEIyXEuzS
ct1D8gH6PUfDQ39fPKB96BouGcbHHztSk4uN7zLLTrdD0fzF8aVlBIt/cyHC0ske
oaUXCe65WGNW3iTKS/xhGfrmD4aMCOnUYcAefByMsa0Qou4x1h9qsv3UOYgNxoUL
+j/MeK2su+UpykH3vCNkw5N9kexIzzi9DNCVZBaMscvUBSG1JmD+02LVSK6/oLL1
sBfbuXah5xuQMLM9SZ1VjXpekD2JyVxCGFcXRczmUGNel3gO6DeCoo7JGEZmyknj
6iVCMhrQMM/3Tt2X/OCjuWYiBdH1JcLL8jEmkA2/r24vU1ThvbrRyuubOGmwOclH
/Jo+g2qe7+uHnr2Xy2MXOWKQcf6ObPo4GadxPXAWAo7xci4KYZ12PsWUQYxCudgM
65ujH/kVchvzUt1r2PuPqfYTELoC3y1+r4OsoE1IqnjYw6QSH0AY/SeK1BZYIQW/
7/qPoypoCNLRxswdJbDx99TbJsmZnRHzArD02VCVV13kcS6hxbcwDjVCSWQVsTnK
zInRV8PT8CY2P109FtKMt0uwQqt+8qeUfUaETqQuYqaZLy23s6vrvSgTWMX90dMG
LsA7nSnc6eWjmUKzl0MSuJAH7SDbobJrTUXhnnRRzPJ7PO3ciiiYpFhbRClzy/UB
L6jlTuDyVIf4Pyo3zV6NYJCU+pZirG/gNstj5Lq2LLNQLgEiLsclaLGY/Ot/H/Zg
8MysHog12Q7sjPYo8na5vNTKRmpMJcJG/xlvtAUdsJUECzWFt89qnYdqRUT5RdXs
5tj14KZIthyT8UpHP9fPlstXzjVgIx7INv5lNuHw3rQrbqZ2/6WwJzZyLSFX4Mmj
vX54KwAZzOWKBPwLhmPqPwoKLeBU2V90s5DqazLkPpc26Puqqs2i/t9sNqa7lSYV
Chu+OtXnkOKmg5NxGoZlO/lCKVWxCkqWlFzL1/k5C2Gilqgag2Cs/kU+wVQOtQdH
UqQgxG4wFAJLZdspVkvMB9J/1CJD0qiPynkLLFEcU0uv+KlyCRLI5R3DrOSoHKG3
hBDn1nD++Mwg+GzqY2Qn3lYDAe2UO9bSUIf9xp/lBUF/QLMTk0sh2PbEcbeuCUNX
XDtql7ah6iUVyJPCrRhLTXS2yGtPwaLhbSjvX+aL7IhalVH08PE1HOaiSrwHbt54
ZGiUrIDHbkdCHIiCtkhLXW4m51UOFgCQx1fTNJJO7dGY6V5bvq4y4woiglSgVOoD
5+kqCwnsNBreUDWAwzTbJrHklSyCxmE9PCG1Drja1cK6tmy01EWhnnaLhuFwnk13
q7+holpyWEWmTYeKuoE8hEYpuojBJEXQSUEKPWzY6hvbzOYNw3J7HtLkoL01+tOY
Pl4OJ8+SCuNCAS9fZr2we8qzM+yjOEyotJnI3dVvkae/MsIZ8TgyR0/nxf505SVE
cj9O1HPEluKu4ou3z3j/7HYRSVWQLd8wXzJ+ypM6mQgmkPG4swSGtJ0IOcXrq8h9
QququeZZGlB8sPgCUMqmedmY/wziCd9zz1k53m8IpxtQBzWCFb45c+j2mb7yYYcB
oVXKy0rXiwjaXNCuhsjgG23XkUO2j2ic2bsYJV10ZKJZaVlwcktdc15DnPHoshPO
rjHL3FbtBWD+reRglmcS7sxtqw7PDASGPsuIsPPC3T1F3cCmzAT6vmCRF2aYJIsN
hECKB76TR+2k/VKV+xdTo+39takchfCdBfMjheM9LvZbL3pWonZq+CQx3H5k9AHM
i3hgoCsxnHTioWu4HI9yn0IG9zta3YSzuJ2y7Ex9/L+dtubYL3OpjcIkT2LpUzRl
TmPNNlDcfz0O2ZSqh+Ce0OAuXwRy5qSkgXetCny/tIA7r/lKCvkDuamfztoTx7jC
FweLv7R3xMbFE/eCjDoYj5J508q7l0oNQG5mpcFfw9otTOhqMGdjlNLFooS4UqSo
49tLFTKMUNgZ546yY32uLYg1qZjcTXHFxrWaKw0k3Q+iHPK6dN4hVqQawvCAgL1+
OLy25arcqZLtmtNFtnjt0tLrrVPiIQI2FpT65yNaV9YWLGkXe7FYRXrhJUKDByrA
1hr/GBDRO7xQLofnxMmTzAaLf0srUZFGSzDVfX/T5XJ1HVb4xcjIL3cLv6L6UtXD
hFD3U45e1O/f4ofRB/Eh2F2lPWEn9xDa9puJXgpSXl3n1gU2vy32hFWoRBo2p7g1
/YOXcKfc/ZAla2BjeFdOcSvtnmET3xT5g24xUIhdQOnXLID+arqD6XrLcm0WHKlH
t/nUewG7ZyYlKMV4VWY5uudmH8Q7NiPEf7O3QFt0sGw8EyTDyKs6b0YhhrMw3PD3
Tf4kAkXZkTTElRroW5UdE2nKV5nDkGYYe1fD1ZfjYW/WgQOK4cIzlVKzaaMGQM68
/QtjjNaIrOf1SMnEZZQ4E5MboOxBT1Lu2IgRQicUdrMKVvGw7j8qtzPs7v3m3o89
k9DEg800iphkqJlc6KstmiDGGHyJ+LTzfJpsuUvy3GDI11I7OYGxHD8FtUsPpF5B
zebF88HgCwJG8LKQDLDHZeHUYkGfNNvbG0GR4jXFqUkNzRFwJtAyRylGt7qhCZ4m
AFexNdnXzPkHIoddAyWCrTNoMMT91xfULeN3Jdiax0XRF+IAkWqMmPVHxE/41/3j
VO53FK2DovmS2dxBFZrSQd7HeQzacvKnvI0UQnaD0/rCclJp/afV4D4H49vWr2iu
mORhyNYV+Cgv3QABLBkk8koQOGCuWlwiLrJEXAn21Wrp1BxgQq1lFHcRDYY/Dlzs
DMucyU79O3aN7Q2r5sv2qNRFDaGqroSyCjBVqtqgHlLXNTo7WWI2rodZTb5SC989
n+NQExUYhj7tWamC5jsAvfj7SeolhD53yExWBLoD5FMPD98+Fg2xVHgAGFGOtbzc
p+SLaVX92GhygoL/MLSI5bhAp5/aQJ7ytG614+/SvgmsRjhOhheNiLDdNT6Gee82
fVg8TUtrZHA5S4XNX0nF1h2d3QeaLy1GokDtplWvqG129xTVxndcndI6mYHGCJyG
xt3WYyb+KVbgiFIe1l+uvjas+guqEbm2DMwkLcdo+0Xb0Xj9TS2rVu6Y056pwook
EHYc5dRNY7yCplrejw6kbwe1BYOulDZN27lKMhAFdcM3EjF9NGMNJcAeBmOxNN8v
AwR6gFXmJizISNRWobQBJEnuJK9f2yZhAUNWJ18eXN+HqEXLzUKJoqVLX2wBBMa4
4IMqR3Jh+UaQc7mT9GNrQVvATNwzK+MvZx6pPxyEWJw0MoKvigc1sj1V7ggJdhIS
qnOSEJg+MTSslOXjti+floXozsz3kA4FVcgpmpzzOsYWwShF+8zbva7/TELlGWYY
dd8X/1ImxflCRCfWyLRtLZ3vvZl54BPEgwjion1zJzSKi7RV1dpM+bA7/FHtx5Wg
d4G1iYZlYHtYSC7yL6kYGwc0kBFjsQYMeyKRqKZQR0Y9CpWD+jEXtjgrHcE+EFXN
`protect end_protected