`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 23392 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/59UwEX+aE7FohaWu0/8IpTj7mav863zUNIsgIH2BWb
Abd9opeuBjbGF/waQMI2vMJTwD1ie1YueHc3nSNpEh4OXp8P5ybZFY89uyGz3ztU
W1EsuUnchJoQgbHZ/sLbgtGRgsrAFn+ZoIeGN1d6RAF2wAESJmYP8zw+p00RvjZ5
bq6N2EMRDBNjFRM5Aaj5PqPvoQt1metcU5PQjjF9bbKgFeetN3zXwTSVUPJ5U+5R
dw69zrmJJl11w76Dlmyq7qNbPCQj7d4IGYjBfNgaJ/uT30DLH1DJ9+6zcnlmD1tC
Js9TsGI5PXSa8t7glQgvfLsBaSQa5KYA5kAsdR3IYbvRxd8jgncACRXq8yCGKgTg
SuECh72romgG/rcdvZwCZTNq35Vpwoe2GxosSYqrjG4wkpgnZx/vm5ECHAyV8MJ+
vaEF8RlphgJ2zl9yc1e4GqMbnskSoDchkxhmClM6zqHtBKT8Y+AguG0ZGlTVGjFv
PXFHDUB6X9jxL5OXrJZR3a+S4txncj7+VullY0OltxEK1Spw5+SRet1Xvz6XANJO
UBOzgszvQQSq1wr0ylTQzbFxCaa3tTqkr4EV3VWu22V+dVT3X9j9zci8Xacrh2T+
tEaTY/8sB/aRbtmmbqE7OSJUWKJWpp2mv3pwq1sv22UZ481eSK8ZK6VPDynNpqZI
ZDIUQaFdAzg1y0fn9DfGA7y5n30s8PYozQKdVWb4PJ/G0UPcaDGIRTFtxA3rCd0E
9bvqCtdjwB7rujpCXsKgOUEbb8YKct9RyqO/Vn5Vz3r3P3KXVEhtiDz2TqkhV3+8
ecMnOHlAwzU2F2woLzy2WHhOKDbBVnD1LkgN3czVQ3IOiaB9PnJ1gXlpA7mL7yPk
wFWVfkBoXzPRIRGjjqhvLynXcw/2tddiNuXUl907LEdLGqK3N8tzVazXDKCeow0l
Ne0RSuujHvAQHTIBoOI1L/GcTFxsrxiwxq6XqRM5R3ijA2EbN3T/5os+dSxuuMD8
uq90OuFpSh3jO1hoFjJTrvwYz2oATPu/hKsB9mH6yFB11IpGwjW5uaMnKe5EZRHy
RgAIBljcnNBzT/sfpilGTjPHsHU2UYcJkqeA/EgX5nSbUZ2LDCNwtOe5pOWh+L7f
SznW1ig8bppRIcRnXnGEC2P9mS8YSIUBGmzko12+XorDMXpGcCRytqRnYnP161aj
bHLIf2PfcZaoHy7ADdfWVjqZCy+wPfZHVGWQl6BnGBj0ZZIU0hLG49m4aNG9ilvN
hSCPYicCR+YdsW50lIgGF1fmlHjaD6+S0FydDN+p0hWC4cuYhi0iPa3bGjUu1KGu
Lpgc7JlHOi44DygUw2b+ShpvdOBYuxvEBPNYo6IalwvV5GQKbNZBmuASydQRj+Kp
jTaALpdY9RQCxkinCTCza7wyQa1THSGMH7IyHGpQSaMdzDnW1ABtxWoF4mF2NvdS
udxRZ1oSWgPFhwanvYtOaAqeiv9OcmFvK9rQP7I0+pj8nEXmOblYVpGwCyZCPaNm
6VGxMsL7J+1OQdlbW5LRO2k4Gav4O24x4T9zJBnMW+QTzW3751lhDhJ2nRLXBP5X
bFv7TgJ90rMdGFUZ4J+Sgtb+/MDcbTuwKvQ/dXadkkcZh3colXDZs2Jv32anr3S/
/RyTW5gHjhvnBATUudIjHhnS1TUoQhChRe9NjY6l4zOClDZnfNHjwZK5zDnZZrhA
2ECpyBNtPdlquqsAwaz05NZF1jMGVZZ9XUsYW9GBaBl6UAig3T532zp72wd0Uhb3
jKOZRRRAH7RFZJQRdUKobMt08MeaNfgMxXDh74i+ZlXqH8nHdrMVLHxyYghbJNjj
ECVcZkMldUq2Kx/Gd0h1cJOd1SWlcY274ikWaCNWiPh9g74jL9JBsmC179YiNWh0
GAlrrcbxaiGHsGuaC3/1imcr8hhsEqEo1sdCNrqJwGbpbrhupTol85aQU/lUEC+z
73o7zZpbT5ifcqrgfkZ386UjLz7sJfnOkn0A7pQcGPpRsldaSeKacjEFqO145AcR
/vKwALIxM7Vyv2fiYlQuKQJQOw8pTMfwNzkV34vmFKwvS10aVAyx4LwwoySeC/hJ
a2v2JBM7wXnmJx9eAqQ5irXKR80m+9zXxRddhvy/4GJTfBL7XzbNnMFff7tJWdmu
fT7c4SyQzjA3+TbENZW2obd89j40dXKzg42VPtwlZEGrKd/p+ntGvgbJcc7JKy8t
9KEc/0z45g6ly9lcwBuxuT0hX9uMwsOP1+ggRxL6UdvExjKDOICWWSiOxQHYdplg
TNYr2/eBXcLwDOfmi4os/Q0fNbnGzlV7agPS3J4CYE7JoSlIU6R1kx0Lxe2xFn+D
ytHc3hNCK04RbStnRLigoWv9uL2fVXMybtCzD0v9iEcX/zJ+jobi5+LUrkBnB9P0
XtS+AhOaS1dUmV1QQ/aG5WKyRH36A6joiGdzDDJ9MRqQYtsal9nfl17OSsEBmT+/
Lh062GRZAYOZuu1azDTbk4zca5C7RChJ6GXXXIW3uPxuxBJche/92yN1j+gy5vze
BMQVCY11mLNtxN5LiMwoxXVhdsvh5cCTSBIFM5CQwm8pTq5nzpl9aHye9O5ZTWy9
6nFhIkXfQ+35lLRiq8Ttxq23TEOi1biA/+yCde2eZz8ED6sHYzBc5ZqR/V2NN9Ue
NjUO8qFPG9p/gIXnsFp85jVQezhISnZKuuEHDQv+oJtyhfb3J7masXIj4VOwsHbH
yR25/opP2FlUAnUPv1Ed0mzEjMrq1EWr4GKY8QF8Km4HyW9JkuAaVsRCfHm5xHwQ
P17n0vOwnBaCAqfp5Rv/3K3h7zaq/q7SHWfngRGtyxtHDvLop5zgOH9fBbdXAVoU
VOWkLGSQ3NIVz1WySnsYfBujbqn9KponnJ8oJe8gjNjO9qn6malnFhDgGS9yLSnp
IXYnvo+Fl+BAirWcYU/d5GyCK6bdWc8A0jvdEqIEOJjl7XdPBQprLFpVPprPZ9c2
aq1QZV3Rpk6Q90X98AoTeDXNDA8HobMKrEp5O9pyLYKChIoQ980Jxcd8NM46bhtB
GFQfvBdQNPRGvvJHxVnP3Lx2It2vZb5DnYe/+TYWPz7npuXHQiPbHDsQjV6if0QC
6XGWpK7BCHchFOVHbsggex/MxiPjwt0DR4Ku53fGY2Me5WulwqBJ5vQ3650tCwcd
YzqO0Rk2TgjnfncFSeZkn00693GJbxAMNivX2wwhZ9FMIyNn1rNiodgwrqSRKq5V
cknlYPi+8lwPGKFpMvkzeANzCF+q1Ltc8YCprne1aklLuz41exkW8WhhwZxnJknv
m8gJ4XCLTqNlA1TdwRNJnHpsPl/bRBGFLK5jyQHp0bCsmwj7H3jfOL+YS/KLHY6H
/Gk2NMIvQyZC4DSgjW6VQV2foKmXK9a5Dz2SHAo6LwRO5DKpmiEQQKm7C20Q2wtT
+qFZ56QL9/MqXUQChU3xOJWsn2sOdiDzeT0XEnoxf43nqWC5RRRJB6eSGHIGgm+e
5Y57SC4MiaQ4f+WgUNU/Htj/odMWHvLxVu8XoNo4VgjVVGahwgfzGmcplUC8jqIQ
V9Q9YejP0Rn/lJA2N5KtJtF68cKh0UbqV8FOLQCe4DlYZc1vxQGkSauxq82hDyv6
Ku9zyoMAiM9RDj93qrgY7esKXFFSmOxAYrnyz9esbVnnsYoI0iVXA4zMQAR15vkQ
3/vriMW2EPZstavJpq0ZrvBT6edBTG0BQT8VjJ9naztP82Zj+ESMNJOoc6uT2vFO
yBo4L+rF8jvh2++WAZTccCq0oPQQPKxiovAjEnOTNIjnBzUrCnpF0lFzpHq0wFQJ
STYn4ZtTjLz6nbx38Xuf13TQ6+/gWM69ZRrt0hzGdJC5mKz1EJ16/xPj2CYOb6jh
9IInCbBpAtyYoDNt1jPB6wFx5YS2mm8ItHvzLQNnCG9s3jDvOf3e1q5THffPKYiT
Bejj3mWs2kzNhArmF1RBaor0MWUzeB+OP3o05lJ+ozTHk1ECm00c7gpxO22md4FA
i4s4HdB8BIxH5UEQ93Zyn+DzQ4oHXYLMjmRom1ZXPiRqAuBGXDIsOg5CMxqcWq35
9uZmtHAwScs2+7uGB+ybVh5sGOZvJ2AtsIkXz9KAeyhGPArzqb7V6NdM0MF3FQqh
o74O1cCop6Go+vEo6yNaQnvG9fILz2VtSAY0mvxoOS5Pr25UH5BioH3eQJEe6gTb
WTcGjeF6CAwVNbBpg29mo1vz57MDWQeE+Xjk0FWefuS9SgKe5ZaDamUrM7ffJ7c2
1C0K4llD2+5ALZfH7Dc/NuB6EG9XfUwOi0KGd0VAQbRw+Vr1PQaHV3e2e0pPPT3O
PTv/S7l4Cz9ReufpGUqgXyqwf4Rr/BkVSQmQ5DnWD58l8n1l0YeurzhpcsH7lI1w
rlYtaTSI/yJrQH2hIb6M+09EGYrBNqpsAEFBfsLqeIldalyAucZd6t2Mg1JBN84R
rYdJG+g0EPvJZ7iSQtRdCqt04zRS82MoeYFskd0j063l9/MjjoU75OPF+I7dBeSR
1NQhQ0qiyKJlMrtSAhEAlnmSSYg4hyyQ0ZKSbXG59y5X7B5LcFEZEt1Zs0YvaoZg
nx8aTbZZIXdPa8F0dHJGMHJB5ctMJdAdm5wTL7jeX0S17Y2Cxdjr3jCVjOXxXwUW
mNy2HYQO2T4bzJ0nhw/b2Q4ej9zAtkKfK+YqQJ9uxgKyqs9I3xpDJtEAVZbZ1kUi
+dTFUBHfjX00y5qHiz2X4ExfG472j1pbLYIjzsuQlDm/MYY96qSFnVOGjhCmfnWc
EmJwHQEmc5os/gRmxQKzh9uYBe1/3qMM56wcFYp4PoDSxUSqam1DLUfF3fzYBB+4
O5PDlVGuWCSrdOA45/A2/mmvaZhYQNVBVvEmRudeKmMayvf3sa+wbvFxKlJY3kAb
uKdiPM0hOKR/NNKfTytlp3yl1vis16AMvKSCXEu/qCUBj4cfQZBJqekUAQSzde6+
8in1eN+/3nAPrV0no8xT7qltvNTl3TgGRJmqNZ/OhikuOhrJu64sJyhndXG11Pwo
H9pfSC/FqULLd7PWWrl2xpP9feL5QiKP92EuAuh9lubkm4s9QMX3ryeKZKmrtstM
ugW2zOn1Vy72zwJYJ6bdRkkAgeIN9vFvDvDehDVPkLAPAaHwvjJHOPAV63W6L3F6
XPpu9ShZvMTkzBcuRs17/GYSdwqO1eZ48rFgKmfvWslgvAjrd+3ROhDwWHAFsBag
yaLxbLtEpRWTxgD/T4MC1geLTn5B8PrxIt3IkebTa/mgeSEUrVCeje/w3I1XP/FO
I6nBdTv9ggnR0+8ofICV8ukrHidKb3tHgr+UteMw3TE0fzTe80kNa/Fk03/j1M6R
DhuU/MWeC/FeMwvoXAXrnae1VA+/2gVxVC9aHAgNkcm9QXg20aIGB19X3lG/LhoU
O1sVtYS03OCwsyWnpdM+dZ8NWchDQu5IKTTaruitEuWdvUXW6zSCaaWPJoMjkNfF
NlwwKu7AbLCw6ygV/Y57R4PfyxXV9nhJxN06vcMijhYFJuTCRmB99LKh5fgeSVb9
h4aeVKwUn5/JxtuYJ6PWNA/OnPQJhMhBDB4UaiyQEPCbrwrfjCrZyGKMr6O8rtEj
pXYCLtPE6+k8ZSrYxVQ0eSyDVBw+4IY4UGNjwtZfr1n+Qid4yj+oTOGxS9teG4Qp
Hbs9LxVgn12cAuKeOJ0T12Qysh6Bk2pq5twUqYYqvgQFU430Xl5iWT/xG/O1BEsu
QBRj5KOPvx7TwutC3Tn6zL0Erbtsdi1Y4TAoqk+qiW0KCdpYlNEnmM6XvI8OtnRB
OxvcOQrlv9xwLxlGMEl6FBnVNVVIRCY4fW0cwsxj+ZEso2YtNVws1VgBT6umlPPQ
yl824TIS3nepfzpbbRt8yEHDodUycc+Svwhkr4Zdj9z4Tl1jjZyRY29rNEfaqRXl
fB1JDfcZcQeSl7xhLJQuV8Z3o1zRJ4whIat9sQxE6NKkufOGV232ZvF4gxz/DgYa
PCWCq+jgUX8JAHXRU53wY6WuerWE+CzA2UIG+rBExospMNAFfDmfhkyLY3RnfGf3
VlxlavKbacmfCGDpUFKM4BFjQW3epz3bIH1s98hF56xv+0nQaiYc6VSPCDLq4JuJ
UjqPWMuRuJSF7o7ioI09OUkQHq+KPqzGTnU7zxKXz4Z3wX+G1RTYJt9ByZTtEKn9
5HVuykaSmRT7+8an1Qyd68cJa62Zqmb84FUTGWxjwJlhunxAVOVTpq66o2DPG4vm
VIVSRJsMXaw0dS01izATNFc4PpXxbnce1kSNmtHp4NSqc4k5+QBDR0AqC/Si9QyE
4qL8Y/fg8n4HZsuAplYlXcqdRcuJT0XQtxPguREEvouihr+M4BTp6yQFeJygIdyY
hgq0tumY8v8f8HalwmUTjbVYtTBIzByMV2AN0ARHiuvoJSKe7FsU8Pg58TuwTW3I
sKjCoDxpWp7IRVdd+m1xwRYyolDao4FIp6NX7BqxnD6rjI5tx3dKVlzSAFOwYZw2
x7C6JIwxYoNh1QbeYGOguDo/fCpjGwVY8rcndTwahgRA495r1F8GxkypLshZJhZI
Z56SbzgW4InPwHXRZCw+kEWuOsDzbSPzugrcIBt3LFPAVFn0myvDM5CAYdRLwKbD
yYGnjle/8NY+i2eJSp71RsS41bcqxNq0+8COVqbulobFe8WsPruU1Vptn63wAcO9
NFHaM5fFvYj0mmYMEoQfyWporFiq84udCLegMfxo4uA384tcjUGTuQbc3G//ySrU
hzP1VQ2sh4yHK1+55Glhcr6J4QDSZRQMqM4/ukGGdt12Ul1Hmxmou3tIv93y+KtI
meh612utTXGMR1WcAUgQ2jQRltJZD9b7ExJxfuy4KJysztB19rSnp5wULnhST2MJ
p3IW+Njca0bpBxoR7U9GV/ny7LbRvllf5wpgKMHEUwr1emIQ9JhxDmeRTN5omif+
iVxkXzQwhxjdMFY3CqML39GYP4PmkI6zI0Gb8Yj+MvJTy1h9jUmeCH+GvAOqc+EW
PLLIwZ9tnNOUhOoUhZjpxnCLG4ElfwUuA/+av/cl3T5vLprjUHo/1udkIVbCEm9e
xTtoBJzX13AqpEbfBAMQeSK9ve1kaV0XbJeM+r7fLxd2L+ruloMt3USlS6zbimSC
GUBDUsL7DY244TwHutOs8wybSFior/1DHfGnvAryi0zggHdk/pMEc16vuptVHSOq
uyvazYDAmuAkohFLsimToqtMTxejjoLliCI1+yDpGtYQVrNpuOHnVusunH6C3sjp
iKnwQvSaIOo3dwfudHcPLAquthHVvvKAxUaQr0OxLOXpaPd8VM0m8wtiZ2/JrjaU
zxBSlCjra3CO1tZCeVAva3VapJn26Pk4tU1Uhz8Zu/O9L1hmY0PNofgxyGH1kkav
YTsuB5snDuCUCCS83Bd3HEiBOZqTrmh/08iHKPks7rtdbmOfRecXEOlKc5Db6+Bu
Ns68OrJJQqwStxvEBnZAlNo89JvsIskRSIwGXjsc2HbO6ZFlU+2jj1DVren1hkcY
y7DyW4F+DHP544NfAtCiJv7CI09zsbiie5iA7XVETwGVfAMM2+R+egzjFhgCEM0a
huQJXFlTq+0Rev5RWISM5ksCnOA50W4gtaicToq3b34q+YhG0YBM8evGn1R5eVu+
lCUDZUzfCwBiK9oytS9oThGhHVytBClDDk6yPeRA51QaXEeihc+ZqfmJJxxCjObW
HEgGDqLLv5HsvQUREI0P7j1E/cJxh9KxWepmgYvLNf3t3lY9aQrXt9SVUbH9lB+g
9kYCohSnyRAaRDCeyjrxcgN3Wg22g2TcdaCOdI8CsuNe2oRvvbUFi3c/GZ7T9iTU
hbO5mB97bLVWv2q1jpRn7sIiQ8Uhcyn2cm9eCy/nTV62lMZkcbseXli3EIh/Uh/l
+m9IzOkRU7iMDHcbgAcnKzH0GL+5uBSHT5JdCBy06M5fjDmiA3hiZlxLYrfXCH2u
Wc8bRG3b0Vgb8PWI6G5LVJEPht2CjlzB6RtuNuC3dopP56MsAh4HQJkLgCMPmwgK
yzGsTuO6D0ClB6KM+udvaT2eQpFDqnoye4RXR0URGJqQXTShvtcED7zNq6xWuK6X
K+Zve9u6zXasAonh+YTXCGcfEwcrtodgba5d5qHlvJWxJvawziaMUEKIJybKdxPP
m+KwTEuxV5iInDNX31ENsw0kLNf3uAbC80HLtcMdVQ0OL5Q0EdLV8HxiZKKD4vXb
ICqBCJct9Z+SwNEGIjpuB/HWImROgJ/TyQ9Ckkh0HR1CUZORYlVZzV6qcm0/zyJp
stKOMuVYSbjzDGACuFq4JIkklPCkoS2uwaeMVPFCVYBUzO1isB81toJPAMhf9r5d
Q6oO5bHsy6WPwyrZ4GFSS1KJ22oP4OwIrRSrX54UJ9UA9aBGHHSMG2luartViwK2
8ZjC9KA973zDqY/V+j/EKKwUzr0c5bZh6961z2iJKZkMoXFK+UmLMN5srQra8XWI
y2lzIW+NrMLDY8BpSpUnBTV963N0FuJuuBSOHb2Bt38YJCMM5sXhGyITeQHoqqxe
7FXUbB/NJhMvDraGKkQGIZDPYR5Vdq1PVIR1SfMOMmqvePmI3bequ2z6ApCq5H1I
Kn8v2r+hYF6nOAUHqgi0vwmZfG1zfSzG0wSYo23VKqYjdSBQHTr5DfknrchbTMBa
40oddiD2Nz5Li3pYjyV01sPFX/2RXhRCmVZQL4lZ3BANTMWLECOjdqydgBfNuiEp
RYd1xrAtBscESDH3iNJIMJ4bsF8LG6sGL1w60S5e/x0PVhuUYNvMecNoJAd6JvaX
uXEe4ZGDbqWj3yXy3Mn5N311YaC4eaVPbo4x6YfZMQD2rDuJnqBKuSC0B3X923yp
NIkjgdvnBy68PiJCrLZMETNKiB0AamFGQ95bEhBvT6JNUE9qQ7Skmm2f3iOc/FUX
PxvbOor2N9FjNb1lwN/NAQeggmR0Dzqvzds/bZm/PRfO18AZy2vYBWb4QAQq9yCV
yFS24sp45cn12NeheRshJCqzjuW1RiCICgQfggOv+nLIvPl7u9K/Pa3qerKyxn0I
lzOKQE05BQ+3QDKVBrFxISlowWkiNJIhMW64NHjVaS7pMuvh4hz+0TLB0NGJgaii
FUMVwv55jZonPgidl8RbvIBJqtvQ8LMk8PRwrYSyuidNmv1Sxg84ARnLaVP4sHQq
TdLUh8uKDmeJ3DVZS5zxlp9P8yZqABJNE4P03ze2CKHMEeGnP4AsTCRtoKr03uDV
mKCNlWMEShCjGe/0vlbagrFC04AT7ud/j0h0wrMiNRktLZLRhuNqzNR/FExM+Xtd
MkYjOCoic9TbB6WnZJ0dln880AD3KO/mChkEM15ZlmSyEML7qqN9QHXtmeCrijJr
UA+jvTuxooQDmLJWy5cF8OLQilOnqVxHAPvIpad21CqARRxS7den0kNKR97zaqrv
SeBOz9T2kbZy4qTNoR3AXv2g+8ZNkhmvcW+ZLDOggE2pfas9s0PUS6Y/ik1AKXnN
W+yOX0TGfrF4kYVklhbhjzD9erDUPe4o23Qntk0cdQgyY1+ivzj2hIc1ZqsYXEvj
PKWFkbHdN1Rwim4wLuWI4FeWXQQJTAAJo6/RkNqZ3/DZIJJ+uSei4OzfFGLqbAu/
oFnwuSRyixXD21ZCVLLnmjJo6atqJpISfhkKAIDyWH/yW7smDv+vJ5TrGAScMinh
G5qQ7eAMRYN9Fs3sm/QuWG63H37ZoS8HvELV/LQrxWKL2Q359mmzN2wXFjp/ycN5
XrNIeeHK2ZRmihuAtVia6pJ2uzPhY1ppE6Zvgyjit8ZspILb2wdO4Mr18oAv6X3b
rAvMOw6LeHboX7rQ0xFLJwJgjNyQFLlNFqppQbzez1M9Y33G7BNdeAzeVUz4s1ab
RabCv6jicQ/mmBXTv/njiktEc3p7m7uX4oQS8NOjM3ccHv19zxdoy9dTD1y4FCHJ
c8yXU70Qe7LduuRE3WR6Z806HaEfgh47NRyUlMjDblGZojDj2z4bf8Gj2yE4RRnu
M8szbP1oOy8QBUrdsQPsV/9g+na7XSDYJ5ZLLphwcGiH3sg9kd7gNFdp/HV8P7js
9YNZu1Xqe5IysiW8S6PrYmIHX8dPrxGE2qEzKu9Bf2aZh6gnb9D/JlH9yPsUpt4W
SeAeftzWW5+a/Hmrq9WbAkpI7CIue+y5v4wUvEPE5kL5f6iIP0jeub9DFPGUUot+
Ezkz54xPuC5Eu19yWr2hEk9+pV7hYi+xSroMmjzBF6zYr+KKVkzJjltn50dEnlnK
TLZQQbZtP2x5MI2nCMF3xL+8QpJAMex4Z80wDL1dBLWwcKetGn4BaS7B+ETlGrm/
CMstjycUGnLNj4MNXMU5RJAF+K/DrM+sbjc6NuvcU/a+mgWTj3ZyVzHvY4yAtTZK
VliZ1FtsvvHBEB3xxyGpHQCKFDIkrilBYyGxNWiNA6V92ivcKkoz6hyDCYbZ3ILX
SxuFxQpk2NPbZU+L4iXA9DbVCa3fIl72rtoAaqf+I3FJq9ZqcCE+tFGO2k8hzUCE
xkZQMUtZu1J2404F4EALN2Qv/Dvsp3BxTgHGyGkadTrqX3KZV0O5yifkeJd2y2RE
Jb/h2mKRfNBDJ6vjMhAcHSiSJyvZF+DpcnJkGmlbbndpf2IB6tn2/yRmwWd3bLC8
+KSdNEwY47MG/H52oVKSUyiunFcwlEzFtCgUun3EuLSFn86OJkQ7MHTQ7Wi0pnrx
A+bW6uEINrYDVBG8sdquHl8RpruOiFEIqjEReA0lkFTHwxu9nCX+3QO8vTduSL78
Fp7R01Ku6qwZhTH9dBm3e+6GJnJf8RbkK5lpcpwsJg66ToGgpTUD3WX0JA77xrKO
6HqkuCEr2quM8WKYJQQEtlCLQdHFU7gb1FJ96cyYcGRv6waSU4L+ztCqXMkTn9s9
pTzaoDdwLKrVSbCmv9OJZ7YLdoDu3a6lFD1YcWJZG3g7TEDlw8BKd5YhoMDsJtzf
laKsuh8wFzkBvcjf3rByW1xEXVh5haR+keREbyhrcd5E2jsjvCGvlHcOtPhUZWPW
59VF0qkqEfgrJM8Qag9vGbWXFsj2MnP31RAYrwBPh6aQdT3KSofDWwlrJcE596ZW
NESW5db6VE8u7z+3PauXkNmt6Bzutn7z6FvMWQM1DNiyEWIGhAR7XC4vSThRaESM
Z4+z3HwM/b+zVc+wH0sU5wYRkIrm0V04tDROCsmYxWROKwOKk3stmVl0KTPAsk/f
AroMeNYXzOVbXJ5syZGm3zcTLDV9bKJUNQqWUXhGf9+KDcLHCnmHmVWRrKO+aeVZ
iB60/GxjX3z0VCVJC6uoCYqEybp6iOfo9SoK3ZcZca2Cu73exSF++ebi68SI/HIV
1wsE6XhWXo5d5wApWoK9NGteEYsNCiF5lxfwUFuolsoTU+KQOt7D9q0OWuT56i6x
0rcRJFVH8Gsj7fOP5VNR7VfWSULDOlznU7/Cz8B9D2DAVungZdtxTk9e5KyqTV4s
wfECS5OinFH5OcFlie2JGepZMcWrUNHbC3M0JtMhyldqkWz313xn8T2ubVL6vCWz
wiK2u4MAjqdDkdk1u0PYf58YNq5WXG3xlm/HBMy7goUqPmcvvWyNQoVFskIqpVEU
zkYZLK76Qm34PaHNyBBzftyPsVbfgEW3p4yCI1nzIHbVtLe2JL8FyihPr1kpu2kJ
he2Fv1hr/h95Kxyi+WyYs2ehjeor/YYVwrTAmm4hI9zCfI7vd94TP5RhB/7s+aOW
j+MRFYGhQVzsIG9oAT2SYSKTTNnCB/DXzj4D+X2EsMsZdNLb6cKmw3UDtiQ5/CRF
PG/VvjGRUMijRIkCQQykgFqUa2MD0rOcdnKRCJhQUADK9tbtzC9b8TPfITwm+ROS
cqw1v0QGoyAL2qybTKDe18kr5hIZccVjCPwPhfqtcLpd6MV8Rm7v2r6SqTMO9+fg
yOkJEiSUoxNQGYy1sE/WeoLV7rbuV2DSFGnMdE0YrqRy+lHQ3/7cXfTxkqXQ0E9r
dngdjG5zWhJZ+15AjKzAUFDm2i+zCk/KkJB4Vux2nsjyoDFTnMAIsjsmAUtRT7AU
xBi7ia1XKk5fqHVZ3B76C3L2q9ZPf3Lrzq6esvyT7WpKkeC5ANCIjzWD0yx9gHSI
PHA9DDcBroa5YDuE5OhgIJBY3P2pom+Fd1vRq1npvX/hgVLRhMq9qJgVbV4RI0Ye
CGgvE3EddKjLiNw2DE/sn/MeaerZFUcr/PhoJjqwISYOGsocVMckAeB5fCGCNoey
dWypJIr0j19J8jcR9IRqpYTANci2EaXITBKWCyJH7dgylfVU9vBsrw90c7x2Hf18
UkEhuAHL/qxXYw2ejO9IvtUMk73lZgc5FuDkksBcGf90z3dEgWCBQubeWewLtGuO
WzenOP0crERLhtJrhU1h4fPQWu5Y5HjwuhQiEf8oOMIxa3mVP/bDVezlS9p3z9MG
LiZErPcKw5i9RvT5ZEAb4J4b/tr1fSaKXoTa14pPx4mkHrH1egacODpYh4riqyfu
l3hZBFTuZ3gkkcxgNj5xsaEM5b0C4tWSBzUxiuEmX5+x1m8FZkrt+HBsM8EURCF8
RnkSskIJ+Nw148crKaKBFYgABqS8wMpzNEKliURCBJ6kUovW2jNZwE8KCsySpHGn
Rca7NywhAOBOkx6a9AGIJmmADb6OAKpflrTzYy1bhLoyuOMe3/Ot2waqYrwaL0YK
i/F2/xB5s6YjoRpF15sTBX7D2zx2NFbTwqaXFZYsiQ5dLCfKuvFOy7PJWl4xcWM9
vcjRj1nxq8se6sqgsGLbdb/Zrs92s+X64pgk81/jam1z86BM4bSYp4hxVfR01XQU
PsPcZXNzfaRB8vM6LWwVzfbGZm+Shw8ytDmTgFBHbZbz993n2WxceFDOFhxPixyt
5FUT+uvje2S0Xl4y5W3rHC2jVnfZHlc1Ej5T7+MW6v9CYBU8vGj3iWn0Sbbf6Ape
T6Uq3XuX2qcpWXA6VwVHEunAQfHk9EPNSIyHmAbXJucOyb12OutOn/O5eLVsuoOL
0QLbT4NDXbDGE5bPH5ydkr302Rbpa4/hXK3y7xHgM86/ZTkmHXEWLM37pyi2LoSu
pLiQa2U1fg2Y1YY/qMohV3Kp3uNT/bBk2e+KoO/3WUg6Pn0IJrzFPoqgiiRMFF0q
GT3piNaKh9wKtVhg/9Cf0GPt+jnGr68CJXgVr33u0vMGgKmZ6lBqip7kXE7xpa+4
6q4WLdMgdSMcpRnkldopon1SPg8AeZP88mKGBlAYRKKtwdbW9MjUsfIKXGrgzXzc
QZze63hk8hV2psDovr/wluYklDmmykSX3VJytX+MXaUY4TcuzMZC/Z9ZJ/PxUXAO
MNYk8RnQa60UCp6wxnF6R96ywXgvOZWN9Rg6kgmD5jGlQa/ylnk9YkfJpDjVjjYj
wAfHuGeJDaSzPFAJpIWkPXiUa4hyHAtWo3wQAgFsn41mR3qrg031hpSbYOhNKrEx
MdvqNrY0kKLf1M35SIPpc6C3yuSytu/INLeEESwpu5DxENmqUoJtQxM4F+u1tNHj
xndSnawLujBfGz6Dydg/mJZdhisFpgv3EhTe1JOc4CvyhHWB/k5n4i2Ns9SFvXQ3
iFkiHmXmeSkNn8qUnBpXnmFv3bRurDMcu+G+E5F2OuEFmgCBYN42C/pDYoVAZCL7
wKxgXLlOiXDfHkMtkry8YdHjY8x0/W06/FUFTULhf1bBXDNPoKBtsBeCWp8f52RV
DuJsA2aUQTG/OP1lLONiU5aAaMqa/dTT3nGuKFeFUxD4CMze9nDixtyLXm4ZaUBX
itTPwtni3vm6j+TzJvZSeTmz/wo1xuzUgdPVSZul8Dq52Pple6E6bb5nzHspOc4D
llqkc9jKhf7yQHe2yN4CKlsXlqKIEsMa89HohNuM8tXyDOurWpy14zkZNc9wOxmA
Y0mYrmVPTQYGisK2zLAPiXtl33RNefLnMhSqK8qobHLYxKHZn4PbjRQeFz+u85C+
KNz2Am2L6tem9xxP2CmqDkHSjXSQzDKpacOKoEb+XbNCkY0JQhK3FeMZ1MY7pCgu
cZzkZ+UyhmKkjGUHyPir2d9Zhsh1jzeu2bSKN8I8HA9+MrIACRuUaoateT5tqsbo
dyCXOdys1aOaW9apK88k2aC2+zLNbHdmHCbZzpN65YHt+zkPH1zy7df9R/k8few5
9cB30YMoatr7k0ZNgfubb3J3YVjAzlH1RviyTYNzkFMgNQmWVywoJIgVmjstnFBv
HzVzx+t7qzCYoOh4VIVNrdywy+pxXXLysGjc09qcQXN8QWNSv3cHL/d8p8V3TOkw
azURkCqghAQuiCqaZceshRD6MUnQ2UPLMYUN1RESa0wR7BAJngzI2IO6YCD+2uJk
XmRONHKHdfSGLGYHrvHu5yzIivwva+KwMEmdfOfWucCRWVcyYTnJa87Pm4s3WMbo
t0VGatAn3BFGziL5kSp0lkGcyF7Xz0LVR0CaUu3mSZaN2UvZ/vM+oZg0Pgd5YxWm
s5LfzOzGkOQ8nrKiqDlkoVKYgM1Kzdx6FCnB6tqS/FTxcwhU1Y58TNqdWeVn+plZ
XD+xF6GpH4gv8AFcbALjHUuVUWisAnxRZPy/RW+dfRXG0cS3Eqsf89Rd5twkPgrZ
VrazUJn46+G88evjliMeJp2TgBLsRZR2mAiCPc1J24D0YJ9S/h/VZFyPili9BYCE
vWZaPZW2QFzPHZWo9HdAYjqC9wgkYJDHD9dCS2FT8j9vBORsXICE7CMIiTvePZpH
YfMglVXk+y+tHki9JViBiHSonSsZ3pdQSPwPNmoZo71brO1FSnvaMoCilh0OiJiN
MPHhN+RmIlHjPm1FWAI20M0Y3lbxk9JJbtB+cM3jFU8K32axzUJZkRjTvBRDNYMi
0R1+0zQVRmVtzvORTC7iXaJxN8P/nUjSKmrasH5F6LvvlIqEEALQGmwarLnVDmWg
cG7NU1yC1PXzbOSpE3xOr/UhzjCdn2TCdNbLbAugiBaFoqRZPo5oP3fSCgbciugz
8UqYzMxX4BYmQaK29SjAOSV1GOragjwcbetgUqBVBJOvLfHuQnKflu3pDDPJdv2x
j3eQvBA8yUezCoY1RnfE4gxuSKkNzZr2CwFJccIJCRrSJMoOA1jkvGlDd8OtVfsE
ly0+r/olwWedKFpuZg9QDtnq7+8ZBi/XuVnEpRpKhIc9NrQUCihDuZSvIgQBnoFO
VXiaK8yw8skKOjuze0RGAqHUsn2JCNagsAkY3EZ5cbn5nXQ6CYnR2Q1WvIAUNPIy
/de0Gg2GZ6lF3n/NZBBq2ewR/maBY69/6jqb1JirCk7fZ2vqDEUALNRBYcHPICou
9z0rQzDCgs3rV3ZLThXPseOF3FR8N25bCNGtc3WC1rW1pdi0zkogQPOpOucFnRde
JLkdLc91RdUAN95u43pxRUNP3NHzS3tYejlsSFSzIDJ5AFizmKgb/XJ7tg0WRydb
k3nZjMZvlk8+49HGMSysPWUpyWzMAi2i6ldP54NAG7FdDjkVtD/pqH/xfXfRtyrt
qreLSIJi6xl9swcyOjku0WtQn891tOyJVpS9mvjED4vWtJWf7OAmHubJL36udxXq
T156jmHev5gPQifdMntEilnXkCyJG99O9RqcZwa1q4FAlmAoKH1u4a2ARxFmyWla
ws57tT69UoQ9n4Ymlr6bRmLMeT1n2bXNTqy4hzWsy+//gXXBPnmAaTF/13DWnd/u
2Hw5sjLa3oWtba2qJ52mQ7M/gaXsGqy3Z1WkAjei6DQkDPUM3QP+M8ncTDks/KtO
6gK7d0TTSnzhdjCYOAZQ/XbGPdwowcZIfH0loZFLYKPU9JxzjPTQm0dYAourpsSR
Kbj78uAfUR+j5I9/rWFVKPkF1XIvqLt1YoYz82raVAxKr/UN16wFHdQXco/OdQ31
Z7qKES1VwOWHAAkSwbHFeNWDfyvoj3r58To+8J7tB9G4YF+LhEe0hFG8932niSGU
r3Mu+VNfh1OqN+1mDUCz8I1dNrpvsF50raWUaCAuqY5VHCzvbq9blj2HQlbvVp2H
DNr/jlfJURAek8yWXMTYmxwBhochW8A/u19eQe0q75mS2QPpXw0r23ah9UYK/HGI
91sWb5iQAmP+TLX6CkcYHin6HJTy4jucbzL0NPfaEwslL9Jei0wBmqwngDrXxper
Dnrr7YylF1WIGVANCq2RBxU9vO7gFp+qCjKfslkR9SYDOZZhYfgPK2MTP7MUYO6s
O2BifpgZFr81r0Oss5+6gT7wpRqVWaNqX0y1JJY+MkqbHalQF2iV33gknlw4IgdI
+YEel36pxV6CNyk3iuc8u4+t1bcPgiIwe5P4IPgJkHeFK+pxRWqiDl7DPAJhxbid
Ou52Uc38EOpjlLVWYM27sJ82OAS/gFW25gP3pIp6W9nsP9svxcwVQ0Gjzx744xOv
US1e4X5gevdXamdNISwNMBOVN3Sgas8xL7bq/LQCQcx+mc9/P3Bh73wyfbVbHugi
gMDMbGqQ9vDitfS8W3kLfeuMLOm/+u6AbReG36srMihtx1qMgYWaO4kbxaidzXJ5
BYcx6ADRiu8ztv1pttPy0FEeLv3OUQSTrNnGVDBWFW3xyesCXo2nr3A6g+e+xljs
Uag4HaJhH3gRgZEmkw+DPMo1O+pwuGlAu5EyEGMIossskqnyRp3usDBvNxZYNsRz
pIyqqWWxpYjVaQKG38Y8bBOfgeZsSuyOJNfpXXPiLnuX7YaoqgPWWdM9bbnnPv6/
W1n9MfIVlfd72LAP3AYSJQSHdR9qe0LyDkiI2PNk7GRAnBDaQy/zbdC4s7RSCyIm
lI9s3wUdVYqOWWGQhEbhGmxJhWO5HU7VgjyufgJwMJewnWxNTImTuwUcef+xZryC
WkBWo3avYAPY9L8KVJ+P+wSuVxgzCue19EpWWuJq+hM9e6lUshenTgE7FNFNozEY
A9WkmrultdwBecz3O6l3Raz16Eypf2xhY4VokLHgo5sR0dFSpVZK7LK/ySmXzz9I
VkG4/suQ8b+e0G5xk1N6ao/2kC8bVrF0NGQDemNbHScpVGM2OdOCir7qW5Hoqbja
UsM+gUxbteIIX4o/CJzOmBSNCCYZ6dj9XIkgzSjvmlKklIgonuzh0ewjGLKftdEu
KaB/hR3Uu2foXCMoTfxzCM96vTYCziT+Ew9vC7WVVS/U6KOPiiJp924aKi+ksMb7
FiS9pozgpgywMbwJmwsKWBSu3EvR/D171zJzFSgVZDMzktZKupcEBjnVbZH6TGU0
pa9x5rmkuooILkJLVlw8dZcxOuD/AOBqXV7DiJ8R8zuO5rNF0TvjSgRuI5v7a/Ch
gPSVoHajF/yYsa8ihR4TNxqut/Wkv9vXWTzSfBSdu4RsXs0MqqiSyNdPUtMX4pqV
6BQqt2yiBgmemfO7Aqi/DoVPxxAWfGIZYHqtwkdOZjpb/V+o0Bd9QsX6jXwfi1f8
n0GkcMBnFn42IDi3TLk5pGa3/BqOlvxLEo5WV2y01y78dEIJJxK0XoN2w3SnpTGf
r0nRkMAqBu8XnUIokilY14c/NG9i96XxDogSDCy8Bgw9GLeMV5BmwRBu4sF8uyO4
u0FG6Dt4eSzT4XXz4RCSHL5s9S/NbCQH3mvCMQ++vhKchJ+MwiCCPMug4GMgMPbQ
hegTNxdsBs4LlcCnkJX4kaK3VERbv+0oKYa4fI57oMVWgZYfRTBbauzo6gZJ+G8W
TAOMTtkg85dMHloXObcuWlt+iEsJwAGPfwYdCIq/qDXWbhhZXra9uh1NnlpFKGZc
/fk6TnqAlb1QMQ3Wf+P5vhxEnh/Kz4sZp24LeGJUSFZ7z4i/Cd1QkNQSOd8Uv2ve
Wcpqh0y5hajUF04l75PTH3u/EYxk79VJcc4OjkYtuWOAEteZ61TBDEP3pgzdhKCS
HUDIYLXBaZZghB7gS/V2B0P7HYzx6Ep/cumRbFeMhrK98WNqamQ0/YOku3634ssX
KuE0MB4XUEXLGL3IKw688uAg+4Sl4+2YQbTxCnLgKJckeE8GtARJcykdcL3RKRWe
937Ao3RTRmogZzAbXieuHqfzy3aAJgfiXywbFA06O0+BYUO8J7cBeU+aRh6Oo67C
jPQ6LwXnawElh73WQNDohPvqX7ngJFprOyX4aP7Z//JQXHt2hWg45gDOqtdJ4s4Z
Qh0hdJXqr71mchI5oVZSBhTjpvp4KQx7ukPZYWSvzpSyCcjnxuR4zVw92N8FWUre
jJlo+RzUh7mSxa2I8fTVIBq1WDqel5vZLqXX9FPpylIpqdGHdTFtQMOqpjvQ2DVx
mp+mcFQ62Au2jjgYh2LDp3Zk9ub7JbQwP0jNDAAGoRK6zXhBLzF7cEmDCQ3aW3wE
VYBTZd9AAd8M+eUaocCTCYNpIhAjw5bWSK9l3v6CGHQcSsiozUz+sogFX2jYMDos
G0uq3N5FJoTEFKdCj57JHoVvZi2dh3NRo7OWmdV4wKaHA+UHsWXY0b7HKqvMbm/s
eYmjXvZHLQgGKIaRH5XUJvT7oGz1Zu/nN1UZM+hJLt/R8aRuGeN1xsZzFXfczbZf
faIwYVt5Ai+PV2R7/49YSlUlgVmwZshNJ9bVap6vM8a4oA8DAPrI6uLTjQ4bn968
nv4Zr9fzleCE3FFbiz3bVAULLWJtjFMbLKedHKfPHrir3mTZbdJdWPBkZbxlSJyl
LPwlHW+gR7Z3BP9WKss6Oe2vK9yi7/WcmVzfkr06iM3eDEwNLTLBn47fsWbk/YlL
8UpFrpOXsER2hbsldwzIf/wtKWsKsdkIIORPrs8SKZFXiHTDk/1wc7bXpfJQJAoP
52FfZ/jo39HR/PB4wIBnMnZ3c3Up7Ja2iUQi0l9U5s6WS32PUM4OVjE6Xy59uh3q
9Ig6j3wbzQksQ7OiakBruvB4v7hfFUSI1LPaKBUd35FQZESFIjhX8ZyMxmHMGUyW
nnT5o8bJdimvPv1dK1go9AOUJ3Mv33czHgRZz0cZhZ3DZo7a7D3x/A7O+AW0RWY8
0uLTMhXRtZLYcvwLuiqPOgdCcTF7dCLj8VMqAlLZ62dXvnaZ6vBqvPwKO7BghpFs
wc+8RcrNRdo/wzLhVicdkUEWywxFnamahYunqfhMG93Tm3qTKWvlDLZVh7bWE28/
kHNyUdZ8NqeEB2ZxgFjrox47xYTViIXE5L0nqCg7z4dTASfSkM1q/iU8lBBh0jOz
z+H0jBSk1NB0v926E3+jltYkmFStRER6myWVKcfASAJdk1PDQ279sHrVHnmFNRjy
SvrNMGr2yPpr19RiJq3riT7I4nOxnklLVuBgGMTPF/Z6vJuiqtoqL3kGp89l131+
ceB8lQ1aLaEtApzgcn9qKyOp6Sr1G31xIkGeeUaPvnCYVfFUzoJ3FuT1ZgQ8zsUo
UdtrES5JnVni6FLuTT7bGTlVnQx2MS0YvQAEl0epeRIE0/KlraV5/HtmWdPsiCAW
RoKnDJy87bN7DgVfrdEzL9WUvl3RmORMPOTWs7VyUN66PKVZlrISRCgbEb6MWutA
36DffXcvYj4YySUu8RnZRFle5tNF25jD4pX5vvtqQhLQ/rQImuOolqb5GOzB+Vvi
oJwqH9nY98QNuzomXj3ASLfcVTOH1KR0PDJDWc3+SeD/JA/T2AHsIHf11ms6P1bE
TnU79QIDoL0FuzB/a62qDWvjUP9MU0yfF1AZ9/9wY3AD98x4Kg7/2famRvKELir8
kVbPMstnJFvLTMAzNhp+FTV1wKKHuYtQYhWXQckYG8xkFkqENnHdbfZBmKZPaZ9p
OBkspQ4FWYidsM6d8FXleZyB6CPA3DW9xh/VReCci9D4Es7OHI+xwH3EAG45Z9hD
djuTLHGdyXq3Z901Yr0tUrw10r/yTlXnPXGKtpMQBjrm495Wp+9tTIUUt72Lgi1f
Ap+YboZ5Yhs+/mG0YZee1Tvhh7DRsXaDQ76ESzZykkPG4erR9LNbVxQO3+FqBdR+
hAZoMUiNU6pz6GdrvgJJ/8NpdzvK5li1kIwgFoLrLp7e0UiFWOP4zlNxL6YX8KKF
jJVZCITG5fMdmerZur1a1/VDM93j1q99z19n16y3NNtVql4g//9yCz6ztN+R0yFU
9Nn37sZeGQ56DfcreXvgLJQQGg9Y/iA7I6Lzw+URhxQW1UnVgAkoxjK1rhg/+2LB
cLMuTwYXxVmbvZH2CwhYaedqmvR6ItKxaRwD8cht9q0vsT2NxIr6oiG1bN98zQRd
cJ35WQKog5ROa6VXSxpSUc+BWf7IZDjEfEMqHbGAzU8hTTXD/lLEH3L+GudEUmiA
llgnvUMnflGaX0G5x9CCl4OophfTBGzXG4IjasXPDg1Zfc7GehRqhfRlutl1u25U
2BaY8fxTv+DLseTDRxGG68x4REmZ6J5wkawS5VGMGjb880MlQ/v3Uvj7l3mVhqSw
9RtZ8dh1AxcqOwhUJPU+YFj8bciUu6zdRJSsF6HYk5hK4Sb0Gcm/Of6vUNyM4aSS
OEmD4G5yORhN3S3RowCSLt0m9FmQJkL4gWIwu4/2gOCI+h23wWaXUoJ1ddGDpg7b
nCNf0Fg5obG0rXSMKKfd4PbMYty+Fou+lDCG0NpwXegHRLBG6TubWyRjXbS8AZfT
29++wiVz6Fs0bVmt2VJAq3hoQzVOlKMnXJRzFjSNEGfweeqRckxjoUY7ScH90b6E
iGF3d6xWKBYTMngbMSbK5c2sohOskw9HnVvVMkKl5kdWGMtvGnElHA81uNFSO64N
JQRIV2+PpYfeT21ENjD02pVqoKDA8tHxImZyqI1TQVhhiU5GwLlC9g43bS7ofara
jY+3doUqhRx8iEOXgEr1P5QaR6iIvYGDZBlANC61KlO3vWU65U1qGtFuPS6S10FO
ZDyPUeozVBTUCG1EZYVQPOtjYEPxK2KS2RWMzBOr0IXW5mchQqJ575ixL4dw9uVN
7HJM30Iw3gGA5s+Ilf14M22Gw9YEFCpZh17s6Vey5+2gTsmH82bkUfOFed1GDdax
zjmL2JfcpQDV0MBMvItTlTuwDcBfFFS9JjL5zhkWE4Tbrx4OuEBTyQ3jTZIfcuZs
vATbhHAqJDkoOe+9CObQ0SZq1GJWlRvdhrqacQF/FeZgq18fY9YsM4oEmvEdtmZZ
SonIyFT058Q0k/hIkehTU2xmRUswQxhkQRvj2lyyCGb2WnOaYomIDAOhTuQoc71t
kLsxkyDM1FphpQH4EczdjyVRKaqpHDqfVm8IKafFUV0975TZvdNJ4i+wHdwZvLXZ
UoPD7lW9/p78encZg/ICZSfq/7IUIrJMPYfsfsUesCobHpQc/JGNmF4Qekn4xS/S
7TsanaYJ0XaQAx4qx1io+WOnQTGX5fKk29ai2UJmqLnkyN61JQ/VLRkIJoSuRDQ6
J0E8c1oolSnfAU2wFy78riSnIKsTNencQebTn0RDZtaRkFPiGmOdkuOdaP+dprxE
QLJJm+Y7Z7knRbd3egSde/itQaBG1hVL0khCez4ou05ELKZ+vRKVurYi73kmfowy
hKB2RnS/Ifx4oNj3JPCkYMhzpsghz8h8PfpMxmiz/yaX0N98ygOeNNCtU/Isbugk
8aFGXh04D870BfRVOAUZZQUsM8L02fWDL7+iWoC9no8HMK8CjvUWzXKB009aifRb
O+LGFwz6HtMdlQwVXbJctZG8znwLsEpjF/bjlWssLSrdSwV0/xXpjxyDTQqM3SQS
DCF/JKBmtV4Go6GvcK5/vRdtkMJ+kkZtuQLlKKLhCcxPd3P9+2ju90QinFuVUemR
75r2dDK0VKw2EmDzdU4MtFbafwBlCIrORU/6cndcsfnYOkka+78dbvIVEW/LVjpc
eEGpXXYxZYRJS2zzL2RpB25RlMOiZecD5R1PaDXb1xIyj2S9RSFOtq1me/kuALhw
8JvBUd0Tx0/1nMhXrMz92v1DWKPTUJefXJnkjLfjSsMeffEE8UWvxF8nNoZK6ep/
+xvMQrf/B4lKsNhgVu9Cq1uHoj9zrEzRIRsF5TpaXe9AcQY98bVmcgIVdfpyCgFS
JqS5oZhxsSunj++9MCefrAUDwVOtPFGDk5vFfC4NuHmle/LA4wBMnxMv+sOwOyrh
P9rNPyzSEXVkjvhpD4ZHqmUnFWxXncRICXeqyWF7peSZ/0RpVnNMUGQtata5j2Uv
tbkaoUkJXiMsawvv1c+gkpvY7W/TYzSju2ePIbWBTOQZFWilfI5RFk8zBkoH1ynM
hbQP0GNvk6fn5IaWjGzHkBglX6odZFqpQOZJKPMWeDroQm2ac5UOEN9wCAurfPOL
/OhBrTGWW8KbkJDPQOiyihhZ7QGYhmAe1ReMlfp9+qRY5ffGSULCC3r8U5GPeJUv
24xC3UtTL8cRxQBt5ZI7G8nubb/P2PKShDqa3LaAq3426QFX/sm7s9kUsDVhC285
1JD2S4i1bCTKIBDidlxKh8Hn+FxcZV6sD8wTj+Rt0juvZegNC+ntCQsI47M4N21m
SLZr2izV5vjp61vFCtAiwDCAbzTqM57asMj748UKzV/8izlHRLjE9hZc2OlGJaab
RNd6yuqYV8Z7p+iCJvfV/cGeUJ28ABcJurcAunrkFEqc4TfWEInQ1vvBuF+Iy3jo
kFgiNyKRX8Ahl2pRQ5hAXq0HX/1tKW3vfT/249E0KbWCnFxWCt2tRECdayeBmigG
GAl3ovABhgxDJS9f2WIuLhs+ozF6LEsYaLyz/7ww7cv07EVT6hwSOqt4/AVWR+oo
ZAwBtdUN5k2FwgEm7dEDgN3h//ZP/q1cRythfotOaJr34b17f+nc1Z5V6ALcbioL
J/YMJ3SfQk2P8rPv3eLbw59S6+OUHfPIJn8BEs1KzGrq40dcOGDD1Ck3mwCYc0ur
5IxmwTq5JQ2SQxZS07ndsynTndOkHbff8mxk3I7i+01x8ms4hdkueR5YCNmhDdi2
MUcNmy3ctUv2+F4qlzxgQilHxIorfJ2p5n0rmq3unEHvGlk3uP1LriCuGDxcYIiL
sF+8GB7XfRmEFVhHFw8jePcJIGLh0CNx2HYxtKWcJZeZqubC8irnHZl1uJutlncs
kc/UG59T6ddtBBIrgxzyQRvJ6WJ96XSdtwTEUMqRgkvI11JGbPWHlRWqFq1HTF64
M3yIccg2ptmQOIlsbilfM69fc7Fbznjg/ZW669o8h+8QNJ/OiAZm6upOAWvuMWTQ
imq2DFdrD2/DSPVM1MKnWQ1iwvWMjzvwDj7RAbA67EZrLJ3pf0v8D1h4lo0OV/kG
AYNmHdJJ6OLSM38R8FATpEICiPLjAVKDwTNDnf08zO8shOzPvJlo4W+xOFPcjFVN
m4wawv9fkDPSgSRmK2+OmGZ8WH6vqGMNTG4BTbGly9bIyU7I0VivkcZL0c+ImdUH
6sKsYR5kwpvMiBSO5Q6xPGQvTvpiAjoGqOIpwH+YlU5lZ/K7/UMsmmUTDEGglvm5
XYMca3YTHi034ORO+9b5ajSbRkuWyYpW0KafndsAaCjiQwCMgUMVYxGXon5sgIaN
bcrH3hOv6faHtxTYZVGjK4un+t3p9iOcihxg0l32Afw1qaUwLqPO6Ltfx2ZuRYIE
nnOYqZ45P9wUmBZDQxswO8i6d8U4u09+I6AaWEwKOHJETmPAvlEaBxU+vPHqpnQY
eER/AvepTSXoG0gT0enF+F3bN7AhwzwEbEAeXpQQE3Zsdlj7UaLcjKL6cdF9DwNc
AKIa4IWvZBUqUnDdNc17ka3v66gVhN1oracRxN52K7fLko4P09YV6fAk4p0+zKek
ctw7Y+BG4LYs/OIX/CRTFPjPGxET4bCQBGC2y7l5nNBXzclQPTyy4lyRQjTQfquT
bT9wi+zmj/mPFORQptOu6V3lr3xCCSQ+uKaM5iP7991RzetQKbfFCMyDJajDPsec
gFLXKDVgtt1jiiWK/d2uF/dCul93dh0Yz6dfToydEC6l91oHCvp+Yt+AUJH0vJ9R
ycXmx9/kNOwjNesAfwqg17pLrtxhcGP9ySImi9c05+/YP/2egBpboqkNrcPgFPZd
xTfkuPMDfgwLcocm0P1hLHXh+iOYdedSQeaI1AqEhP+7jBt11oI9kc3RdCjHw96j
XQCGTxxgCw+RwhyDT9OLxYI/auxsDJ536+aqhNtx/zRSAIRe//aWqW9eVJ0JZ9eR
3cG2E6q0PGUJY1aWjV1N79ua2SSawQFwzprqU17/QRTQ1Uf9K/jmVb5DY1LtJa1m
Z19s+gsNonT/C8Fveg+Flygy6VFtTtq3dP0Fr1T8SKvfRTV5TMgROkzcVAAmtQFi
G1wE26aLXBzTnAgIm8V24S6QKcptC8vjLy7TehH/i2OeYbNevrFAl/XVnidzbIsn
Mh6MQ63HQ9wi6/JeHBaTgGPLFiIkVKhuLA0JoxBYTp3FUPe07mTjhNWwFD7mYZbC
PssgrJgs/dU5TH+60F9iJDwwz7bHh/e4XKMwGj2dkTgjLfRAolgawt8N7fKwFDr2
Kxpiw2qF6hS+m5rlo7HSW0jO6u9Gy+qZHQmvi026rA3qJT7d52uD0cPyKRBJnobG
IbGgvr0oxdYKR+wr9ZtYBN6vBqu6RMkjixfpXhAqEmXAkHcYW7YX0bezjqvGir0S
2lbwa0fTmiWNT27ebF7/QYou370KW0fY9wyz1GRt0CZLxxHb+mFFr4Q0s+JP6r3q
8ZWNjCQGAtfk1vjOAb+7fyuQTMhj/hP6FaRiZSgv94++sHgCPRu+2IzSM8Eu1FM6
M5EBHP4veW01bhZxtHX3hu9k40WY0WWoo6FnA22US6+vdlSAOYEmVxoe7Duvu9lI
jyPrlTEj2FdVMpl5QVg/M9Y/1qkXR+8UNmQS3pNAoRCSklDMogVkiiJvbfYFH+us
2os657JIfUTAX46AuYV2zU4HzG5EDqb2uuX8TYOszbNZbX6IUqRcI9xIKH7RPhhs
V2EOcR1A0RwD38ORijjWGAbbLzKnQN6JaREUThS85g80Y+g3WCuRc6wx5vAM6HB9
P/epOuf/3JWGWoOFNWd8f/H6C4roluWlhrhIrb6p5qV53ShoZHuRKKk9ozFnBYRC
t1/jYSdxiRhkARxmJR298YAKH95OwTzFT51GpcTUwoXc/cLQHE4G6O0LmnXvsSCs
s6TaCdlkDX3beeY0rwpfEDQzVh29MugEsAVJCwlXsK3JvqWxC5C6eyFOX/UKsBKf
2kmZeYOBb+x+AS11aSSIHrWrt52aBw3+yFaoOGGAITcoF+x1tN257G4PE+KcS3lu
FHzDvtWchm2j6jMdtPnwTsn+35L8UMyoViq/gd75R3SbLQh45T+hCD/v7zXrbnRW
IEy/FsP9Dxuiy3GiUj8EtPeHLL29nMSzx25213NQMuDV86laJ/bfHMi9F1xZXF8/
f73j66U9xwzF0wR191Oa1QCtco3LD4bYIV1o5NmjxLf0PofiO/BWw1Az/SlDe8dL
PleafhEukpTKhvsepwacbCR8vBbvrDbrGSq3x8IeiBNks2Lyn+eXfGOP6xaSbOh3
15q2lJGfKjZa4+Ef0DY60D/Z9eHfQFl0Dk+s/GAbkb4Cx2hKLCgvqbqJNWxa6niQ
+garQG2om9f5SzJWnTYqsYLmkxPaMyIy1B3wJabHyCG6e0A5gOdciogg6AcKi6/X
YJsjOrgQ7bOPciNaVdlbG58zhWasstNyC8DnzJa2feg5ayKr25cD2o+g3DvXYyBQ
/3YNG3NyT5k6wtJkUqpIepdTAKFnez2cPRUYckV2BzwowLk44bzb06b2WCd7kTt/
sjxSGZXMJo6IAplo9ujYzIZ4VyInK2SPrYBnqpc+fIghs8c4nkAmr8ERjV3zGidt
fSuB/I6kt8Zj0wbFHSo+zHUi1/btyKMDuwvqAcv3eUZrQZFZMyyZ+m2CR3UgRb1k
xXKo9T1QxAIKCWTGSzfM8KnmpdYXHplfNXCsJahE1iVXD75kov6eyzkqCZPEv5R0
xi1OtYTT//TqS3umFbkuRof7uL5In7eS7Z/7LDHIVZpjS7UJbXxSzDQvJAyKJsoT
h4N6SIBQKInDcYsuRVulM6oz9R3WKX1AnrXXNFJOwGO+Fkz8xwpnh6Q9FQDglsEs
ATrXYCEJSSJPht0SxCFEzD+0bEL7bkuJ2FNnDz7RBsLIDkv+17YfuXXoc6NM9BYK
6Jt+hpGYHUXxsYJq/2lVGb/NShPmkIYguuv+8M3uGcMvEwBlIYNwwBtroncqWGPy
9QAb0Swzck0Xg5E3nL19/oZSOZrZX13aoqwihgs56gAsn+fqtu+c6qoANWq7zz79
CpUxk0g1dB4yYutESOQYa145GD92a3OuKUElSMscNrwskhldVd/hZnPK6I10OOPZ
W53OPOApQ9K4ao8vmjZky2oq2M+gCff7rWx/DrY1/SK9RLk9VqPqciQA1rFh5Rsf
Gx8GuFWOTi8FjbWlQndOJW/IyeCKVmHpe7LL+vimW2D6GtNJC+zShUrEH5qYlTkt
mXjR8AsYhcw7xBzfKoVOIPjmegOXjkEJoLZynO4Y+1+7oqI+Q+5KORcaTj2tgVyl
u0taF46lcU6UIll8wEKUGyqYiX7uJN+mkRu7or4rxi++XwKRrK3kzS46gGQS/Nwf
pgOd438W/mnD258cHhc7VDgefEUnjxiocTLeQOIIwbW/fGgOlCJSkGY+Jyqq7eLY
C7eHdfQ20ShYBWO5DTTQYVEYS6IhErS37OkbaG2jwt2ldYhveeGwcMvprntM56Cp
4hAhF65k7+7Xjk6WfSl1GeM1ocwMIaHEDnJhlkEvILsFN1uN2Ar9oqJrTtAWgOEf
z1pGI3VOGBox3iN6RoFQEUUjEmlUO0MhB1t+h6Qw+lRtRJlXzZosVKYNymWonWHb
jaH7LUS5Ysm+ugakaZmTSNAIXfN3OAZfGyz2VmhGfmG1tklXCWJtTt08lb6dUHmD
JreKJVguwiAMXKjnfB38jIZCX5ssGcSGBReeH7zMD+5nAQVQyA3LXwrAs0NtOgAV
v0ZGhi8KLAy9ob85GYbtUQvomESP/WM35Y6NHwI3d+I1HjasFCt7tuCGbWs+6mZC
QBYYdwqvpl3aJ94qQAxQgouzGZx7XirREV9sS7Z49pzT2n2++PoJwQkTQCWmmtZm
RlrOT8/SsJoiV4nSpdzmyebDjjVP7Cg7Fm1xi5hCvGv1/aVaLYZ/Gv0jZvsBrAfc
OH06p8FFOkjJPyNS/KXJ9wDqFTt5mde6iBciL0XSSkoBO1YeSIoIr/GdQoXsOIol
sqdcyZUC2O5HNY3IM/E6ADWxDdPAiUbEfMTHwqKCz4trBuvkm8osN0+4UjCZGu0T
OBtqPg+1rM/PUr42dI1uV/N+uiRibQjHHx+BDUBjrfmOtB6Y9TgoapqXc3dPJ7qn
Qw2397yRFArF7L6GYf8cSsYgQuwe9peKyqdqnPRmAs0EEiPUBUqB4RJQNGQwapak
2seLzWNy55G/mw8uzCTzWTyPmXBwS1xUa5x0Pse4n707FkDSO30k8H8c2ueQBA2p
PtIUcYSN0DJyIg+hxehehZQ5alqLCM0vbGBV7xXL5O+rB88Vpc9EDGXYv6BGTSbQ
HLh39jLKqc9Hzn196Cw16ssJUflre2y+VpD3y+A8Z5adgYoXl6BWLy+QjluyJPJp
afIzXe7eIT3t4KXXB+82lxCIchgZdCD0a4X7b0wTKZMFGQQ/kUZ7QUB043jP2b4A
+UUXFVJ52GfwWpDBZADRf+28EtAQZNp+wJ+uj0kU9cxnrTfNffjNjzlLrBv7TXhf
7YUR0Bi0swp8JYWDrMG6MgskwWjOR/WfWwDExEAjKILBVBuQQWPigjVJKeJFhWsg
oyovM9MgkbjMkHNuF0iZtOY3ZvYhVKu9O2d3m/bsuJEqePSK4j84QLXtdJNv8ndk
ZYXOKvwjIatofYjdr5kSIPcBiqRIUtq3wVGK8jfMQ5LoLxlPEC1+8dcH/j4XHUKv
0sgJnMebi23QLAR0tepobnlLVDx3LLduUNb2Y9Oz4HFWlEdZThkdlEtFZ7c+Y1/V
eTBDKBIPp+AsiUmSue5JtCEeSEUbcmbykY8qDJp+xVq/CaOvnrLF42m9H77BDGOL
mF5jO1w9GpVB0uWcxzmBymQaUHVyOPK2JV3pKQ9pDfLGlN71I8XeEgznVkX0jNyJ
m3Y/USWBgoWMHuMEnE3LgwjyJx9ron9+QwLvhTTjQO3ZGk7yxO87KnV/phwrBZFr
SF7GqT+nhvBjMrqWF+ue6mkVg3Y5fG6QrZg2jqQmXWdutgMizbRpCOeyqm31Aejf
s14wBqW19RhvUFjPD6a/Z1OhuRc5gcz0qeTAgi/PvaLPrWmW+HyoXifOhL30K7oU
syN04rqTDlAYwHMkuefpoPDO4KGc64+a8zV3XKLuLqeOY5Y82FM8xKP3xlgJ7QRW
30mDMF+pXCCMEhlXMuOzPCXs67tklWp2UWYQw9rVJjmxGrsFH8X3tI6o+DofrBmc
Qc9Laq3NXcsScAfL0R4zqmOco5Eqe1jEXGwf/uinJr4NSjnoEDNASdBWg8u0WpFW
ZMfWXqR9G2MT/4poIXImLnX6p1XzHCHXHCFfEDenAmYJvV2EDn7StMSF10Qf7/lc
tuZpfwXU8XV85u8FBvoszLnaJcOQZxDezNqGzVU0wt2xqoLVaOHVnWDVwOk2allf
gv9Hizo+95UjcDoxBLLAuBu/RseF5l0KLRW7ECRtTDZdq1M8DzxK4sPj8d+RKR4R
8py79szA5FUCJRD2X+zXsg5lcSKOzA0mmNaS5ns/9iFYlBDNYuB42ibfGe9LJeDr
64rmt52hJKq+vV+BeSf2gg631JFl5JmerrmKJFsVeEoNHHbyqxddU0hetsZ24Pz6
lR6xgANe1RbgbBPJIDSzq9vOBThuevqIi8v71BxuqObvzVoeg2347nePVD2ZvdV3
LJ64id0JitaE9QSwApYpKnzfGV4idkNGYdzFzimQbHCr6KHkMtDDqKLNQkwjUO6/
mkMMRuJ2W8yt8F3AusMC1kgT8L57s4w76NEe0o083dzaF5kZNC8Z7u08G4WPcZfA
jjLBBsOrEcBUt4IlfFRkK95kqnvjqJBzeWf8bse7NU8Kw3KvrA7hr1kiGz88rjKw
wWmhXlftsN/cUWeb1CDOcn8H3PptWGiwDSZxQ3xSoHygKKPiNQjUh/NpsjSGV/Ad
MHNYBZf1onH84z9tIBc4DQXvnjvvfvcWbX0a8YDU7fmYuaB6vO23Fg1B1nxnKYhi
MJnF4T9o0nDIHBX6b3rPc9a4gAXRDLe4NmtJAEYkw/HoYpNAh1Gng41eWEieEN2m
pNLZFNTN22Gf66sHEYCmywI5EAA9D/ModW+1W/Hh+ROpOmYAK+0B/ZSFp5KdbR8h
icfmeegcRsVErq4XY8oXHagGfofrDfz8R6PGS0Z2+TWuMBCUGM+Oxvw3aTsUZb9m
m0pvILkpXdKwxnoZwm9J9bb7DLtfPWWF5nKO6kzzUlXOWThoLgQ7tdwFAsfZdGgg
ZZyTMXsDSl7XVOBf5fVBQN6dqh0KZL7mhk3/y0o40UhPIDiW7ji1Pgp/mTflNGNI
Yr7tRdTtiAFhBA4+PMU6SDcVOq/dSDpElC2wpFdmxxaeIfxEcUTVJ/AvrnYaXa1U
VKui+oL5qIe+XSfqUVJAi3j42nq6FwQHAOOaIZhahvf+gS9zYiWj8gOjydmyMic5
2yWR8fVsjWtL3mm1HxhZulrKrYofTfvSfuGytlo+QEsS6R88ar2WaSh43lz4Q3Ez
Jp3WHnGivS5hmd453ssil6IuDhVDcSmpI0j7NR2ataStr5r8OQ5UA77Kso/jdhQn
fN+nLAmkl7fWyfwF0fvLkpatGtHWtCQFwlLYBefMY6QtIRQscIlUIJu2WK5wKb5L
Rgujr/tNrqy3DxDYYj/7uHozhITsYe2RVPjWhlkZcfWdJt2/H7WYquM6cC1z+8Uy
XuHmq6iMiA3Lu1F1FJIRE2aW9Wb2ZRGAGJ0xAYIMrf/71NtFPcgpgfDn4vHmZ4fd
gTHWMqAR1Sqwh0+GOv9Oeb/LlKZUIXTUKSmvKCGLaDEhdApE72IBrhuSdWaPcbY5
gEqdbHXoDwslnKx5tM3dp+cHNcK3PjODVN0EFRkY56p40Hzf7y/zkAA1+h9qr3E8
HP8RO1yYO3wFDSow7eAKtD4MVviQ42hZfJ5k1ODFMw5BIEVGNYmngk9NE3UT5++n
aUU6M4n4hZuq0IxjrxUmv4f3S/wb/YwX0WH/lPs6zQ1ZIG4BUIhQkaka65IDd+Uk
35bsglk6Z6TxGZ5oLLND+Nx1L2eC7GuW6nQrY6Tmyq9AWqH1nBvtUJiMwt9gKJcR
leeoejk64T43D/bcj9oT1DwDOqX//5gJGv97/hCo/aX5+NTAXIqzu+2wyfRsYZbA
xdJKPUPcixVWJNWdixlX//XxHjUOUq5PUiYdBathTpCG1FAmKQohsuH+W1TaCEPv
eFzcNR+RBhRv0/eebJ2zA+FYRgfZkONTstLqwA/ruKpPQArobLyG05kE4C/XgZEj
3IimaLLaLl/FiLuBjLPmoDo6TMSPn5NzZpYdBmp0FQXqXYRA+0ND8aVF8WTt0gjg
jHgWMzEHHW3Drdl5LNVyBqQLY3OGSsyQ0Or3xR2df0wx/HEG/QPo63xvV6G7k9yk
KykuWBUDbA6kuYQyxZAcFoXAHvE3Bcq9JwdH74hzMumx0cX7MY0oB0RdBFpnpTor
wGNaQ8yzBnorl4A8scfwKgF/BqqxBuuR8miTA0bu9R1X/0GMx78iE3yQ28/cxiT6
w1WxRk7EIvdxYA4ExLN5kZECdtwCfdeQpQEKzQtLOKN9mwITPNjiK1lFEoN0r5tq
MG1Tyf4yGxF9+W02zZBDrkiHWVY40d3Rs73f6i2oYWR5YAq9X7jCrWKQ6Vh8okB8
tXE1qIPH4FeOBLdd76tSfWu5ojHDMQcXnui6+HMKNWTQlN+aC3aEfCzv/B5hezym
rncXpa67srD17YEc2qE6Xh8xcPxyUS38Ugo8w5Y0vrn643zn3F+Vm3RoPg4hMgfl
mapmYwgNrBJa/41/6nfMV4CZ1YZhiKFcR/iqW6X+FsJJazfHeXhz6R3esfuL6xvy
XwQspwUxVMMNCXhjWPA/aEoynJf2C71/vCpcNUs39X6pYlgRfiQG/CeUJq5sakmr
y22xvKzBFNumkA93JkPGkp7wMrExyI3729fB3LY+3euM5RJFCRFLaK/B2bDMSAJm
6DPRiGYO287v8Bh7N0SX1A==
`protect end_protected