`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 9600 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/9huKRhRMtvnNqb3Z+UU7TahEoHV+T8U3P3ufru7l1O
3DlgtZzb9QxCbOjthp9+wDkjygH0eUfDrEl1ovhZG617qdJ+qf1NnRVd3F5Vjp4N
Oc8v4VwIOg+zcFZLk9TG27fjKkVbz5gELvynB0tY6gywds8EltZ9UdXPSZYt2ZGP
YqwQ4c9XMjUwNnyaenIS5kPCgzRrOPk/JXrwp7B+cb02+iJSaT7pGTX5V+IsFrmd
pGQpH1Lq1LjhTNksoyRITCxYyvKLE5cn4e037wq4R4+nexc5Nu8MV778A4zSyHww
jSqW+ahm871pVHSwQvCk3ZPIVMWPQuhFfSVunLOSmXcbwUnNnVHmSgP5LJmolKvm
oJth1gjOToeRKLo+k4RzGX8zqgcvPF8JQWWHl2ruvdo5I9Wj9gr4IJG82hSqjp4m
qmoXI/BfLDVyXN/9b7PCnQ+GoqauC5R5KC0mCXIm0MX+3gdLI8MLlahDxOQDAr3h
ocl4R/zxs8xt2XwiUfiRPYyBF+5/QR5VwY1pOVZSiOM4NZDtItTFMtPNaEP6/Ub1
D+rVF0nECYO3JHmkfjabeOaQWSfSsU75iYwvA+RXr/fD8dMd8Nw7Ws7mBr6whIkC
qdUu9321aKokvkCzwnyTJxNut6WObDsJWSJ+M/fR25DggdUpAuSPtupLrVfftS/G
YypNzSB+kSNlxahSqVaGDmQHoftPK0SaL9l+ZvvQwc0lStiDvVqVso+CfyiRN24l
vdVlfov8icbxEqomIXS4M2Z57mxcRWRx7dJx+i5Rtjfyg6dY8EuV/rmN1SisDDDl
1D/ekwX+VWIVlSX9mfU1asDsiZN/8iE6imfJXDiYP4KWyNcZoNReNsu9RbGt9vnx
6C9SdZM0dPQdksG08ivCh4ttNe8eigOPTQDL+0aHv8uojIcUqUwtYMPp90F7fCmQ
K5uCkb7zZbZr73q2Pj61MxQAtsBjfCdWRJa5VaWksTY/YJuyQy/8tDZIBYqohCv2
7CitaCYdVdp7xwempbSjhtmUSxSlGuDk59kbOXOTGbnHzQmxagXRNVUAVTTzF3Rz
g+ZDw/qWq/2yCKUYSdFe7iPADv5PVuPxhhuJ+D9Qqx517tf3Qg7fPHdQBdfWqCrX
4vyOoyhlygzT4nVVq5d5CWu66W8uXuhwTlNLrI7+oEFwo35BGFtuccCQEKjoREOJ
runUtSSfPqK63cfRkE8RKtR5uEkArkQLhfkHScW6OIfRhKWoSpHZZbO9Uj7rq9C6
xAOdgpcBgALdzcROqdUVIvA3L/U2VDwwbwXhLzJfnKVOmZu/ez+y/5DcaR4TmFYk
NMS95VMcTErpkZmc+PfhBOnRZAayGKyxe15lfiB9tPDGRhxaWiCv/S/Cvbbiy7al
+Bz4qm1HKXArkYybtCevZEHJQKhK3mx8vnVCI/ppPeu4uH3opXiiBW4FsS3ka06d
MkxDwwrIC76B4L61yRJAFgkqetoa2jPBbcsB+Sh1wQZfLOsM8kQiIxAfoMfoR8PY
AQ/TwSeZ/EK9fr06KmxDIKxaG9/DZEoScpvQWRXYYz9cXDr3F5OW0uT3svqIiQ+C
19DSGRX+C/mbdWgJiTmY5fnSXJ4UAT2QL5u1cgX7rB8K3wsdNK4X5IkCpz7kzkgA
PQzyY+eNp7aKeJ8N2fhZSFIJCHe/v67pDniraEvz1z6c1vCLZOdTJRlRs0u8KW6c
IijeTQkYE6ki7HEKEE4RWlqFCjzjNuFanWVnD1Nh5nD/cdrxhVGFXQ0iGzDM4rtY
lfRTUfueqs/JARb3t3LPrF3HmxPeUSxEoL06b/rpgGfLyEokBWPn8McZ2iaeDnAi
MdP6DSsuAKARF7GY6oVqerKCRz1Z+w7qWD4LbXTbCEbo+U6dXDkD6dYvtr8szb/H
+FjD8GN5vNSD2mWr4dhAj2FmfOKgWUHz8CFE8N+RYHXLYIVnrvrX+paVZOhXa1+u
9vdR8Rf2sQ8gmOxrgsGDwy6QH+61pkwjXHhoHOXwiLLyYpXs7t4Sl4GwL0i+QDS0
8DO/6lxa0dToTB51+Ci4R49oG5kReBmTykaoh3Jh6NHYDvbfY2dvTLTQ4slLMgxb
NREzPG0dp9CcOlviMRKG8SU50t2nhEG/2Rffcht3Xv+EpyP1ZAIF9EkF1PILgZPe
cYSiQ9iAy+rg+JMznlIYdpIlGtryZ2ghyWPfHjVkDj//8IW8kTpLCC+HYrz2YZcR
CuRdwitmnXj0qI4xEIEyI4K1MOIKwfgngvI1yvUTvA8jvYzFpqEfEn+fCoYzWt1I
myEUC4aL2DLgEJUqE3w4DPcTTVVINd7JTq2OS3J8CjwFPAlh1QGcKPDdwfFCgPdq
4WD4guJhBcqvmVbUDNIGfUGtEWJmqd273v8b4zoqgtmlnhSvFIm9tb1QTzG7uiJ0
e6bqJn+YdUCG1s5aaqmeBBK9n1MMNP3HRJ7zGcQlXPmBILBEnOlQAL/DbIYhzkB/
LvrfwJAGBiC6pTGIhV6WBNMk4I/EyEFLCWAaONtwhQruezmTIG/LiauTrks/KQaL
tx026sMf3QW+ufCHvSGleZ/3fDEml2etYM0p51b/xrO0I38SM3jMFCGuBVv9LQTC
b06VoecFmIwcZ8Abi1Pn2mnPV/Od8sAT8alMDc4lH3Wv5QR3bcT/g+d04/fuJlpk
mnRr/D8CsAALSMyI5HpHbuzWMYkNutf3j+1AJFTew9gUKHpkvB0EfUg6cOaqMi/C
462zn0mAkcg9f2CICsm9RG1MlyJlW6+Y7eTqW0ThdC64kfMHitbYzUH9D33zdjbn
N1AzUi1ElH/9cvxRBEeU3p2IZNhTHr2dBZsGIU8/pJxfwlkfi/QNLrQyk6w6QrW+
5QkTZOR1EG6Br/xYi/J6gFEdd/0rCVyhXTdD3aobEdFaQV07G5kcaN/Z4ggPpUdl
xLen1vF4a+Vj9504/cbmIk/jYI9vRr+jhmVWkU2zFXubYkvkZ6DalYHfbB8MJ9Uu
nlObiS/o/h5j66el4kFnCIVw6PCDS5GVgAA6E9QyefJOwp4E/xHA7HVooenHezUc
qpo1vHoCAR+GSgg8TN2nrFEKr/L/zzckmf5u3N1+BzuMjF0YFpN1f7j9WK6wfLST
TbZ3M9aTI1cTjrCflb1hsHvwU0bO0d+9QF4t5ZjkgzeW/HqA5N6AoEKcM72dA58b
k8THo7N+ovtSbWQksgTJ2j4V8tETre/06fNunPsDj1kqoioUYYNeGOWg7CEeEUpv
8Kh/XnfSRMaLNNkMjMKgJeo6GWHWuY8WLg+3VK34Zy9Q/BLonNI9eAitZAXb8/Yl
CP+57mwlVQeceLb6WN0QvODnDKYXPN8B4CxbVHhI1xPPIyqjzxabKydlqkUMeicJ
Lzl8kyeeqg6tAHL9vSRmPEBLVhijmAZkmVowiYftEge+Fxzc0NU9lsVl2tnxOHFG
LwQsdgTkxO71UucJT9XSzFSQh1rSMJNnffsVb3z9waYcsckSEOjaZU1iW6PtBlc8
wH2klzPMreqiwDucUlxx1xLrgkJo/inCey0KQpuMHo+wlXGkLMI1C7Zkcx6lCsKn
PILcDbgNYwc9/yG9HG4TYjc77nHAM0UJH2xmG2tHO21xq7V867ioKITQJztZ2bqF
/kiRmpcfU25p1JlVDAEK4cGd+B+mkX2SNvGYMlvPSrHaMngch79MCNVvspQpPRL+
OHtuz+Q0Q86fmLrzpmw3iDR+8h8ws7L196WFEKNLbNGbEtbOpLA+UM6ncrXGb2hb
hE6jIA+zYq+8dquQ4VBLDHj8Lv07L8IHL81ggD/gXbSEhDnG2OZtbg7UPm5Iv5oA
I9Rgf8E4Y+JgbvehpLyNzZuBAQLXwBzPjFdCw/6tbiz99JSj0tErduWo/Uoyi59x
8XS+YAly5GpNo1V/mwX+Dk/WTEGKmwrygOIV5QV8HpFVx4pGR772QrOIRcCWhmPd
Nd80Gt25V21UKlxzs1wxqlTSeBsFpu79fA4DRQ235Z9+MwNQqtt1cyD5ySj1y4+7
S0jWSmngLINpQoERE+n1pEyG7kYUD+CNl+t11uH7Ie1n5Msc8vftu0qsBsfNgvcS
ZmI6tN93As6jYmPDFxbCAdvwctrgOfH0GLUTouqoyGJJH8DiIn+CPKUdYLAuPWCH
TQ10OjPPDY2/A2fbw7cgtvMPIty7E7KyvVN5ZlU1OWhYYpIRXvHTpT9IcRLecYWV
D4dbLkR7VQf+rxs2SNUG5K8e/pFLcZ7jQMxaSTGKW7uU9oI2P49eZasp7Lk38GQQ
5uViCpVSrbKwrj4mfAjlUOH4NryNG0j5mZQv9TVYWe8tANaxL5qwbebXW7spyqTt
zYNTZgLAwI1YloQHZNuA0m3pau6KeyFOV/VhNo5PGjw2GCxy6XZNxdOGhbsBf6B3
1bMC8I8E3iM1IXwUEwnayLOtXp5pD4ZMTm13GN4feCBlu7pKe9qWAsq2OCNl5Nzo
VtxciCTErULSik6irBpsf4rL4Ys38MIxftiBvvqM6g1v+61tlMREbWCc5eyosNhv
RQ1rUKmdEQPyz7V02WdjNiMGn3y8l/znhP9hQmZe+hONBicnst+Zjl5mEzBn/zbZ
/Bu9F3uoakuu6+IVhe/dn7Jp0GSabSkmO0WbJ9DtN3ZqAemAAHGkxmTvu6USnXi7
mgOf9u+GUJt0DcoSicqA85MVKaUlpW+KdQIZHKrszH+VcVgchWss5zfY6lm4mJqJ
WspTfc9wqkf+qRoR0MATsyDufqF+L2q6pmmUxoHoLff3WOfRCtfu9CEfWziFZCgj
g3sUSZmGVxv0b62B/W9t3mubLghxN5azB1krTdYpoT0RiVZfATpf91jxem2CHK1d
R5nF06XlrzK4kmJ/umlDVGd7qdkbFdtpO2mCWH31ZKOrqcm8Q6xqrarsaz/AjxPn
ouBmhxLpkCH6nY7kl+T937egm1cemnav4HE/XcBBenOQgFp9fD3T3+MBKkSlfszQ
Fp0WdSIeImTSc0ja49FW3Pm8Kvo57PMhFEwkQS7afLZhfVnvkcEhtYhb735oe5vE
VJc53a5Lf979PqTJ/T8ZQGDFBsZ4BEDUOyNHDuPI06ty7ZIL7glscAgTvD4UHRzn
s4mzgt4ESASCmOKmn/iISjDqvELB9aPLqDkQkJ7zRbzIUMfMjpxPFvRyv1c8ooAA
YxjQU/Qa66IFPC0i3uge7zwkivFYN8R4XywN4/o3S8MhY9JDSP2aQOnAOMYMW/ao
nN7y3CyHHIJfFujchMdZc1Eoek38nIsD47LW2nVVqTR/+RpiMtCX/3tmoX0LjbEQ
aiIgy0FvPjrurHtHf0qaXi7wMB1A7ZMCuFkoG05jEdlsZMu52qhXMWYi88qTiGAr
5xAAn3LGQkozcvAOPvTbVOQ2+P8l9UPjVxmVCoFiuD1EtjmsaJ5u540fD8xc1A39
Re9IUPouBrFbtWDFV3X6+hrlTuTrwRCF69EDJxlVjDUALxQ9DW4DL0MxJ579pJAB
vIZYGirZ8iY4/g6Tkuoz00JStYTuZZfCLl+zYKHGKYQDkVkqH/wBsHsFkP/79vel
qowXVpOwoMhxIKviC0EWmhRm6wp6++OyTrDScMOqCyIX3NNY0sf6ePEN6wnRVr8y
z5/A+gWwG+TvgWE8JJW0XhPAwB5SyzOYXasFODWOa8suyhPrcl8sOLHFh99QnpE+
7izFWxtF0Sx48qHYTCkj7s9cGja88sUGIeEBU/VfTv68FCHinpTU53ipv6tqeaQl
jj/mOOdJ6drdJLBMgZClxYpeV5/+JfrEu/3+nBdQTJ/p7o6DFpEQsZZiExVztcd/
7QHux3eX16nFbU6q0uw4NEyAdwQKvtnSs5Z2jW8oVHh9nG3K51Qh+W7FdVzhT9Fq
FgTezg8f5yn0CKvxhpebunLYADhaFK+DZrUXOKyp+Wwiw5n2tBeY25X1KUnFHic/
r80PmUQe5ItTRI/QRqpyEhq8xWQH4z4Re+r2HSceoUsQP99x2MgK0YZhY7Ki3Vbd
P0C1toxpJgZgLpWt+lFYpun2b6jAnHfkWfMjhwzXg5J/cpPMcb8g9sweILzMsr47
+QcoqKPD1ipHLlGN5pxCDAC20SDmf3EbqEAKKs0DnxvQfhkO/nWn+VvGtX5HRl2y
xkv6BVIFmwfr1/kR7it8jZ1PuCguNdG3c73BHQGKrjM2ItBUhH1PzC9mR+V0XKJL
liZFLsmF8asnCOZ0D5owsMiV2czxY/t9FNm37JQEVMTxbDQm+zm+RfV6qYjZ3TsO
5+lPN4IqwKKC9qy8yyC5wE5aOIHZJOR0wEwwvpLdZv5/ValKHag3i9bRUEUZzR9u
MScyLqDDSSYSO0i/KoLm27TrIjg5tSPytzV6LxFif2CWHDnCCpB94Ogdg+WitBI1
ENRGejhTQcim171d/kAZD+iqgRYfMdim9ZN1nl4gK9885kWZYU9Hn3S2ljI+CMGL
3h3fyG0Lv2T5ksPDj3dOJCtBkMKr7kRPCRc0WHUf8dBfuGs5qZZgGiutUayCkPGK
mgNYJpe1lv2K5eslVLXlyIiuHMjO/rVqdHc7kv8+1COFG1nZ+DXElOdCP6HV1qfv
kA1tFUJBTIt+wlXwtLRitxxNhrSX+dCHDyuqx3BPm0lhOcxffWoEOD8UXlrf0rpZ
M3ozUfmKQH6TCz7UIC3qmXfeYJmIdDTnbFlvdqUOn4fjLHOtBm2b5fbFZl6aEg/1
JKl15tgz5ihJ6OSY40Mt84/wQmAGW2wEb2sDhs6MR/NF3dN4dqgnxiXUsefVQ1J0
OajDfJnfKMjNiugSLUx2z/h67dseyjd8gYE3m65OkOQ4xk2wIeB1Ge0PfKy+AslD
f3T2T/FlADi42bb90+j+XNeYVSrTwe0hWRrey0wJWgBGlndEd/sTX/hchxr09wZ/
Qz27GXhlZcFjnKWjfWFX8kh2JKbhIXHpnwX8ZfczWzRcyxvZy5EGqkmlM4QAvVIg
tMVWQNSvysrKV9EBU0u4o4lsJzRXJkzaDYCV6xA0QOl1fLGcH3XAonz3XoZAx8Xm
j5B4ct5qm/Jk/8ZUj2jpE5OuP5FpfqLCwtF0K85L6wNFKv9NPqav8YfS1pAnjGcI
OWWAiBLZGAybKljJAcM7XLEB9IeK7pR3Eh1SSaI5sNH9PbyH5+lcMpbyaaSrcqxr
s2G/CiPixz0ssYzlCsjz246Wmv+mnOgUE6iOjKTj9EW8JKfGWPlwf0m+sIQuoCcb
SnP6GXHHATWuxsP05QO18ZBO4MaSptnbCzLU0Sb6Q0YXu+s6hVHwTYn+ULgWT3/O
MKniRjOR0idItG4iC2/VWnAx4Nc64qp6AgDgokJJvVW8EVqpx8qP0nX6OWgcCA6c
Wb0aN0MRIRlLtZbsFKmtEqFaPnY4qzrAPvyoAikWhxO4JIS+yeBBaOhtcnIZTtoI
k959aFZ7c0au9Mij0h2B7q1AuftvID6untjvoxg/AUGpwl99gn9fXyy7hOha3LTa
P+m/lYm13vwkfHXCAOYZjKOBSPWRPwIML21zf9onBd3xvGr0dL4HQ1S35RJnyvLE
i4UzawQZvIMtzS4FcdwEw4GbyO/aPQJdQdke+Edd8QafS8FNN1r0OAFkyTEwYUgH
wBIV9DF788paqHH13E21ya39W69saa5L43dFymsd+++ZJzShAf6pQyN0Zc3dnnI3
UYkzzcLuTpOBIlLkTEVv+OKlnQJWYp1FJoIcI2u6MWXoWxl2nYR5soWkNxCCFGWv
VLbQV2U023bv1l14/Y00TMzlNOIWFTNjWyVAZxwF9fp94HQganOmukDZiCGLZLYb
Lmw0GRO/2QJsX17vD49uXsAsg20F/HgC6OrX408WqR64IuveII1uj2uKqnGuX1sM
0yDfECN405iPNP4AVDTHK+Tj5kbBs+VMGJ/HfUGHHUzWpnqY/qGRtdCZ00zpnePY
ScBccJrChYR6Xw+Ye20wu6g12YNr2xOLQsMuhxwLHYvsSe2rV0MIXF7RfDz9Q1jP
+qxz3r78oT7T/XuD2Zxeg6oRFSeqFRuJGtTCv6Du/uXm6Z3K+V6RZWoHk2f8zFcn
mseTaStXJD2NuxfBQH4VyhS2UIljlCd3YhEOq38rvQl96gJlMIduiM5jpTGcL7P8
RCS1zCJXj54qEC768C2QmBP4VqitDpnoU2abTcSTVx6/UcAA78V9xIgdXMpKpl+0
firyC2NPekaVYRusrEs0fzp/KeI/Tj+bm0gBpvCqCfMzTYkjgVKbTrRwxgp1h93F
6CAhtzKfFjLPwwP7rBlt6KF112kNl3XJc1gv3YILtfN6RwoInNZLf0W/wvGS3gf2
WvyCjPpHq51x/ewkEOuew/kqeIx7lTZjqJVJ144OYKi9z94r9KCi9ZiKo4TYDniA
TxT0/4TlbqUEIA3gvdC1OIUkQ6pXiJhtSJFLNEFZf+IDyYIp2fiXqO//zBduUFwJ
caI0Gl4OTNYNPxCWoorEEESMpjE0HMtNZuIe6a1476cuy1IgaODwXTYmMVZefE9A
iyo3fmdvqC9iVUxTCNM30lSvOzhdYmnnXT9HTCmvvoDENPj9U6L96kJajRIRjbNV
NeCbNyDHqUiYgaBWYldlFin3Zqer+0Ua4Sh+lZXWxPM26/DWjt8KZsHhEcqmV84Y
6KAr7X+s6MP7jLy6gIQ3s79k5OHj7ty6CH5oYVKBElmAgMxeWjCVt5GaRhSMs/Qj
qOGy/jnZm11+a+zTpA4zfE9Fob86FM2Ids2DAhY1autuE3OwIif9fjzmGLoOLNUO
kK+4S632fhrN+fMa/3h2DGNKff2kLuRveBrobMJ6Nhy+n+EwOT/a6SYl3AUKfkA2
mj4D1IJg6ahLsDnI80L4sBm0IvtBBjGNuGkIW7D82mNpjCaY5Yj9oq3eqaVWviIH
mxR0hlzzeFCBowdS/LXcJFB4A7Hh7EFbMj2oPCHQ795ntTJaR3cJ6bbYHZO8ydJi
opUbXAE7ezBfnZie4LaqKs1VDzQ3Egh3zW/W9NIR+ZY06edsIXiWTuKeg/X5FxMa
Kua1ZR7P4oho76yKHjJ+LZtNVIrtGEGVtFXA3RttRgvxt7Sfpt4wj2ST1Tiybkzx
LYW6POLGkUSA+YLVeZvD+AfdEUyArBkq74mN397kw5LcRpR5e3cNDlis9L94veYI
jhj+8fob5zf1pGH1cjRQVT6Bm7PexBKTneN7ZKxIibD0cxE+M53FYKi0S8JQKFJb
nJNcthfeBzfwsmzYmVrgougcnnlbRHv65y2KF0ErRsLKYqIeuLqB7MTd1+xW5QwT
mj7jNExcF/F76R58LSJK1pR1xRsPequXRFVY9voybF/gVev7/CVdrcNmW/838X3l
EzHDpXmiWi6l3Oz3vhH3245fDcKc3YqRoWkiZF1Go7flD8clRqm1z0jhFMbI5/EK
ecv09d8+bmvHJ2vhTqsrffsaEhP8ctoC31LEn0rZdJEzkX4d02j5MASbzUbBjpaO
x1twEz+4qVskK2pkN3Z0D3Gi7WTf761Rky3A3uka4PZp2l/CmsarTWaxQATCPMP2
RAvEI+zxhC6qXyPX3gPzYvdzGOnmqitYdo5icUxrECBl3PrJFgNlUOyLnI9+s+e7
rv42fTlaRympqnPcmaXrOns9U4B/s5ffJAwk3ijDaGAGEf+eqpNgsf/RZ55GhCal
oxXRC4EDDFQiZxx+voAw0Oo4M+XpftXfN6Q/SBeYDtP3H8Hv1PIVjITACoxb4fQJ
PugX4zc6hoD0zEkLqWib580VpiDpi6DDpFr+PXZdoBRewP5EubCdyA0mSNMk7q0Y
5ramNfgKI/U+Ou/RXf05yg2r26W1HKSpZY+L2oV6tZj7KvAw++1ULDCahGXoaE4t
fObeUzQHLyAzmWMbQYbmUADF4N31cKZv9SrebEcRKqpLfy3933vzeeZ0zyQzPCvz
5vkArgg0/0z2qCoxsgIYhnp70jcwkDB/qvVO1Tj2pJBWqve7a1SrqSpCb2bJ8iNq
31/itdimvS+ye0YfkropZs1zgW1cXEYZjZGMJ8M6mNcDC+IubiATaioHTnw5ZNEc
gTat917WK1nTmPZosMeRCeVV1pdhHFC62LkxqHqmbX0WwM++B8KzmDsnvyOJX/Z8
6Z75/m33j0N7WhSTRXF5sGJ2okYbGl+jORmsOwNvmJt8LOIGlKMirbJB5uGLzp3K
UDKqOLQzCFR3Qn+ASxJvwJ1QzQJbvcYfp7BFRH6N7AZir46sxqWphERAaPy7htmR
/DTK1YDKnbQKFOZO/E61DRt11zIlFqYlkXGYTtxzG6QxGdChHwrOH/NbuURtUF3d
Ko++HKdsNIVB03E3pj6OJtaT9Wk6UNJlP1o5NFWJc+OfvHzUVvXSVqd13vL/MAxQ
eC+lRGhqXV7aoj+obwuMWYw0GCMR3vsnHk9v+zwu3BZtwpSAv8GgX6KXIHompjDa
Mb70E1tK1BSXvEzKIyvqnKUbWU3pMvhu8GkzdukMFLkaxOSuvBx4mBfTmmxFC8oY
YqTVO/GpGKU4At7HQTlESSWjAxejOF31FA0hDBuPh7Y1i9ojCjslF2sX0dPptX5w
/+EPasn62zdZFWcR8wp00e1p9WEjK8H9b6sn/o9iU3SVIC99+AYLG6FfdkGVO0vi
Q8n2jZ0kgMIQ2f8w6al+/dZ5CpJN7MoISXRCeExdyqSnHwxF1g3siKlKMJHsjM2u
IgAXPMZ3VpWe1ZrzQwjHOkM1V7gYEb3RNRUbMgS2gffLUHwuWTzTdyvhySw27jAX
JuSVInvLniAZgumNIFbXUFXry7NYjOwg0EpJSZCVO5/azZKP73aeb9eO/yBFXhHR
9yuY1cAXIM5agnQzFFDGhtMp39vOxDh0K1zbO3WB29Lj/APaHnTDqYqNA+YBn/G/
Z0Wr2UUWMHTQSowM+N1Af41vzH32GS0T/FQmzOIp9FggkQTSRgjtgrvMUVnGi9Vt
9AKU5NWQmcDa6e6kwZKfeoCOMRJVDBluyCXWxJHH6Zg2VdbcPyh6I78wVNzPMrbK
DGcylJFp6XJkavTwT7pfjz1QqA7BPIlK3LgFrFF4xj/y/0ymBqXzz2ah1kA0Z6GP
R8ae2NjkkB9F7uJN3Sy2oE1LaByAGsXFaV8SzJfdMi+tdH9PIaN6o5uuqxqHC8kT
i+H0wtllWTBQ4U8PbYrSfJ0HF7rn+qZeacSZ+MSRmh5O31Nrty18mGKts5eALyb7
Axwjz57VY4cwD6fSlyL8Lx5/l96b7ZH/ppDiwgOIVUt6O2y2kTAIMPO9EqvvYyqK
yTyf04UpcxcQMFPPmY7JemsyAANYMtLDvPEe9l7MaHdIUJ3nz+mzIXfgymRvNGSk
r2B8Hi1trb96h26v9bzOHkoruUoWxORmkLxcYuPYtXcGsCJtMXjpuJEQVzrEA3v9
JdreazVfWWvwXjZQeUG3TmkjAOJfQVIfM9uUVJfHYqU0sTdI2L/YvlYTyiDkLRFh
2Zp8v5+cex0QKkanKHtH2xgqJraBPBuMhrAwzDblRdrZv0qRBzQ0k7FWPSUcc7Yv
WCHHUIGclBN9lmhsBxhLnCvbMvdWEOHJFIC5v9ARlUz+gWt9tEzFr6bgjUGe1oJu
uYp/4nJc+1qTScn8rflDLoP+18DCdZod2ZEjVfZhlYILatqmRkpVM6pBfZX8Enis
v+V97Y4UOvCvRwLeZZ6fqok8L1XweRxLdYCaI2GEAP8nOmMu3zF879M1RoUC90fu
2zCdfwXWcTwVGbcIiW5KXlmH1e11uXxMlH4Y/GgK6wwohYXIZzzbXXLK13P32SRv
kKLMq6lc9ZrgmqChLXdtSsqYEP9IF4Qj0J28q2uUPBLMypJoWmfPWG2zPHAxzYwF
ahMwV5+/MjAFu03A7+BBMmm8P/IiPa6qCgq6utb+r65N7sk1kx1hv7aewurzLxAN
+VK7uDXhfnvf0owEhqHX078wVh/2xNl4VyeMas0fCpN2KSHsJf3AO4s4DQjRqxDl
wgkP9Qlu0sqCVpgY0fYRiqbcgUYCIhmpQyNTArHpmVkmyAEBbYLkzEstpSPb0/4/
DzQdNn3hOvluug6qOxStg9m8HO9S9oiseDeek4JRDJCHWCJcKQaK/O5gF8QwmUxR
/wPPRTYQprRjhPKxkLUvDYyza7OI0RqMn2Om0B3zeC3yhmQPOy732N2tc2Pp6c7C
w4SFow9Um6y9B+h/VAMOnGBth6I8T2b+8yPJRR+f5lqahXzGk0vsk7IDS0UjTb0V
F2objBQxFAfEuygj9H6CygEb+uYli+HKXl4bP6ICCYj0UNjYSdyYjaqD93mY3DXJ
7+H3q274iDKrQmJ4qq6b+nXH9c1hGAsGRU87mhI9IkE5UbXqFBvt0oJr4wZ8gLzw
I/FRqCbg17GSB5fqaBwtI8HXvrxbhx5X3pdvF+oCBPVUMeiRgy/6/4XoAKf2uQe1
CMuFKrZ32dilgWTJu+Su00kc8Qc9l3HS7mQcqkd9qK4BCXPosrxghmtLxLZKMPFl
zoG/eJtpJpWoz25k802OMS2tDBX0pSCaPR5YnrstNTIbGvDbdc0YeVsN7/THSkUk
jsRcybEnYnnf0NPN5DVrigSx4MjzTMMnLvzsTFXNw2eVxS+epBzspzLTnPNepC/Z
iG966YaSUiXjMQldHy3NfaIKEsSpFIgMTcOzKp8ALSHnfKuVKb71QXv/8qsainF6
O4YMq62SvaRWAPl3k+XP+oXF2nbGABWtN8HrRcW+5WgCDVM52+JSFAB+u9fYoZV7
SuFmgGbZp055x5FtJWnprRD1FZuoAhP0XvXOBUFaQpQ+VWiq1ijcVY3k1McEY+DQ
`protect end_protected