`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 8640 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/9huKRhRMtvnNqb3Z+UU7TahEoHV+T8U3P3ufru7l1O
3DlgtZzb9QxCbOjthp9+wDkjygH0eUfDrEl1ovhZG63HDzpJ75aaZTdwxyZ9Dmh1
SOqsD8j28kqCD9YYu2eFNF18Mum5m9JH96PU5tNGLuPXWYPYvZjxvQSyWc143gag
Y6+sqhxt+CqGtnWGByEcNsAzYP/WdbmT/91ld8pRmXxx36siToXophycWycKzGNT
TTJRSMqaWSYXJGuGUUNrr3ESORHLYvlqVysRKf7GW34O99Ln0rvSuR38Aw2jJMoX
NiSZ2VPK3KomN8vnoo7o4K2f+ag9tUKDxokk/0oH0/jktnJiEsxBsWlqgdUGNLrX
JWTE1RzVdjsGZdESCeE+wbfow2UInA4HVzck0FbmOBYjEZNqBFQ9BXpwpG5Ol4Vl
KJ38yjsLOeMDrPJo2HHZelrVuyF+V+yyA5NyeduwFFeYQtAWMj2/s6IxA+QxAtnU
/N3uPWTjfnOuqakAFYhARofGWF2Fu0b8valK14GE7HBlzfWX41/n+dG8U3CSodZd
la9WJ+rY/dVCBWHi8IcDcc+tyZFvX6ZR+cMg6T60pj75690gYWN/F2Hb3DxV2cZI
vDYUaTyeLEjmm71ojYnAByiIUPi5yV3jI6TmpD/ShMSyUgottrUgLwZDu7oBvc3K
nJTmJkv8ffZueGi9D38PTkBYwC5ig5QNrU+wWGBnbjQpNCTtGtXv0xyLlXoLu7Wq
3SUEdviS/woqKcfrUAWITr+ObLPz0R2fXl+AMZ72ujuLSE3uaxwkkPiAu4jgHdKm
5efTAmIpAe8q0rwjZqB+awHKTdizdFNj612oMO90V3tTUAlMpMdkXm91+nYRO9xF
ml197yyY+f3L5uZj4y6uVYBng9gB+MSZLDlLQKAWZsk3ZlJp4uYOko+30xoYndYE
LYZ0xcGYDWzu+LaVHLMsTrUwPuJd8lZcJ0OnBhNjmr9rhMfbwQEtw8/Jv2hCCuLB
r5DLLoo6zaPHfKuldLfRQ5ft5dvW9jRCpct3K1k2Oive+sqFiMcAy2+Ab8Tl/sF6
ErH28ZNznCTCZorP/cEWLOhnv6+SSid1o+ofx/fHxFimwTIANp5OkiKhkAm4FvZt
P5RkdwZGNith81B8ezt+0u6LC3vb6Pz8WoIVfvMJ8fb98UMT7C4YgIJ28Dt9Dzix
FzwncR0rRfiGJUATp/bqVA5fjECI1qB00eWo66eV+eB6B7c9W4qRdCqSudUIjn2h
JFlCdiZ9BzD3J1PalQD12rpI41kOkYBlVned+b/Yc/9cnkPfr28vgUtz+BaxXt6W
uZuYV/OobN4L/j42Y5d/A+ElQKNsCSyG3YeC7SPRHYOb64HnENJ/zAOQtUFTGtQT
RicXJMvT9W+LE3GZkUwSTT5lVEYIKm0X4poULV1sKx2zbV7KObGmV85d8J+3XqCR
n5HhigV5Q0soD4MGN8F0pvyZp16DP+3mwPUVVFPeh3tJpIgaKq/VNmObSx6LbIs8
Bf1ZDOfzISLw27Ya+JTijIrZGPAR0nQAH5m1+e934kQZsZeR6+bPtesfdJx6ByG+
YfLNOfvB29ESnKt1y2LLKyyYacrXzSxPHzfSImTMR0h+iD9YqVnZ+G69UOvEajBQ
pBF2PbaLBPsX6hH3hzADpMrD1pNBWQMYiZkgAc6ECtz2m2pXnYXR0R6TKMw/wdNN
WxkW+btEi1vbjBagDBL9E0oC5x7xY4f01LGDeoLckuvHGBB+0yEhQUZbUGMr+2dT
NOwEL64uI+0d5DBUPXK/4BDXQcjl/tUGRSi7FigGieznCRavjx0F0mOm6jqy0Uoe
TyL4hWGeiXYGGppISVHh9OrhgmT+DACHjaQqoAAX8p2E8q3nzVJ54m2GufrWnzaA
sgDBiHwJavnHuV3m2i8Bb0ox4SYQMepQ7Uu8X5s4mnWpibFmTXohXNfApwHdhdZ2
aLSeDenIaQ2HwlBxn7Une4KslP1s54+BjHApB+P4ekx/iV151zvjor5Zw8bJ2Hf8
bEH9TGaah0+uJSvA470vbBJXatzWyk+DvvXBrADaYxrIusTObQ/AXCAddSr3NEgl
OJCDixB/XO4z02PN2DeBLq89d8PXIe+7BMxfuHbQlNETsFPI351DrcIiULxXtBB7
BQ/WiRDd+EKSBUb0eIYNw+uzbBmO0m6uCosnroAS40t8wSLoNX5EXT6mpYTF2Y8H
MTpsPa6uRmn2YWKpfkWya1oON9aGSFHGPAJSo9PHJpYou1CCTkErkE3f/vlKwgBd
zH8lNUj/FDuh5e33NZ3C9TX8GoDcRyag2oiCykMYqxYamxMp0ubcj4NfqvCVREqA
tJMHdMbdM9EqDM1wfsRghdWaPCOIwHlsxSVIu69NAaGzx7V3X5NO2q6EA3lZhlj7
XEQaoLfD0SBdQD6P6hO54NUrJ6CNHUqrt3qJfd5tTxMeLKvNwBgjNpIZKcEVkYfo
LGxl8kHqxSGXt4sHT5Np2lpIoqUdwt8XpAFlgS+2VrjlsGXVdm3DUuQWM4Ep4Ios
lVt0p/9AOMduLxssG3xS90Lbx6SspZueTN50d7r+P4GDjL5nMbh4/Q+a3GG41UbK
4B1ZK8nWXr6gCytB+2Y59d4yKs2j2JTrGCLRBz43TKq0ywFdgcUrjPXZorCidF/k
iUz1yyYslhk4fX9pScmAPyZW6Wvuh4314HTwKEKfGP7JDG5pJLYu2GLC+8tMDwNb
pFnDHpB+8UdbNMV8K5hQiZgTP98RM1nf8HA8q2AbNTHO008thJcwd/ngDtAp4uxQ
sGBAYwphaDZWclcqHLcV86jKy6s4pMzLdnUPGK5TDoevgC4GoPv8eVcoT7pNIJXJ
PrvgefqLrbnj/RFaleAuoQk2LQ7qSye8xB2s3sRA6gBEhFQGcOz9fU5oEDvmamck
H8bbnC+IzpDyxlsxq7c+uN30G/dGytsgZ0bPYT+3qHfFRBwVynQ5D0NGA+M89wp4
0vggRdk4DfHRYCo3iy5Can0EIFNVXA5nbooCm8bxy0H1gBQxAdVqYsvGs1Gg6Wi6
Didvh765B/9ZSJLnVRtd7POrpDuz0+C3ME1/DivjT/zkkPuvx1OGq4WTrkHvOsF8
B1VUHOHOMGyFFbJYTvSxZDq9m9KFWjbTEEsdvfQC+vYHSTKupp/GH+VbIaSPrzpm
Ol8HDz3/nm8LJjaJXVw4S34IJzJl9JYo/hugYGNAp2Dld3DTnu/gZ9j+aj/Byw09
FDTbvq5uTSAx0VzMtzobhn99hMhTqLhhkChRoRcL+JkDFvpeXJVEu4ruPt1blsLY
+Fj689SOWF1+JxPAaW7lUTUqsztZeAKHhkgeUXZfa5XDFY77QXF+N0oTRxT1kb77
zpqa7aI67+2m3xq4KPBmZPUaSNSYKeeR0MJiR5cWrFRYMD8ldIrfu8TtmXSKM+Zx
CKnk2J1TqacD9oohQHgDQAx6e0qTjsZeeIVdWTy2HG55q59iVdUW4QAaeelMYehf
RclbIg2sRZqzVBdDR6IQq9CQ9Ivuo9SiThA1vAT4//MxBtODGuRT2imWpB8Hi7au
1BUoasaTowqstSfNZR2BDZTVY/NadJtH/3aK8/hcs6D/ZRO+1TI5dZHG9ZdO636x
N0ZlEl/lm/JNBGFy3ahJmnPpRMLT1w5b53FXwe104550ETRRzfKxf/jzpPuvLnGr
B6xrKBJLrQKOBXmh8KE2PldwjnHdoT9gYPvhHVjeP9CYkfl7D0/nUeRTgmUGvNzF
TuIbyWKfcJLTw64GRQ5AgoQf/uaUb+HykBP81dr/dwMxoYTrWuTK66xnnauFXflD
+BELRT9S8fB2gv3W/x6fsWzicE9DlhoeK7JIBPtUTl71A4Dt1ASzEPW9cO/M5hQf
jj7OMc8+Wi2LiHGgvIyJYHTzW0DI5vypdy+0G8YQiWf/84YlXmo7Kvg9qn8yJOoO
LF+IKTh/7aROBgMP2LtSMR9g+lXsUWGC0G7LweJ5LYqJMfHOJMh2MGKZ+pFM37G9
YcpS/UAwQsbpHAklDUfbrE8vj4pZl1Bj5a5uGjPROYwLpl2pFwiAraV5IKHuzxlL
7h04/9cuBj6M3JekI2NCNmfH5jxN1/taajntNw00MyiHh1lt0v40jhOg0KQcE7ZD
JagdK8R+nT4f0y4gtHrsBjoOaHRyo7roD5AQZ9P6dsdFToo6Jn7Xa9spxLJrjnmR
UCo5NJGleZ2IGKBH+MOIyyf0A5vu4vSMKy+uaMs4f6BgHLHOAKNczkRjUb0r4JGF
mz+tkaBpnmvVhSt0/Z2Moj/RI6le9u1C085uUdIAQHiJGwma0D49+StzMeLngSrN
rrQJj9rTy9TWbupR7yiPycsdJQBg4yXnANIn/0WuVMdiUqH0M7xbmpnl/dmgxVGR
rR116mGsroh+N4Nmavsm29p7YOiCKdC4FhMCG38JLDPSTQfV4If93lx13Zfc9yQe
01XD6w5i/uB2G+sdARCC6E07XKmkQOEOwQq0A19B9D0mANFgn/5fu3cSYJuwrUXJ
53FGVtKMla27Bb2CAJegCbqlCQkmvkeBDpSamWo/TrtzD5dPFT0o/crqjNMCBwWA
XLhJVTqEiD6jULEextyjhiMfYdsVzBJHey4QcmRSTwNME03DVAQuAIDk/SCTjcuV
GtH3LbHHxVQe5pXkidITyXPmpS94mzo0QNAdToSDXvnkXUUufiIzwL074W/zRPzs
VDF1Kk4QWTHfz30tRaGYWXMkohQjogD0RO6UYp+c3AT0vdD8Hz1RwI6FgMxXCaD9
jEIUsQlSnh+bXbkRXWZHcIiQg13moHMVLaI8swEHi4AO+pNUT1ClxALEfAuU7aJg
lk3Qtd4kG10HdKMNgMsqLGhcF2S2TH3rIqYWWHLXBHWrSvDJr/jinyI/W9YX9Tb7
FcU9V9bzsfZIWqKrlgjAbVJKdRMH5f64DUcjhVLOImm9hQUfsv998VoA6JoollU2
mNRYk/Wu/rD393cQsU/qUB5UvsuFR8yytIf/LvOtUnESFVzA/XaSxQcsXYBX6WNz
UL/VGayliiB0+LhbiP+z9DXnYwETTI483CRx0MMj19AeXGLMT0AAJYFt1hUZiO99
xFG1PWTaPi8S/QwB71KB2h9gBCjtBAn3QQRxTbXyqz1fJMQEOcUmqH4wOWB6sicS
ews+e4XHOyVSOtWdcWrUKrzvDH5T8BXFRAevqJVQlGfnh0uK5sYj6uD2Xha0AYjr
ljSorFj/206JPqCOWP1UY/9TC/iyitojBAY9aTQpwzOtzuBkkjrIMv8M4lFQ3iB2
FuJGCFe++ZKGU+y572ehpdZRYuQS1F+DeHuk1ty5MYE+YvNa/5cZpwaIj67z2iP6
Tkdc4XgP1MD+AYeGQs0q7o7YkumYtk68opqxLtwVCfSNKQIoznvxiqmBZhWTJ8yo
ku5Y9qBA/5KKRwG58yQ+1AniGqOWRPXevRzil+Y7IEaeXdUm1+JyWlwf/y/DlbBu
8v7riVGGgEDvdhz6RcnZ1O1hdj5o0kSxgbvR0NRq/O9jEo9eYHvjHyqtDDqGRLLF
YOq3zbZrnHE82e6yYMAtj/yxP8E9zD9CXFsqdC8Zg5pEXtGvOD2Zchx60s93ARZK
oHJ+/hDiNJ9um3Rf6i2wyvP4b1pGLd4qa3t08um/k89T09y7zsSp8+suAi3JKPGb
jHManxXY+/Iy95J2GS+udpr40plANf7zZUtMr35WxXjxeOMHaPB9tLsvkcrzCFrF
3qHWZ1GM62bFvX34RtefgWtBAcDwNt6BhOq9/IcPAlVMm3JEQI3SZpvfm1KnGxI2
6I93oyLb2XCBjBS2WFQ8O9oDdMiNIVPCpuMBtX7jSiiwPR9W59GXn4RabMnhP0uG
Hd//X4smFK002Kbr752GS+5IpvWfk1eqd3mXI0gjmp25uIt1Wgkefsffmv4yvCFV
fFQK+MfkMRW8sWeupZVokvtZ3xE73c2Mkyd4a+L5MNDGZSWU86KPp7mfiyF9CfUh
mvPuuizyCltqVvTgbUa3528QA8kh+UvP9t4XPXYQi2HC2uHExccL4U5p2R1iv0N7
xEd4e5SFbC3bav4Ucm8QCZYUW5MMv9WdhF0OUwutB587gYq02i3q5UqgkdhZ0c6K
L6HhI0+Ubyy3U69kVvYVWksx1RMtG83xOeSWoI06lenj9LvdUZdMoCltncbERmpN
qdwPjAvmG/CV6+XhEbAal6rZKwjqGSyivISuClJC6RX5GwPj7kPLkb8GGORFkhWy
yQKSYwyQQTBkDeriZiecDrwnl/pwZD1axRwCNlGOJE7J5P/BpMBEBc6bAEnpQxsY
BurAHoieixRRl9kFOxyjqJ06+Amy4DLAM9JpFSpIBbBEPyING/tDBKL+vqteS2L9
p6DRjy9CJ0ADOwlHxlTaUjNvoWQDikf9N76iRUscURBALNpQ5qUCJNPDUKlh4D7u
0CBdh8VgArmxGF0hmVSUhT7UUJgU95IddG65+yZkSwN9UIBIKP15ZluQ3vf2XX7X
GDnqw1NG6iYJYs3VNhwxlXFEyxjRpubF6r2wJVw9mfWM2aFbXoCD0t91e46gKvwK
v0t7OUsGl3cfNfxMMmge27aOryag6ZYdFuEeSMomv7Vrro+qYfSvrgYkCK4qVag8
CtAAzRSfQ/l3QenX7crQeXVCCO0GmVxz+Do9qQX6A0yNHw8Y2sqG8gH12Q75fThv
YIv/KtgYwNh/CXjfvMWhqN0HNP070B7jrjnBDM0UFIT0Bp3DeB/BkbQl3Fje6ZRf
i7ABgyNhkcb+gW1RyMFWl6R1amzfO05XSrVqu6L0PhY03O2BK6jMjwFCxulwhZ9r
vT3phf2lUE0vmDr5blD7ITRwQEHMJtYp2sVMNtJD8X8EaW/Jam0K/ZljgAMSKTT2
KqxTtNHLPNLcdMFIAkkPlCxAGrKqttVPTH4U25hqkEzYcHO863o5i4OJvPVDp/Wp
AH8mLYC52xBBPmzJDMhvgme7ILBA/lJ0Nn1h89sVNblIeD+Vv7mIktOfGJc4M2Z5
q9l3eDPh/UOWoKKjVWLJFRJAwKFeQyRK2SwjnPf/4Wgi3gm8V6OkjkxGODdTfEla
ukPtkk5eCbhnxIz/LqIWcsfw36YJqQvASd97wJmYFIsOW8379otAlcWUSogBlEWJ
wfNvScvcEOakeDKTMa8Ed2875dTRO6WfzNJj5woCaCObyRtqJ/YXRNMaDb534BHk
EEuLUUg4tiupqZkhlc9xzDsTQD34HVpCe+nahZqBV/jXSoaE7vTGJnGcaDJx1uj0
+PhRuSqbGQnAa4aiFNgsQgiaRU0pXAzELL/sdIOTN4EDqZX86WOUyrDBxwV6hkfZ
O2xxciCukXx7yXNDV3upCVoM4Pbt9/voW7V9nG8WZlstbEn2VDodPws4N8B3LlHF
LLlTJPEt6Rh1+79kAE0/jmTkOhXit35hFSrrgEUFUaX4MVWQHRj10YezoQJtIMLi
r5LkI1cQwUG9a32IoKMUvZ8AayJQ0UqtLHEWsN7z3hRVX6pK3MBnaeUIzQoXfRnV
jKcq9ErZ0eGFx+wGtKo2LZ/WbaBr1Fxh9xiuk/zVKArJUk0JxQzcCt1AI1JIa8K0
PYGGWm531pazSq1n8BE3Tq4SXEaQk6FjazDUhi8ctHoeDj/F0HzLdn6MkxDZBmOK
wtBhXiKt1VH1S99vaFxQHmeuuS/FN/kSymE/Q3PyWbgDXn0uy1cb2IvqD/13lljp
k/dN5KaQ/k7tNK4V8RSJ+HWQvdiXy7fdEKT4voOAPaHtuXbuFWKINJyTmXbTurZY
+nRUhZb92WIlUeMYDMnvt6cJV2X2rgDXPmGRhJ6GaJpmDzaMI2ERYIykgmi2wGFZ
B5zp9ULrRl4NirYFiV0TV1daqspcVVZKsTnbQfZr3XkEoOzLSQvSlf22o6u2cjDl
GsQl2lcWQT4UDh4vi7+TVQ4QVvFHA9fDI/uuAA4zY38GrQt+wR6ACwj1GhnMSS/F
AkFARF0Cq55JlTKbDPKp7U5S5Fei3dNi92cl7Se4b+/Wowq+JypCkIoKyWQbe6vj
iwDfA0IBbyeiK0glcn4gyIvpGwo6eg9NEqymQ5Ynh6rS1gHLCCv0T0mzsP5oyXB5
hcgictZpB8NaF7MUZ1bmIrpOeboZij6+435yVAABpA0FXbVA4dN/AN+d5u5W/OEi
ltnlzNOnghNFRJHZBGDmIul9OeLSbtR55U/6OFhKBG8VXTjpvbBiiivh/fdSthw3
Mk0vEDAgxxUFU+nBRXMiCqF0IIJjgEhNtRsOFe3Wv54vl4zknc4icehho39tl47K
+RQCsW5cex8zfVsPgInj4G1Q1lTa69e65PxXzM+7d33ls8eUbiUiNN0pdQ4zW1N+
anwuUmiBY3YP4bP7Qv0H1TDDvtinxwwnLdZiejL2OU7AddnURyhH6zDXFRvUiXxF
YzZtLl9k7XHG1FgG3HvDo6MxhJJ690qWsbVebb2dHoA++kMocKKTt4tyLZrDh9Zj
dEqPmO0e3NS0NNDeI6PLV4A0gtcy+T/Pn/Gr1gaBoIlJmWLcLBqnA/eq5J7aJWHh
NZ4FOC5DW51ZKSvRRWRib+Xe3TsgZHe8Wn0UpyIOSJq9R6BtL2bwg+MIyRP9N9pA
OonPWvxDLyJwJLNQjxmKHZGA4XafRK7QvGzzIYyyMec5ypRmmz2MN0EXkKvJkCU/
pEVhPlfeu2U4voMz5nbAekDAjgAnzkk5u4qFbBfz8ARMe8pAv1Q+gqdhUJhabkxJ
JKfQeUTT4mkM63K/wykv+JOrvYev0IHxKSo9Hv+I2KQezsg3IDRRWasRYwYYHrj3
z//id+4qV06ThVLWze0Ols9/nyF3kzZI+H/H+bVQFEzdgBxgjunI4BipO1YTw7Q3
2AA+AQTjg+JyoNapueKqmNoQ9iSwaIeatJC0W0orZbCoLOdQYX3ykRIKiRF7gGH9
KLdBhFlpkRFI82tSO7Qk18PlYTdeWwJN8EOmw0YqUc31BRQMPN3NHeMffWGVWy9d
AMociKoRzWT6jtvf2kJGhWPaDgC/Y99zjb4YtEqcekUsfaURXS1m3i7pRCfCJIUD
4UQb4rfh9rke6kh23Zrb7EMTwJJqXae0XZ2a7oxCc1r7VGhs6n38zllGOeTw04Fb
pSG+fldx1LgWdHihoeMEkohDbvKq17qytJ+KiPsRuOAJ68VYRSEkFDstyffxXiEB
Zv0bywOums10Rd6rWgzBK6utH2eMqM6UUSJVhzEBMKAVNBilhoBvD5fjlC87uow0
qzplW6oORocgLxjjRGfAudmObop3JiAX7wS/SN2/9wiRM39SsNKZRL6GCPYQgd3C
wQrb8QIZSWPsNXKh131n6NvvJfzt+Riq2UqgnF5lz87/efEXj25YQ6DUkB0JX6Js
tHZXiHn6ezda+upJR3X7u0uCs6ocsXs2ndE+sLd2dpPJIG5vQhVsVRCJ9oDoHqmq
Rs4CHey/2gFzejS4Ok7Kjwzd89O/nZv+rVHR/kamAOAMmRofyVfE06Zh1lIIQyAS
93JkbZsKxFRQjlzwI2Tqh1WkWtLoyfYpG8sY33+noDErtk2xGGSEeZbPhmYSGuDl
nIpWSIKoOvzpQWCD9KCThmmBBWjz8zy5xms+XgLD/GXX+jSAEiwqSF42QN1HPifW
KIlPu+PTD+6EPQm1MXUq5qLiYCVRG0e2oSRk6ruCFTxbpS1LFtxvWMEgGL2x9j+1
lKp7Rk7vGnaaQ9kxw6d3+wfA9IW9JV9Dne0cDF2SZf5nFfKBJnzR1ym3mJeAoi2C
HZzLYDlaaPABctlH/ZjBrvnLUm2znxUHa3Y2Be+41nb+GD/dx5MVgPr1EXFgBlt8
PuJKbA603FKq7b6TQU3tdTN7blhvNiJe+DBjcZNM5TI7xUKEWk/Lhl+4OO2BC0PW
sMEVKXO6LgdTh4kxmTVAMKkvy4B6ucatKGaXtcrX+ndTLNUvXfouLECl7QDnbn9j
uUM2f6JmGjPvqu7vOJC5ixVHCGzr7fcZsHlWmZgABRVSgxvKKWzQtMyQSe9ZRF7B
oB8itaIGqFb1nNV55F4Pp6kG/VBbqyuaBdiQZwjAJifOUKO07X7Lv5VBvqZHRKRv
8KRmRUuA7axFWOY7bj6hESvXH+Fl6fRZRT3lY1ttXxQlfoORWGxRBlEBzrgksuOb
uWALB+4LUC1Lf0W2V+3cL44e3mShUJ/eYy59JBVbcXA/OdY0EnpX5+x7FQ0xnTh0
STPYPUPQVucJ8HPX5RQcKgJaEBpSNnXVpfZC/vrAQI9Zd5t5MWleMFrOt3NNsQXW
1AyOla9E3NQllZNqC49d5G6Wms7crFipUO4cwvkoYQAbr+EYiR0RRbIBxnuDA3zB
Fkr2MNKT/8fmY4hedlkVUMAWdo7/8Zh13+iVauYVy51FPaCtgqhCI5AJBhaHYRYw
hGxaDifmCm3dssw0LYL0xDTEG/dzWAQ2rWsz7PZhHelh/3d8vV/ye5bd9SD4wqe1
9/POcjkSdKtcUVYHD+DsIFiQB/drZJwmPRnsvyt+0ZViGYm1fpe2Gf0Z2ziAYRny
SWNjkG2wSK9ZUT8vf7xrQZgkl/hIf6OjrgDow2oLJpEqB7F+QRpzbk3yeBTZOEY/
vZRXeGZg1335FAYh9J0+yBdIh4TP1oV42vCSQFSMvRFOlxAbtkYVIqmizfgE0xY5
rNSYyyDNdC7vtZ9em8iaBr+r66eJhyU30/dR9JcX/wArLvtCaLp6lBOUiex/4a/2
/riV8r9UgrTsuGda7RVz4Wffp8fg9CILLHTKZFQPWX9tTs4QYX2Kv1i8k7klYCot
64P26DvdrcvEe7b9cinwd6Z8v98EolITI+6PxgkovgFS6gqJiYtvmDVKXQLt4GVI
12f3GibTx/j2WWDxvSBYt/uuDpN0AVGHTFl5kheIK5zU8K7GI7MhET6Klmchp//O
xsKMQ9WVGntPPkyJxNHJOtvNYP/pj87IjzaiS+lkqI8DlN2nTtNwsDutCIF44dm2
cdgWBD9mM7Gn4lbAyP4D/ZXTZqmUgUovM1MKCxgQj99tjapkNzCc9bCSvPS0C5gl
KkmR15ghkFsY63emybS5xA/XKpZ8pgLM4h93S44lCm3Uaho0lOVfv2IZwAzikviJ
1CfWR3+Z+haUVzBEAogCVG3GTbHR4wjfrMhin0FR/CNFaHTOnFnX9yrkErzFxLuX
5AbEnwbce9+a0XHT8Vzxm563UhGP/YrBBjuaFdawxhn1SeoBGo2tTeC9gsGue7qT
ujdT3Jyiz7AaZvcC62+d5ejwZdTE8BPfOwNKQkKopaQI4Nsvup0sPhQ+QjgCQ4yV
De+z1LjiGIfqVHdW6b3N1OrOHzZ9Qh8WXmjkDg30PPqVwg4NM9spWcPPD3AChx/s
Ka64TfXblNTJXGSK2UpAvD2LlkAj0bPnFzBBFaHhX37v4GRMYZCllnt8b1RXCoe9
IEQtGW0JUV2ZVz+xAhClo16AOoLSuqzveCmSAgtiJ0Dr1Zp0SX4EPhH1elThm4eC
`protect end_protected