`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 4800 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/59UwEX+aE7FohaWu0/8IpTj7mav863zUNIsgIH2BWb
Abd9opeuBjbGF/waQMI2vMJTwD1ie1YueHc3nSNpEh4OXp8P5ybZFY89uyGz3ztU
W1EsuUnchJoQgbHZ/sLbgtGRgsrAFn+ZoIeGN1d6RAF2wAESJmYP8zw+p00RvjZ5
G2ATm2jrAjm+J6bPpiDE3wiIQEsp+c4GG4s3G/grGn54V89BW7q4R4jqV0Ubt5Q1
d0gZpZ6WaxZJhI5vUh0iuurgFRHNiP/KNj0Oxp2IbKEBH5ZhSGEes+e3MVv3wnQ9
FreYvopWDBmTCL+SwQSAXgX+RYMg9nBIaOK9iT2Z+vonTWPUQe6a9Ce5FaL5AjT7
MvE9niiPQNrO98WE9QexX4aKmQIpAbLmJmgKqepdLvmsGELNHCK9PggEqKLFPC27
U9hQFLo1nrdIoXDbKAT3KCJVzly/EbqoMIEa86AtcVxEAFJ/bZ2x81ja+liowxJf
VUfnTcrM1H4hI123oQkRVBybT7B+FFeURCN69PjyNy/38dKBpNPooPGLFncmO8Rk
SJrdpNm5KriW7oDfI5c8OjdmyvQuNdF1r2zcyuiXR8NBqMMLUmmwTT+8nP7Cf00d
Al2jEldLSbOCeX5H5cJmPWnzpyFtSw4N0wPrvL8H4MuGezFAM7aXwzYp4F3BEn7+
Bkbo0/Y0mlIJZOTxSNRRLxI5LFfP9Nz/beQFmz1W1L0e214boFubCqYbllY4G9A1
NlL6pdlj+0eE2/qV3U9EJpG8eIqTQtu2b4fbPtgz5ZLTyycqUipdSPz1ZnDTMz4h
CTsi12JmOyCBaz+mzaXp4hZRSWYm9F5vIvYWt87ovBGTzruGFPlqfPjBWbHqGF+a
vulyeBLC27pYjdGAc2LQnJsIEOo6B0Rlg8GIzHWTX3P9sSRTpBaH4XlOKpn2Ddte
fGjifRJRsagK+7UGzmVnJqjeeEhTD41fsyuo4/GCRAA079M2z9bYeFZILv8Xgr0r
KBmHZwalFZhLTxS1kZmnDVlm2X+TiHrEn+bbv1NslTyw1sN9nZkXaqiXHRq1Kqfi
D6xExScE+L2dIxpfQpc2RBMoJCdMXFI/iqposX18zH+xNeNRygWD73qNa5OVYq4n
eA49sT2zBd3dtZUMRd2n15Bof0Ux2grEFgzMmwPHC95ydlMjS/WPJlGrrMqsger5
kVdNAMfUM8TienTTCzlI9acTgK/BRGk3z9fIBMkbY88cbXrPEg/OlZOrCTn54pzf
IN2ziDidrDCfNoLjxHiVyxJoUUSF1Z/zpd/HbO0jpocugeZC1DnF8eVHTzILjQ53
VqLZnytJrkfq9MUsLduHVn76F4KMESBjF8p6X2LHwvQWxGAuMwCWFHWVa7no34SD
rYDdcJPeE0jU0IYb+HOAWyQvwKNRia7jHCk8p/W10UvMT5SMlMRFiWIUX9KjPzv/
rSHj8B048kxSwPYGV16/t4bYNla0yG1CrJc0p9IhuykjgFyEBx8OkPhB5jhu1E0I
MU1qxgwI0CFqd+C1Mhqo47kXiVxGBLnO/9baeuRJTamjFHlW/hna/30gxct/K33n
bnsls0CKLI1Xc1OXcBAyjtund8UcOQ4n90P88Khn1+PxPmacJcXwpIQEIYxho1Bk
XDunJOEqBwqnkTs9s6PUS3n/M9EVIYizPObjNaeHwB2il0qH5wYK+OIQ0A/tNC1O
Zhon09uA+dUUJlUy0+NLNVgXbaxnUsMO0dpJLeIvJQR+XLvhpV69v6qLecQPXnQP
De9Gqm2OtCi75Ac3gYPYkNAgFgtWOcOTQF3Rj9ZlsO2e2aulaLBRw9tQPtV3RpO4
kRjv/b04y7R9p+y1e0vgyUiY4nqDG7wgHH11AQRIXlY3PDANkNiYL2JCZn9ozRuo
0f9IKIHOoAakvdcZQ9OM+cqyb8AtLcAhZ0iVgbTizjmolMdmlGNZGJr8VcEJSJne
Q7shh24rRt+uaFUpuGZs3OQEjjNf2YEfND6VjGCwNrDme0LjtjNsFmzdi8WxLHoC
uqjLVOIe+sxVoMnJR4L8ADvX/esgDXhALdo0qxRQhqwtGI04GQsPZoisTviTJy8e
X6aoCo3PCOtdEXqIc0Rf+egXigkUyETdBYd4EzXSfccrFWawh9fs1esYwa0ZcFVy
oLnjfNHwjBgT9QNadQXue8iHxQV2xn2myOSRFrQWRZ9slyP3pB5w9iv0LmuWKnSS
Dw0fLrfMM9ajUAYdfSwpvbScB3aVFvVrrh2NGdqaDT8eV6yDAnb/8rLVaMikU9mP
dphXXbZlVV8Sf+D0SPGzCkbBW7IpAg5X405Y/pyxmmJCQ8RpdEhp4OphYQWvixCM
vI66FJ4M1sNBygaWOratT5xlJ8eWIVRNILvluksxPxHkY60Rq0gH4R5EG1G6Npju
z7iNY00+OWW05iUBrkYNI72ziKiqDi7M+iyhfL/3Enj5t+WjzDDJ1Is91As3GpNj
iLs6pabw0uIlnD5tGE3xYCbRU0hGMwMWTQOvpyI8s9WhOhRnNeF3fvCa38lGPrd5
oWbno5Iu5fKlUP/25AeMim89GmpH/UzAz/TiayyOuzT/pYRCRII9RBto4PxwSydT
SSaM/YQv+Np0KCsnnV/eIx9UcINd8iVcB6ELE77upJxUhW95i8waKfbMbcSsqUOT
7TjIXh4RunYFXET22kzRawVZ+iBv0lA2lZ+4hhJDj5r4LjLZBGunzIsAIByZXqS5
BI/Ci8mLbDQzzJuMJqD5BW1+XRblt0JKHs+E7vWI1xHfryLaMGf6NncrxwWrQ/Zf
zWtQTwnmOpqZs29CsOsMqINhw4oa7bIQjZLekjVH8BSpql6YfHJHkT+Ic9pbgE2A
5lsB84WssvMfTomOePvx84CO+X7og6vChf/kabeyPrl068F8kFkl7tdZX0LY8bBy
U+dF1oB2tpjkoqacvoFq4KzKDj7Dev467V/MTXKSrHNYrGvYaCnSgR1UTSSKQQgY
CvKgCRvuoF+P4OLs780FmA8JSjYORLR+/t7dFLbdIBklAIEPJd9AtAu2wQeFmh8x
XJXGZBYeDywiPBX2RKDmZQLp7CV4oTT2LvtCQQ79lOdnygC9bFGIbU0rmSniSfiB
enPCBgugZlw9FiY09EgoSjN4QcvLreY2wcsXVDO63TpqwNnhLDYjs4KL1XWQafZX
qus4B9fmitJZcD7l4exv3Czn09fBFNKxh8Sz4Ou08ZypRIDuuqUjij3i7T6osmuD
yXdFfKNLvpNH3vN5UQF2Jt2zzhFgNFFOViuc4qZoQ8d8gErzzhTQQJxjUef0kipp
eE6eEsJa79NbdQ+Y/9GMVoPxfuZjP+YKpLaEq+KcWeT7fIlFYsP6I5g6m1uwQWzj
31cN7OnYQUPoi780IwWJotZJ5tvJSlyOfH0knWvjMCgbC/tQt2cRYGa8ZNAzA6+L
0x+3FsC2+xPTd1RYedkBiumkcsJAdORVEmROlf9mxPuBSVgBGBD01ls2zdcN1Zpw
/s1vmtYdkcEhvln4xda9sCx5x/26x2PxNjA3HPH7UaklehNx474O75jVR9roA29+
supB3CodbYzlFcnVJNj3YrnJcyLoCj6QWG1dJJBIFplNFxUhF4lnfmPvv2rqQyUc
/0lP0jDp0r1gnFOuObwxpoJtMhYkSmbd53o2eAHM6b58MaBjhxMBR2VrftiRIJtM
fUAQv8P1khDqNPFK1D8ThVI+h/R8W3Jwjkj7OfFDm9Y7tTgOPC4czRfivqRBTcQv
cM8+WvtZj0btQ75c+IeFT4iNo/DkkUZaRys4hib6azqoetIRA2hELfvaKiConb1h
EhW9LZ/11VRgFIDCEe4zC8Ywr9aqXpiQlfiw0JyBeQvKRDU9WyiFfXS0xY03oBRl
C43JXT1rliLhyjujLa+5ykZdEm1lI7KeRSUR9LBzBJBKDIptaMk7YYqA6vYxxWf3
3Yp5MP3VrzU1OEupVRgCkMRWQtabckOEEoLQ/jfSlgShyKpwtejxbbwyD5zB7BrD
wHBPH52pegiW8hyXWNMW+k4cONFISlE+bnhNk4Ze8zfZjNjGAY0LHMnpGaz7Qn7n
dyZ+6jywT6mbh0BdLB0j8Nns00tOvUytvkS9aBsDfUvkli+62i5vSgKtnunfrxuB
eZmKTe20YEFZ5naMTOmIcbj7ltx4eatxOwu77nub36wHGzDCeD6xEMsLs7JoSifn
F/URCLa5srgF2rGdVVnYt9dydtF7PllhvGq5l3NiSoraDojm4UN2wYYFZ11iUjXd
arhyRnBkoNu9ASoCmy6ulCHT4c1xF91Kjtyig0PERs+hPyGYoJpzVNRBNrCAu9RH
XjIscZy4n38XKOUs4A5h72PxKH3IGphhwwwCdPerVWe+azjQnvlTIkrs+gqpJSKu
smVHVE8VH+18mAaVdF9WT+8wHu/DeAtok/WsXnZjVuSUVoU9vFyC5mtiwh+WSru1
4JtbmJJo2k6GAgQLVcbmTHTBCW1MDtxC1KD1OzNaYYKnDrl7kc0b65fSLbARFnO8
ZfSyZ7HmXXOrWuiiMt6BGX0+yxtVm6vByDvR+KPY1LHjhTEYZisWr7TotMbx/En6
nLo26tZq1i9PPGKBQwvbbwIqBWCHhD7V0F52OcNM0EM6DdMMEM62gxzEWBZQkitO
phE4umnxj4ymU/nxbR0JWSfGDEDyhhFPUU6GYrkovPmgp1BmBThqV2I/A7b4uC3H
bEGE8QUFR9Py8LVTaC1CTaw3W3N5tzAPcCsQR58+OQly+58lN5+hBvqfy1c51y2c
pX7cUw7ysror2TwGCCg/K1LxQa1YVRCA/2T8Jzci/+GTDghgwC6VzgjslZhRAjP1
7joXKuDXOdICQRkbn67wwtmY9/hsB1a7Hhjfq7iNmYA/QWQt5OqLRASes2WpE8TN
qw6ybMCtRChtSpQfbvoVtrbDj9LROdpOP/XDYwKXbfK85H/FIdBNkWhdAeR2b2sx
TzmtZN+nnNK4a3AFWdj9pFRY84B0UPEbotrTQNOiL7n/5GIp5xN4BOaLW1za2Jp/
QhrrftupX0aEknwFTeVaGmg2ijkXiUoMTNRtRfLOydH57ZOCBF/cu7kNorYyXUJK
aqQb+6Qcq+3SRnexWq8y3Q5ii+tqmKYqH81zW0dlRmFtApz5QuCwn5ptrZhu6h1R
Q1heLyqJuZwMj+vfyliynvscmSroT/F/rdrFvrTa/S/3IVyLiRuUEji+LFCMutkd
3dTLdvuVTF/C4/K7VS2FgPtZMOtezee/BDyWBoRB0TMZWk9Xz+YuMfJ0yjsHSXbp
O/vevwH//PlpTG0LOcDA008v3jTADBX4IJ9lcJXHEBnKZMBZ+d7iK2/FpwER5DZ1
d+Rwds7nh4c+/NRh1Q9L3nM9/snQ+sYIwsKIsupNylTFdVHUCx1m/6KlE9ggXo6s
w4dZydVYWkqLWMj2SzCh53nl2k9ZkMYjZpjUvYjC+p72Y6zhYZK2PpypjXxlASnw
eFpGVbyRytt+M1KVuwJx/SsTvyfCBOdsEvSP6D/eiG2I5NMunkxvIiYmjTzzRv9I
p4T3PA4we/lbXuEQP4676Hh5nz+7IC/gh6UyFER36pzbscpNrEV6dWptXrNRLJ7b
GFBRFTHRK/raj9qorJvvM7sRmry4Jtu6vLq4EV40TvSk+zqXJlpwMK6nA3JNED0p
M+MxTWEfLRrpl8j7zkQx6EGElCeFXpUoH4v/hpyjhhJhaWaSE9lmwRYCQc9IYcz0
GLRgBW1cr6ZDNn8AeagIBOiRTJfqxV73GnVdhqixq6S5MQrh19wUMb1De+hGbEPF
/JOTty6kqwCIZRU+FJCNUF5SYUDINXeCtVji6dMm1KmyimgCmdn/wo/DzmgX+BXc
ewcyaDh0Ptr79f7qAirsOOv1VLSalXiudlGsN1DZJPCrJj0Yoe3mIa5XPVk82+fE
5nT38cBMZk4MB9PQQyBoo31dEN4pvgCnhrcR4I/md3T25pP7H1JaY84fiIkRGCni
iedr1j1NGmMnsZ8rGcM4SsDdFXC9CH77awkhnacYBMCuZ9oME5bl6AUxoGEln5Tu
XfMu+4WP4EMdURLP19Ve9QQbh5cvPxyf40XeoCiqrxv3QF7y8qbSpw7pmUii8mgV
5118bT77MwTIOaBw4jju8E+gKRK4TZPYETR2XIvQR2OwrzClM3LI5dnkTydAEUaX
iiC+qsax3ClFJT3GrhMt1aVSISaitnd/8Z3P6+Fwr8cwSA4iGfBjU6yD3M0Uyevb
VdqzOt8mac1dpvNlhBtXW9lAtqW1dMHMG137Zfnva283i+trFaoWk4YjkWYaPZkc
weYEuuj1SbiYJkg4ejunyvyUtkxuL4aYha3WbmmC1GuhN/NWiUEYDsbmgtVBQrr3
`protect end_protected