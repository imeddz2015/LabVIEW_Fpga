`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 4352 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/9huKRhRMtvnNqb3Z+UU7TahEoHV+T8U3P3ufru7l1O
3DlgtZzb9QxCbOjthp9+wDkjygH0eUfDrEl1ovhZG60cQHmUfNumtGrMuo0v8Knk
/WDS/Dy3Lbk+rjnjX45XrGfANVj8dku3vhwEZE8vTvO8PcbJ9a59tY0i0fEy/4Ri
yJrRnRXZaXma1CLoOpO+6A66ynLDQJ/MM1ods2Zblci7dOBEkbeE9Ju5iTyIds2x
Y2FjF9dVosUUekLRYQqtcIho5JZ/LOxDPBdArOLSjLBQMcvdAvTlIe1AfgEyKP6e
JYvkC86zATCmB5sprqbfl79eMqVBsBjXqd9nSi7CUDEwEeKhp/SxQ8XaxnAXd3n9
OZmPs34LlsotT2fwfPoInCJHc2MjlCzcMKD7g2b4F9LrVBd2Nv2A9QrvAhqe6D9l
btygL6h+EZK1FWAQJ6Sbx5fU9Z2AppEMkEHkCizPnDB5tjUSYXnp+5RM3SfG7EVj
aRU8A0am5RZqHSeyc5xZGqAATpc8Pnb9cEPUKuUeuy8JrVANiP5RabWVriLWTkXK
0N8MnbMSuSVeiE4cIcVCdi/9obPc3QvsTIogjGKMKvwrr8Sg0V+dpqvgjWxi6/rd
0fWEj8RLWOpKILAYUAj5A5jgtUuV74S2X0EyfyWVh/plxlAccHVIkBpjE8qeK2HD
SksE+f5qwQ4fvB9rgShUkTdL/AN0JU4KJkRf0ArisiNAj4DA5hx3suuMUmLsREkC
X7yGHqpHa8a1Xa2xwi8DZQm0jzCcIzfODg4MDg00TPKgW9V3zR5XdTnMB2VWrFKu
zHd4mLf4MfTRxgrpmn6ruRBv2wO2VPHPh4QpgfYh8kwyb27dBvJtuebdLPVD6aAP
C9Pcva7M/sEEAGQUkE9WyP3k/5rc32s0DJcBHDbMP8FsgzYPJjfi78d4VZqKfoel
SFAA/Y8sHFcInbI/2F+RJJB8Ib/CdVJpnLO/dZFo7A7qau/f2lZLkfZLvrlzQ2+9
B5j11t/YGTwZ+lkgR8KfwY1J/t97QFGv32ezKWSjgzBoPikoTk20nyf4Lu26qPGn
4Bgg1O/NAJTfM66h3jkVA5YMNdqs+trqgr3BXZAMcSvPRhL2lUf0Qk6tZiAxvCJr
d12POcXoIhjUHCLcpK8q+1B7I1R8kQ5HksicN/ryQgDDRwyMhFYH0z51lq3HH83p
zmYa9V2+Rkg7VMtFqCIMGiKx7biykaDv6yzsBqg/f5Q5YJYN+vrgZy0lZcSzdJFg
lmoKr8x41qjVSy8jGAq4t2+63sZZwkiJyJIJGzvE4xA18IymR/nKfsbRtpla13Dl
geUDNvc+m0ts0UDR/cH1f3sWuzuJ2dt8sCIF5UzBPQ/KP719kCrHT0pwrLMjvty0
yamobFG+XsaCznZmflZSnY8OwyW88uOPSw4kqQaYB9cjxoOigKtTE05WdG4kbTEx
x+PHXxtR9XFUiCQP20ovcWNoi+UQSr/xHRg27CJvE8TsCOhuUStm5jaZbOKnAQF5
kp3niVgFB0dG4o4WS00OwEERx5UIcLdxm5ftWH4kESoBcYoquGK43OlePLFE9zJC
YBSaokCWru4SrjHEaFMRhRQbEUUbJ3xLsgqXG4NxyzdqZmJsxeoCRtSJhfG0f8Jd
hW+eb2EuoHoq1qj61eoU5lJ5Yj8OKtHSTaYryUNxH/sU5Iw0HBfSwhgqlql24God
BQE2x2BFCNIswiHOFCPvmdn59VyQi2z/5HLAmSDVJpMkX/fVVQQtKdGQJKY8k2QZ
aHytYsya7KDeI7S4/DPUM/kqNWmcbv2kEUCI1qTy9uHy4C+UvhGBJjfwDhXqe8MS
aTB+vm/ytJwmeNONEwUQmaenH57ImPr3V5uVT38JQDIVqH7zxsgkYyfUx+swb6CB
3pLXEBSE7wh1LW1JrpRRA7jQ/7C0cr4DIOPc4te4NqZz9051XDMvUnmENK9fPyaw
w4Y3Wm68SXp8jc7eFb70Dgf6wDbyMBIu3hOMhADEteezrSSCM/KlPiw88+GsOIHi
GYsmCGEOshcUYXacIcR153Iq4AWAW1hUzudhh4SRAWa4nh6XNalq+vC1AZBRFtyB
EcgcujpwA9oGoLEeQtIItLHLWUed4FTuN3Mfnxh7wi+Hk3IsDsJM+vAaekLq3NYW
mvadnI256r0GiejI8MElZ2pzScd6jH7alwIylwsDlaJQttWEaNqA8AIGfpKP14Zy
fHsebLSASHOr3goEBE3xlCTL7pxFRO0UYG2w4X/1KZuSO1y3iwwszQBkUz5vyK+s
asNUp1eip7NQA/HLMKJdMxt3d1lSutanfVHCkdH3qRX8agi8ZbrpgcaEQ+PTCQAi
nD6f6Al6/YpqWCaKOQdl+r7PtwwbMrLWx3tO5MXob6GkpeEJwTzhNP7uqoqTpzuq
sovG0LJh9LK7+LY5Kzjw5SyFuFWsDhGoso75Bjhet/X6FofeOvfRNd9Mq1wrotMU
DpD1REVchnw62glMZk/MMVe6v/BAblKL58p2XEzcvcTbP75BxusjOdUhvsZlbAE7
v9HA7pjOMTxFdJhfegME89w9azpoIECd9p3yiiPXuOFrdpOE7ua5fT3sCld38K2U
xpUbSFWBsYojOs7xD5tWvm3+2aMBRGQ14cAf8y6oOcxL5af9Rnsvh3iR3T2nPzkv
TmV9TfAaX2+yPvH4J7Dy/aF0ultn10ZjV/Te/dVCmUkHVuBtWnVumOX+NxcNGTKY
cbZD2v1plGnI9ZjYrrEcigLiWiAcPPHuRNHJhOGIXSgPFO4wZ2ISvPYVBMSPpOwQ
KnrCF6xaD4Pv2SQo3kTNJ1a7dfsgHczcSMazbPVyQl56nzotGSFvjt1G+In7f6QL
XoyPes3ZdLTAcP5JrAsDKQTliqhyLwzg8e+ruhxMSLrF8+aRo/T0YuSxw1dKYRME
BUHCvpkb1YZxH4dNqRrcmlDkvtsMCrnPtzNIqZ4SYvIpBvDVGB94WwjWDEvugFWH
8JYq+oOfBcqI+HS0Y/SzeWDLYfMrKkHSWOvK35fRDUNqb5y1ab9QnkQECrNqeI9e
PokUwYEpaBKDBDtbVe9ZnGN1FiWorh+J2FOPf+F6QHiwLue29B4CbNGxQMUwHsjI
fc4Yg/KC1MZfOuXvDKaTPeTfmBtIMd4e6ipm1Wn+YigZuhQKFBjqzbq5uTTJ/264
rwgAA4yZf3w2QtpiiEFSg3MYiLVm2SrTxZsWGe69rn7hO+rDuuS9ijBQw7WUxI9+
wAqo/vUTBIyoHpmt5G8yOysXi2CRZK4w5BFPNqd0IQTQhVedQXSze3XiNWesLa1o
9XW0XffPb+mAU9fK0Sfjg+vErKpk2EK+Gs5rrGRR5QZ/n2AEwVOmNiwCoz3NVJYX
ablQhvGeFmZZeCb3Yc0O8UXWcZ/OzlNh43H3ify+QIRlmFJvnzX6dXxfsPFcDYT2
zRgWpE4gOeKm/MRq1G8cGRP8cgd+XqVWu30EjhIpBoRKgsBk9t8CirKYPuvc60+K
8gU4sKLnFP8grzM+BoPaxgIch1H1oYTsDe3dZw4+NommWoKyR4/96BVhRr+cXXGl
RZ4j2LEiEd5f2C6i4wIzOcpkgFYMo59jedt+Lz+YqPe6LCowQ831rQj9BgcGmX5v
EiSZMPaMQKQcF6E/cmyFDH5+xkSofEb2Y5BRzhgmmb0dRyLTL49tSi27RQpVGtzs
1111FitTqPavgJdWLO/VM1yBro/+v0ZV+7sUE0yv7ByfQyJQ8EjfUvQN+19cvU23
cczbhcvqNOmnBUhrSyxKbRu40zUf9nJXz1udfCwiec3rlTU7EOKqjBuZuejA6BXR
OOuqZ3D0y9uxQUc8u//cVWSDHQRHHSN1iNFNMmyc8H6LfTz2D5lzYbJd+N7LDwD6
53PyVgPDOYRjJyXAXbUZi9FS5YD/4WNk4o/vuGB9QzYD7aQYRVK+kZ+LVOOpVk8M
XiCnqFo3SkBGJEH4VncTb4maF9tH/svrPrM2huPQqXW4Tl7xRbnE3zktTsBBAl7Z
XUhvUAV/lpmboZN0dvaICwanW1TVk06EeAQkl8rQLXMW5NvvinmCVelLd7bH0oM9
qJh1B9znk3IMSWjz/UIAkY4X72XSyiLkBmPOLcARtst4LTnAJHmffIskQWjN3gt1
GJrqeB/1hcBpeHKaZvXnWV+chYuWSvSmRGVcLdy1Xcbb9x5Ilr88FLmaWBcouaY3
FF5S7VX9FyGhShdudPdYMFpA3adOLRqeW9QueR0TNHjco02JyO96AZzeLgrZNBtW
V3ejnlr/AZr+ON4BGyHCEKn5ixAZGq/JvDX1sMit13wvGoZBv45yKOz+HeLYHm7s
3XWGPiAcA/wFKxreQS9ZNN6rEVtkFuVjrpwwpnAB1coubreUZxqvXfRPErHqPKog
Wriz/VK0kOrGvJCQgoRdw1h1FitWtABZEVvBYSCtO9gvmajQtZWREWok7+CHJk+x
pVQpdhK90mhUqTASkwF6QYrwPFJN64pu73lPfgw2P7wAgKY/y65CWqiA7C9QViA3
Wj3+LXwQgYTC2L/ofytYRUyYsUvF8SYe1VSmyHh5imjuWzmlgRgNv9RH8fQ76PDB
XhXKGvgmgKimh+AbqUZkrqwro/P99mnyXTpq3WNgM0o4wb+uS58nxv2rloaTojYZ
r4wbvRAp4MqdU1s0axu9/0pEEQb3XqTjTOydySFUVVEF0bjvpXVbrnNRi/bqndzb
5iHJC12Bq7jQBXCiPPkjqKwXG3C5AYCctMZYvxJIWw5WWnVaaH+6S/bpMWXvO9Ko
3YwqYxDLT/fMjnpP5/Q/AENS6Thxu0f7rjHfSAK1RtQZdiceWMfesma2v41F4t7E
UIgycK0MFhQE+5Kr/EhW+HQGVkioJ2G3EeSLzDbApzQ7DmnH1oV1ZZ+Tk2KRX/uk
ct2c8wglb6q4bu9EeVQRgzrWQtK1MLvRi80R9Vgk33tUZ470yG8ExH9QzzGAg+Rz
Ugp+5X+f1lF5bRlOqF5PGBnHJ7NRpqADKxtIhomV9RynvC+SwFzVv0w4sVvlzCcV
Q+8VSjH+WER5kZCSjK2fk8rAvUbQWE2g2GAsg56JMAoVnOu+kctnxrbjVgiT040O
VRolIeOTkBENreFOOh60fvGFLoUfLVykAru5f8QVdrB6wvQ9bbAy65+wSBevzceY
dJekN7s+gIbMDdtL0dL3EePIgId19iGZh6twcM/vTuMyEyqExQcmxFhqi6LJ3McS
UAd/kFg90Wlq916n2ScKfCANigiYxY0yUisUYGiOFap8VSp2vyN6DgxdwrRbRZIz
Z20TRou/cISqwHz0lGTzUEwgfx5hXLdV3WQt+Ch+w8Km/cA2NCxh9xzHuTACa0wc
LF6vDkMfR0eZPErSsjK4lbymmb1hcEHCi+/py6U8E50ylVD1a/CbIvRRgDAThecV
tymdNfj1Wny9GZZW6b1V+y8q/kpktWmhynT3dXszScNAC7uKNfTcFeTv31wz8pzg
SFx+ppfLJL0pBdoXkFEJucCXjNzUvIRUlyyIA7tcDZs/gUGWNhttiqhiwVf17K34
Xmd6r2Ci6Sc9ieTErcn6pUHeXlpu45VsFUr+d8xYxv6c9U8vYG6Ou5jnvqn4MhfG
e5jbmqQbwrQahTfixp/NuVOhBodPgQ2YosGxO0TfCAI20E3nKn2Ai8XVQwfQy1v0
xHeHgHwNynzleojBdKR+TPyO1PaplqmoBooPeu9YY7u4AaGSBxrLqGL9uWuGU8lL
e2iAqBdsl3/0EDkwojpF21+Ta+F8KKlMDa1LgLGQXZ4=
`protect end_protected