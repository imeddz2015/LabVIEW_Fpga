`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 52208 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/9huKRhRMtvnNqb3Z+UU7TahEoHV+T8U3P3ufru7l1O
3DlgtZzb9QxCbOjthp9+wDkjygH0eUfDrEl1ovhZG61JQ2OcQDwSwYjEV2pAWuEe
0Wm4wH9KDATZe4733kRLemF1JTBC74PCBh0vcYtWhqaOaQKUJqKpMRBMbNpbMaLJ
56z2ZPVIql2jztuFta+EvTpKxvPpdm8J0QUOCzzXwoOO+GTrTakIuEW++7pdM3Cy
5zv+UYWLxr7kh3yY0wkBkFc4KLk5E0TftblK6Qn/hwe9FDmM7ftwC+8f06xFtkuh
GNIrlCgQ52rLuA7fNgCIxJBJvtqrCb9RNeJSFcg+qIlLsx0a7c3ckIyjN99p6pKy
VT4eVxGloyOAGHQreQZgmFQQsLbbgzstNzAnjn0lysQcbIt8XoZPqggQsqU/1yRE
UIqfzRitifYWlTKMTvqw07IRKOeZtscfXafjHK5z48lQwRITHJv1+jHxV7auQMKx
a7sHRLYep8vyBntLoQAQfJ+MLzU8H6vkUB8Z3FxuwiKEAyJHAEYFuwPXjEULconT
heobheRDNZyp0FL8JGJZGGunlGwonrquz0jOzozeKcAL7sPwOz6hgfn8zZ2+8iKA
WmPNBUjsC5Gqy8wTO6axiq98dplisq200dIfju5tHPgYeaz7Z1n1LErna/gRzsi1
0Z7swJegwTL0QTjNn2KdWYjx62kfVxBkeuiE3XEqKYfKsW/RbxDk2tA6igX0IPTI
5nugAS1O+mWeQ+0WvbqCWUd+4+dw4vWa03m5aLz07ATbUPlckqhTd0SmxC2WziOI
AAYrbYc3bm1Ru1t9xmR+ugunPHJi7tk0ymQ5Pbl+3Qcf28AJDXMHqUFLuGn7L3iz
nQvJIO1x/U1WBxdGBK9eIUL7z/CIK6QAN2H9Q7EPVbIjnl3tHfAlnJHULrw+4JkH
v+WAWD1V2ziTI8uWn7ZANWdKulijOkIzpV6EVRMZ/qNHRy6UIdAGxWyULXUxd6Nj
KCOIj39QDclFpOm4MEII2mqYfRXIYfrXgKfo7xY6BgBMP50f4HXMLxKOm/BprfNb
L2BcnGjWuzZuCpZTTNtfgD3qCmMX6zaExJ9qPk9kutwJ7FE2XIqsEGFLYdXteoUA
RACdsCW1cMnm+q3fZrQtTByzTwJsQs5JOi7UmWICVqEc6manFt8pQE4KzZIqm5ss
EyIVplsE2+bekyMfBRbsubvT1M7dHlTirkJbUwmwQR+QLua8BLOhlX5h8MI6dQ5k
kaNkigWCOgwGom1LHgClsFCNoW5e44Wc7jaDRLWShokG2CObNVwpyypgnhXw9WSC
SYwgkL/zQx5k7S05+mexUvLO9KYBdO30Ypsw5q0yx5YWZyeCaBPul12JPWdfY8Uw
ZHW48KsScPpqE3wvuyFd7CJ2NoNal68k4+ZqWIB6tKXreFtbUHVqt/SxZtTwmUn/
YawhNzjp+hbj68xYbQdQhAhiO4XmDrxfqwNYwMzACBM0bTitsXZbwh9wVv/xJTGp
zO2hGvHVMxkw2qg7l7VIAASr2Wm9yeC2QZDpzKwfXTZRpfxS1HB3mqJDmaj/yEhI
zrYYVomNV6CgQnLBe0/ZhNteoS5wWJIgAR7q1f1DDIB/1L7tKM16L8rxysq0jy/2
0AwisRsNyQhokZ8jTyhO8tRfhpxEiiz6Uji21jWjexPuAneka4XaVblZN/5zXXU0
2jVIhHshC+vHP2yAX3bIilgEVm/03Di1ik8cJSfZvFlyg/OKJTQvWadQxL+IrZA0
d5DKY3/PGXa+ZngXfiPsBq+Wq7aZrLgzABT5WciWqqM5bif20Ynb2yTtBxtEkOA+
D8d9R6gqVDkJsklL+K29QayiBgvc5eFDEn2FTSCCkM7C28ZxKwh5oN+lIMVntojs
QFt3k1NvO7fynu+IDAos9cf0PBX4MGO1OEw0oh2cuKKQZv1zdFTV/Km58CfJM6iY
U6xGRExr+ff6eRjiI/FE8FPlpv8Jyd+6dprrsL48c5agtLqBKTP1uqPeV0o+w5tS
+ss+5n1jPatk4iC0cXl4n0cMVvCIdwsK3oNzc7zRZN+K46lc1SkMkweM3HXtydZN
8YH/26EEDtxzxwarnEMUTEBUDuAYr24RXDUchonLZM/FYZ5jE8+YFQMequtByzNF
SnwLbEoq/5+Qy1VwKQRihptHMc8M0llRv2yjGhe0g0gpY2lucyzVPlO1W22QMNSl
/OQr+tSvQD84Zj3i0276Jy0pdSREh/2lNrKSS2+ckn5lWZiLUjTalyKZf7GpkadI
+ycI4cd5hjSfeOHhtWmPE/HCeOVa0eBsM6uFZLVWqlE3DNuQO/p8jAmG9OLjlNfi
8kfIfc9XU7ptG3DU+UlHk4NnlR6pWHJtAXF5W5XQbRWuwpQPQ6bIV9lhfx1I/cW0
OzEin+U3AW4iOprKL26PKO6xDqjOOaWgFjl/xLky1ukNaxqFJaq5Yt1/y1FYx5Ey
ileiyigBTmeGPpXDg3ihLa8TuZ7YzieIQSg/eobO1R50al4WGc+m1fQ0PAsP1kYQ
wAnjEgUmfSC4VL+i2BTwGEWOIKPsgojaZmtNDTJ4TS8xQrKTSRUtH4tOy0J/gwU2
3cHnQ0NDppR39wVLxjrtQiTrhpSb0ZKTK/0gIGw3IqitHcoELLo3PIKr0jatbdvw
Yxuuk9e0rzpI0E5yyVu2fsIMpx8I1hXldVbF+PldrW/Q/PFOparfvzrmUoLscvZ7
jbz/UQv2Jh1Sp3We6hny0CMAV9EnyuPqZh/E7IpnmKJ72o9vOzr9H/gLF6dB261B
2t1uKqqcx1B7/m5gXcgV++r5KGZgydPZIVtPZrwpCbiFvVAd/agPawUl3R8l7Lfe
mHyvFBqZ5M44arlMHP06khS1oX9YU5ebCTqgtR8B2JHpxGIkP6o4VmDyqObHNtBf
/pZhAa4iLa76OMIXrDVcuRzJ0tJPqQmotzIPKx7XKCDygCvDJI7DaX0AJuJE5fqV
UVZOmQB3NBJXJl47QgINqDKMcWc9ircCKSLvgrkLVkbMk2bOLwkpTdRobElqkX9u
2D6/xPalDq0AQ9yUQ2MS56/4K/KIxY6TPwJd2IFMpi6ky2/r0qEDGo7ExkTlgsy6
4q6Ra02UVLN5TGltp8cY45ZP2DwEFZU8Ft49TJaWt0tZenxzvACTQTvtkHpsTyNr
/UD93ErNM5+QuLhx7a5nKcxST4kOwbUN1YeDQgmfKjjxIxpJTEalMnzmuaMvvPpb
CK3CggnUydn4xVZNeutRyUytPr/3YdQjNzf7IUosP1Z+A05yLD+tfiMkz/Q0D/GT
Q5IaMFlxyo0erh+TFvqtSP2zM5x85hbzFcJz8qQoD41rVcN7hRuPkDcGV+sTptn1
rsxc2VF/vwJaGPBERhUZUal43ih4FNAPriHkLTucNWKvchWN9ubMhDh19G+AQU/D
qVbn6tGG2eWr8dec0GeszdS8PvHoAcpPmRutGQhjy97wLaQwAl4U0Uf3xaeQ/ZwW
oleYwYeK/m+eUnMZ0X5QOVpSZngGdW5xSvd3OrD2Je1+KtBQ9cmjmEo0D6AFJoYS
Cpb1IGen4tTNtGjNXntUpfTDzlYVtSwG9h7OmQQbdmJkYczWDOI7vRPhka0hUhJQ
+pd5NqCtxPy2cVjw9uKJ6Mt/BobLeiFMZa+3DxEmYaH0X3O1/Y4D/+0QmtscmTRc
LKdOIrHDsJVMxW8Rs796MGgyjHLfQY2wiizpZzhxgsurjyIY06pDS5bnkpEHtop0
ktIC+YdoSRJUs3kK0JMCZomrUqgAHYMmSL2hxZ/SJF51mQTqJi528fVDKB4ZJ5Gv
7ltMQuWYXrsfmRF8kS+giZs5At3+SFWLCUg6Ip4trtQ9Oz/Gbmt84LcKfWZs9VAs
jKVAWvcHE+v5hFmVkQ39YB7QGYw/4wY29QNIRiZZXlDptWpDo+2bSwFyr7fo8zfX
ghAud7o4lT8uAKiaLvu9P/4vcpeQXRLLc0TKicG8PlXzMGETtUrSFIVe+CLqtmmX
ALaUQlWG3ytgczXFsmUV45CFX+c6bWtk9xIS8rR/pJ2ZNoftVIOe+HxgKu1ZtdHn
RgkWPEEwbqUl01IHf8/3IKBETyMwHwNGWXze96Q8EQV4tfDp1QmEhVcobto++zqL
uhCss6AfRVdJDYH3ZjcycUW1pIZZ3ghmZvs4JgIO48YEANmaXVJGYh1inWp5xFiW
kYkvf4JQ2ATsx7h9lfRLnYIYvyIo4/zN/KFMGa/Z3o4mLXJlo/0HeonSkRjVk+j4
Tr3JkZuZ06ukCbCje9NvPZ2wqwYDMDdxKhyBFTf5HTMKm0PgTkcPk3pFeNBUE1Jk
As4oM3muHJlAk1UDflrJPxm+1w3SSvqWP8VEoPxm3w4wA4hC9UVF+zUx2sIPChq6
UDwVD16yTHZjVD3UmWlKqo7YqB9k6nImUNzsRsTGPFtGqfHr30RciPOzy/h1eI24
Hy+77hknUpjCZ1GThcRLrafFB+U915qhmha6xkC6kGDnRTDmCatxKn0uROtPPn80
WOVdNWvtvMst7pVQf6SAU9rM7zxY++AjeyUQwwiuI1/mSd/vvzyskLxJajEJtyxP
8ZJyGC4b2VwDtCjaMZUgW1nqbndZQ7HzhYM2+I+bS/FiVboxCXQEXjTZWepl7655
nvDDC214yhLLonqPDbXekJiBnktnObt5yG+TFCeGey+kR7ZTUx2BCTKQDLQBie4v
M9UyIO1q+FnRPfcyyCS1SmVB2txGd0UETgr/IRjHF+m86icgZ8uHdcCLdEdxHPrB
6nQczmB4YEkVMU/CYWm/2Dh2af5xkcmEIsBC3+PCWG2QLQMO2P3lIPxYXJZwMzSz
K3uhe31cH6oJP0jgZA87ZRXHg4gHgxBvWaxZ9kIv5Dwgk/0jivh+bhZBIVgev/Vg
VtMEgsgHPOx6bcWuXA9GVIXLkmABydbk/v/Lx5904huQXUAXr30ODM747m46SbM5
ELUUV3j+37rW8rzoj7XFazButLrsZk9wXW1VCXPb8zFXIwtkQboKiy5s6mtB9TNm
Lkub7j8VEpC+C7FRMd+uu3IWt8JcsUoNWyBUG3rXUqIDO+e9N4EhdNkQ/YcmsWnz
1lzUv24v97FbufWEflwhKZ1NnTMrggQlsBnljw980xYycGdE4PD11F/gg4KLnxPr
g9RDoih5fZIHA2sYHQwea/o9wrxQJ1VE+A0OASbTNYIzkskmOHaoIw6RI/HjCT1O
7iAiceG+yyhz8RezCa6yr8lx0rzdlYviEV+Ha6Cay+uSs1nGbFzDLm8lc/ldq9GI
osmm8OO+d1C12eBlo2CPQaLmMYqhB2xj1/F+iTU7orXvVGzMk4WDQdaZUdt2arX9
MansvXxKHy0GIHH4qbX29S3nnLScrP232ZJIJUep7lVPQ2xgifVn25t5xIxtvHBR
b/fjLPrNilV7+KSG/TqmyT2RfqV3h8+jowrNZxOs4T7EO4JTOeyUEZ+bqn04fvVi
LXTop4GK2cMGqEwcnRlv7mOOgX57IVCkvYgKHSn3KewhIq+8rjOFm4h8EIuahDrX
dorHT41vqaOlII/pGq9xoJssV4+ILcRQ1KUTDJuIEEoAkzgMuY6HWnhwN/AzkY1Q
4excLJogabAeX74Px97B06aQwVdjuen7Yvik3Sph40MgzBn3o8lUAXkwLrHGlls9
I0iV6sSdT7cmyR6Kbnv8AnyTtRiTtLhwaS4ll3rVl7lHaMzfC/NhodS6G0omaiYj
8PbMAZantb8wclGhNc/qVJ3OBPI81VKVqrQdr79dg1LQL2I5/9nEfLyNNG36PBa5
FUikShPVxgYL4lS/M3p3S/cvO88fM0NINK24SAGGbOOU17fGFzYHqtL2vcvg7+ey
w2O491KLxjSTt93c4K9vxNxzol44T4FFZxHhlFSZPn51vr7/ue0HueHpPElZTtgd
FzfVzYabCOCsQ8CeTfHJuBSS3/jTE3NYGd70RlPudZ9mG2hu3RjwLL0YSSbsH+26
V0Rbe2vHZ/qOgT+CVATiWePt6qXgE/moBLnhyos8ISYbFke1Ow3YrMsXhiw8UX7n
a+J/0q3/fak0ebduHywXEMV7zDhpbfyfBtMWp+Y9WNoezbIwn/FSctHImXbE+g3G
5OXLoUVcPlwQbx5fiUD9g/tr4aSMw0WQdiu4Aa/D1DCVxAl6NozDSmVoa1RpS5H1
ISoEDdDQ7rfCoS2B3pys8KiL2n8EEskzD0Uur/saJAaNCYo9IyNvgJ3okw4qrjir
Dk5Q/K/emUj+iIgNmdtYm7+1K4JHa2SepjYNs23Ajmpq6GhvGt+Em6ATjCL9JAJ6
qxNDrDRiaQJapJoEV+zjoawByQK0DDGgwwriBxmxwEDFeSro+w6OXT8S0HC6a/hB
HhWtnZaPkYIt95/SGL7FAkcEQbXcwrvX0QdsmHRBtnmnWMAj3FA+4hf9DAoByqiK
3MEuHEikZ+y07eK4W1Gi1JXfFQkvLPl1m0IYBeDmEilXaXS1VqipEkkZxGbEn34g
6I2wsRLm75zLtnE4OTXerTqImPw5vrup5RpdRjgsRj62yYhtbvbffpF8PaC0DvSc
SAOWl1WCqGfMMtKLU4Nq5JitZYFpbSSXwaRlLbr+JYbAuMazuuohVb21Xgv+yxJM
Jffl95Z/lxFaBfmDYwfUB677APly0Xtkm0b7JszQohyLoOw92eVJmEsNlKzdT+Iz
KPBe8kxz1YDjZPI7SwipkDeQgQMcMYki2iTtgIaqhHqEB2jePwpTWjOWCoCTVVvr
d9IwUWEkPujYUePa/gyddnvx7/+/UOHrCryy8P/iXD62HreypiWcsvp5dQmZ2XpQ
x+3uYwY0PKvxVd0BBfU0UirjXlalqJ34U1Pu9HCtYL/Kgx6aCaw6myKPGdjB3L/5
DSA1XnHCotswOyNjfXfXAFdLp0rqr6Y91e3XHLwt8KS2dJ+mSKLIkWc8wLHKNdQe
MrNiyogF7T8I9JmErz5in8dVp0udV+GMKl7zJrOIdPcbeS/gFOdmRxAbYL1w8KCB
qD09MPkKYJJKdz+XdDql8srYPco50yl4JF6FJmu3nv5kmAmFmacWPeJflOlgYC/e
H3VrvE0Bt8EHkHj2/XFqV5rU10Q+OHDJpGsGpZ2qrU9ebupwUEoTFjf52JFJSAMP
6fzFSpJ+hvoLSAfEIxdYhZ8wvfL+FBuzUha+4SJlTvm9z819P2tlUd4Z4031Nnfk
xO7g5IT9+MMxp8QUMfuxwx5cv+nJDvx0QGB+DMXpwDe9n4NSNeMjg+dVxl/5baR2
ZPRv6qWMw9J+2ohY/YRGDH4/AQ2eANL/2/UT8kI9cQLeT10fdjKhOGaqN9yUrEHN
p2hXA9zdB1fIUIhae/72JT8p5OjyIVCnRcnnBMizIhbJW/rmlv6DBqV4xn2emf5y
4g9oCwhMQhgVUCGkmnrdu/nD/undvd5KGZXGxvD94PtzJ7ZB026I1A5DzqhzFFAR
mZqzbs6ZimL/wYtpeFOgkx3Kydg+hGsOAz4Z+p9I6z9VMjjzBmDBtHh15hLFynD6
k2bK5terEHiOKv6NSqbGLKvKWFA7GqAfCEwKJVzas9edLUR66zRAjFSvdn1B9M56
X1BBh8K6sMeIXJcpLmBGl0HdnSUhkSgKJKn5HFb8zn9Ncd7waYBg2CNhdDAS4qY7
xIljREZ4wrM+xz5ZTTIhfTRMv0Vcd6N2jXqPQ8ZJCN+aHoIHkwDGqx5oojm5fObp
p/mZ83/VRf3OSxaCDC7FkDkC5dR1uNF8nVSA1q7lqj6IYOoqgUfndOHZPeGGIKYm
xg17THNUuwKMQiDwIlctidy0qylqp8fesqAvC2rEzCdtGMoBlKc4lC+5rwDmHRis
Be7GW7SHAqXZrL8izQG9w90Bx9dX6qjd3lrxoZvRxd6PKk7ySHabPrvRIubleAeJ
qiwjWN2apWAhtzb1Jbsm3cS1wUaH70dQ10zNsI/OvtmBhbGhOeuAjZzU/7hapMU9
XrZpoddNzOmeymzI7tV6gypC+opvjq/KAC0D4FUrfL6T87X1DcKfdscLpdZXaGUO
6O+wkqEuNQJ452VHe48+UOq3eyC4N/iKbuGOlLyQzUj+2yrUMOHHFh/If+j4Wi0b
CL0v2GOYr6iARhzTaoN62lCot/hFq+i5ieAtA14SBPe/1F6g+cHsa3ZKeiNN2TSC
w+/H/84A9E5EQlIsb0d2wH+w+zN7i05s9x2M1gB2x5sk7O9aPVtPaUtVBABhslFo
+86kaYybQ0FqoeBFsfXyivtONyRTNjy2kTFaB84MKK/ZaQJuWrw7G+WsL7nWnSzQ
8a7fP1ZaKe+y0dOEbVKqycN3419IFWd5k/hls/+OW9Hjs2ooJ/04JPPlSsdmGjt/
LOrVCTeqaZOGtCoJFVh4DqVLy8fG4jpd6B1k4vmEyWTp7PqqiQp0psLc8R58kLmj
HyF1d2iUbHTDP3kwjO0ihtv/hveOGzksnIa6Etuc1D3+GUnnB6vJzTihEC7xDjPl
MFnQ/lrF0wh7w5I5nmV99R5AJcHIsKJuhStsYY6mc6h1y8NKuw0wvD8hhjvgXhbg
OdqCMnODpGsEFi6xvAL+S2bAbUcVtC2mFCuu7Kvoh29N6Fvv4EG+/xKS7khzeymS
EmDIDfJbKRyflz76011Ov5/KCKTCrUhqHUEG33ZLGEHUfHBAcfNWR5Fq0PWUOgbD
EFFG0ojyG/cmZPKjjw8hN8Q23SfIBE18a1cWm1a3cLH9r0mTGitIFem5YRlQGEG9
2JLw4sk1801PoXFJKKFJJRjMO3WbS/DqBaF+1XwGWhcCgnQqj/2Ot8XR2rfUa2gi
gsx2su/pwOIW05MtXdVf15vmPr6GSUDFgoxll6/e7R8xnrOEujMAUxgPtC/xkS6N
NLXyqD94VKy1ABFhW59/iQP84WpH5yeam7hGwPU/qc4tCtlybIbDpPtVQmIfTD+g
TNdxCcA5/5U1EUzECdb/QV9HheBaW7CekosHgLbCk5ZvjFs9ZzQ/vUm3onlvUXEr
ntwirWZaeyXD+v/QxBADgDq/gRy5U6AxGj4kcU/uLg3RFhoqKhLyson8uq/6RgnD
KNbHhfCffCLciAQ+81zo8KL0kCzPaINX/Wj24JcFtw4UUSXR6uXMhvyGSMo5WV5K
OfdlzeFc+H4rZE+qPfDU8CUbt3atiIPFhhPtsjFF9w0CilgI2ZimjYJWQcsqpSta
DyDxHfR0qWhTYi3bD1fVDUWEIaw2UUOP2bAa12HXTqRdyGr0l5YIdZuymQuVTNu0
IKVfIBxTvzK2px6utGmklBLmf9KvrD2OeBd0+gCqiJRYHrLz71KU9L1IaqhKB+6L
U/DgvSKsw0ww9TpHry7dsytfVGJuLOFm0p2yCReE7e9CN9PJpJLIhHy7akwmRHgF
7HimK0G3tL3IUPpBg7J/2+KanrAm8zoYrunGHbcxePMoklGEmuvqo10R4wS7+GDb
7DgtEUjESw6XXx5HVYmnR/NRje3P101ej7cBzp7PxJhHxLZpmYA5UQHEDocO3FW7
YoADNjUwpFnDCbkmsK1rXZmiJF5TSgVtQdpc+Tt5l8iYhV558RFsmQ4JmxM1gcHL
qaIhgctUkmk1GmHItzskPv3o0xlxvQISArgk401iZEne8yBMrS2thKajC58/FaTa
Tpfp30f2lq7pHq3e1ilJPlYtnThJ1TOaMuQ1n65+X3tmJUPQzX4UQKJ90qZLnGOS
O3qu7XnT39w9+YTTGC0/2tqFtXFZfzuxCsY91t1I1zv4PqPEnAQ/8+iaOFolLrkB
prV1SfvPItYQK+ARUwoSwCkbcrElHHinksD9bOw/YQ9Iwx5MdWsRTTmssQg9hQKT
wDOCQ3gdsmoULhu2m27T3kVzurEIgsS/mXQ2sdYFUk/OcGJdE/CGqjnz7uoe9uzs
1TRYCRORnhrc0hOY3Nrap06i+1WlwZaXaA0472sodWgj7TBXQE8VaHdXc0vJuNbv
aRqGPdw00ThEtrpK6SIaxKfxSIgxr741K4U41r8C+hcFkNWmblPaCHYBnWOq3+WP
R6EByVbiVmt55LK3yFFKZbFThwi/X3PppQUehsJXlICBrzT/6O3L1feBpFK4PLQc
leSBZ4FOl7HmVSYobhIcIpqKu8ZxKUwYE3WZqgY+a7R+64dfT/vQ95BypFYvk10D
L/oEDnsycdIr1nOZ3VV9aSOaY3WBJ/Ve98pwqXXtH6bZQS3gSjkR56Obu3LgmekZ
x1bmHiqW+mkfyZ6wCKDosNUCZcN1srTmfyIt41Qq8em0eA9dg5eaRtj/nzvVtss4
Dv4N4hdpJgOi15nN+x/vTxQbOc7R2yM6VkemUujrxuXIFdcDh+RXcd+MYsdBt6Lg
tcBLZlyGHOrcd212X/mMoxtz2EClSkXlkfgpBnPis5jqIP5un9CHaz2oNsR2Dhs3
qz66aMmxcDCu3IhqJEiNOh1SJWr0rApKLXK2YuHIXz2MNC8fVNbQk1l3lH4mGYij
Esh9Ai2d1HGzo23ZH67S+p8K3P86g3hXwc8Vf0i7WwFy0SvZJXUuXqmm3G0ZEUPQ
jcT3FV3hTbwVQFnYiKMNh3EUXuwXo0hZSihOKWbZ6ju+yHlwydgudF+J/p1PekyF
JDRPg39TKRNqm/qeVz+uODAxbFRyITNiJe1SA6F4God7pCIGQz3aD/QgSTPFNEUR
TPEdS7tr+qc1Y5BX+lVk2Uwynuoc3XyHFcrRCPs395N59oXYbVZRwjlShCNC/rCt
k81vQl81Dy3SjjBaGtWlNLRoCYUm/L0dsx89ReMxaXoWbK3g5jln7sdUjy0aP0Wk
9kDCNbrEOYHbAnyrCzFXxwn9gf7Tcn3p6rV1rJOa1H4cHD9KppVJnUVyQVeeMyWl
RvyakLMo2NhQweGVLkyC/2sYkfM85UJ0XEmaGXWdBbo/Bdoaq6ClW5z2h1WLbEaN
g5ZVRpmzIuh7pfNe2UyoB7Fp4r+prlVd4eveX2H3m6/C/GZmpiqVfvo5LFPtxhCz
2WyUfzP/DGVb7I0eiyGi4V7DgaKKiwVdxbZmEiegypGt1FycgJXYpTz8hrpppO0I
/BZkLkBq2iZ+8agJLiw4UaaGv7mMxaYQ2jTVXzu+GhE1V3xmCdDo/6JeqwILAIaz
NPheJ8b7ni8SLC97Lv2eV43Odz0zWW4JncKdOsYhs5sEx5z4YCiTKLRDfU4sbv8W
IK0EctY7FZnO2fMe3+u7rb+geJ/D/pTvVHGD5Fb2v9NqHqJEoZ/qzFK0W3TaH10M
4pkmI99XUvynH3jKMxMLq8jTDYdoP1SQFw2FN9mbBDzs6w4hAbFA0L5pkKwY7+NH
PC0cOQzCJ9IgrHvt7r2RgxqtGalonKGCpvBpXSQgsIuRSQnkSJ5fDtS2rKhsWPDg
aWpwRVMlmdGqvup81VG948JjqwKaljyJpSrHqyqQG6qpbyvF6e0SSWvZ2KjVIFMm
iqsz47xf42y92GtJsI+n3zrOV/WdkfrczPd34JB43L2GyXfDeYIpyhJBFWYE/6oH
LCpnm01TEvRgGFUDZMYblYdmsKi8lDrnqOjkhqMTMNrgWAoburK12ZlPVhTB1aqh
BTz8B/7Sg9Hkftk+23jlFY2iSyeD390+gs6XjX3Nn2CValFzJfbMfiYk47GJvj+c
MFbuv0tRuiY+W6vZGRlqrSQ6RI6v/c7aErquSTLU1NnQse2bk3Zcwn3YvWBgtyKG
PIvcO17YF4prcuGxSJcpIdcqAc/yRdISemd243rH0lM4sGYjeS6t5hHbHwPBUkXL
43tZWT70+dQeeuwd8thw+5qCsBmFdCH3ZcL5JxH2pPhGAj35DdGkuZUzWqqB7X8C
bU7YX77mRLgEXXtb6ZGKXA+GaoqKQ0AiKim3EBUHFBP2E0H6K4bq88rjVdcxKlgR
hOqMeRqnHRez9tjAUfwpONsOznw3bwa6EXmt9cr0t7vRa4JUa0xen6pRdSvixUcI
xIe7DPOzLJacpwFdQwrOCBpqZqzXLtufZrNt5kYi6lrvsxCWsZKp1XlPsjyRxjQL
Lp+aS77Z6ahZzFh1Im0HOZe+XT2fM7kc4nXtHbpTfGWR9WtgrRuPYR0ICdrGx5Qv
GJBo+HxfUAJYfRWzAOmWd61X6nXdywJEkR3cKUolZyrENx3CNw0SbW4AclAMq5pa
H14EcdTKwcpefYkjIN5N6kmCQnEgyAUg1Y+kj7YnMoIM00fs148mTvMPncJJtRCs
0PfjSHJDwbJmbF8GRX3g+IXcl5RMgc8FPPFT+kIghzQHmMSAWODKryWZTRT5HE1p
aK4Rm7wOC8HO7GLWeIsSZL+1XDLmfypO4AxeowOs8gOQL5381WDRvNomTggqVFRy
oyI38wxoYPvpb5VPthdDASu3sLebIz8PXapS3fx/Gs4cRYvXvqJgQu6kraOiOvZE
PMplc/jNyjXzQq8YSbojbBTnMnmG6HCNg/y6nfxvKlrPZxQAWSgtKvQkV/cx9Mrm
bkvOVosqGvx/CUf7cZ+Y4+RyxFa5QA+txrxcFeze/wZzKbe9WJjRcGNeruoiEkCK
yE3n+QYggUYKl8VH/0GGq3u4OXaQsR+FDEjVruRjaMfymuDIFjGrxJ6Ll6mZgki2
DC/Wat2XBJYlesJGjUh9vOiQMzK6nCka+/zcXfJxLwoPo5jD81+oLbF1sxnyNkRC
HfasBu9S0egbKNmquFP9heMrIFr3JRUrKG30s4R1L47NXcmdIBIFK8xIvZelhOFH
+Kr9G+UsAjqGCRvQgOwc8iFKZNO0P4BIvSnVPKSkxuDKmbvE0ic0JMFjdW+Udtmr
swSu5p7e/xGsPbT4JgdkqPsuX/UtdFNl9XR9ga6/hKPrJN9kP9V07sb2JngOyfqZ
KMksI4pab67Fm/ZI//4MYPim7c5KCTQNd20BW3n/J3fPus7NilTClq+wsuHa/r8G
RU0tHccvvtlbGE12ZsHRhM0Hi0Q07GUBZiUABKiiI0lLs6AeOqosQssp2U98BHQE
heQZLUkGv0oWh1xTQlv3RyxXbJt2GCPefI4Z0kvbWelx3ry9rSM3+nBGyVwjaV8W
JN2OBIdHHasAu6JNGEZamHww7IeGk1l+9tjfk6jZ99q9EHVwsfnCRkANLr7Cl/i1
giKWtZQOn9o0+yhya0kotrd9FQGRkn+yFiq8WVTYG0TGFNT8AoDk/8/dMaxiffkg
aM8kC5BtKKe/kAyhDBmcFvL7nqnWIVBnWGE9N7VzoiJPFcBtqar0vGpEkLzJGzLY
vG8Jr32xXDcvx9xQbANSdOC+akhF4Kc+qb/KZkmz7r2lsJ056RY/lLJt4KqcF2s2
q+ttk0xS3r8vN01MwAgxohLLQm473cJ6drZRCNvA2YU0oaD3XJLppOU769dTTudD
VLehiV0PahYU6XH+9A0UbQYHwxfQQ1LFifKk9RFvTwmB6O7BtzFLOaUzg9uoy3hR
rzeJ0gbF1rGHb2uGzGsY9lgCi8/i2BBrAAspch8hqQndutqCDGuhpWMssrigygUW
zj+Yxgh+kki57/CsH37KWgNrnZhFkSZccKoPD58Y0i2U65z/JzMnfeWxG+Qft4Le
YZJtJNuKd5/SZk6paN0npvTvUNXI1KjthC6Lq786KDDQ6SEy3t6kCIDsjFGQIS1M
JMTb6zRUvKWlH/rMC0XSdG7pTuKrOmuubvXOAh8iVZHNjlvCFJToKAlCiYe5LWjl
1onROOaTqn5Ydbfw+470ZETEEkTZDThHqt5GBUe4Yt1ESuGWldLLiadoAgYSyr0o
iO3D8BHOsToD5XWBBEZhmVjTgCn/mPbSJ4beR3QRI4EqPLWhbstCLyoQsA9roLsU
wiM95HDl4GTzFCLET5EvMGU/9s/KR0g3bxj0gxWRpHu4425cArhwcyHkvNQq8xvj
v3XT9ygyGqKfvQJUsWLhKLVhnkQY7ZG0ZcRjjQBUaPvdoukSPP99uEzNa/aEO67N
GiVIh8tUnt4cyl4GQsh+kQjZ/lhESldlsw1pFBqX5kJEMQcnle+1w3blaJxA2Sf1
eixEifDjRcjuLLqpwwlhS30KieM0aF2WEIbgRMDCa5Jf+Z1YmzvaTiOvjWHs0K1B
DrtGH3qNHaAX3kaw0y1K1UDbijqu4o3VIqPNB7gvh0Axrx5KxVYwEa6G14zb+63p
ovsJwdsPSMzhyZf9F9lRu0TdsTBtIKLWQBP2smb84+wfzOf0Zk+cYFXyd1qEbceE
YRhyZtmGCGMNviFD6r5DKyX8mar8Xnngy5uw08x3wTNnN+Ep2kbj4VfMrH2arcO5
+AljjJX0gcf7I7CSQFSdYKg5OPZFWly6MW9BdDXXrGfQoGh8vZ9/8kHKsIWPxqv2
Jz/GBcb/No3OYcw5ITzkwk+82L+GU9YostVQpLjthWQi1Eo+roQtgso7MPdI2prF
qa7145ahRuRPnlFUWUG/1wmFR//EEVOfsBLo+EMAqobIXeFdjbMcvREOB4TkK4lQ
yxlk5NtltbUQaJN4/CWwfbs871XsT3rOSoX8TTv5pQEwov8w4RJCgqInke6BO0ol
F/BHuRTer+e43IlSe9EPMvhY4VnLsSb7J2oL9LcV6enLtGB2Cv7jdWR3VRoi4Q0y
mQizr1Fw265uEAliQxLdfK6SV3YnpXRhzSO+1nPqUhAz/JItASqt3gjI8NAzCjJj
ZvfW+LOfdB4mAwrR/llFFEiE0lzOLeqBvD5hDHy0GI5ebHKmn+EixktyL2QQhNgr
53iRWIjBOM40hTxwzPvWDr0K3IFL7Mu7oTNBNyMRGhvEpZptjeKaofrFwRdeEuIm
MaGvIw0FKVZZb7qXt/XIb95HU4lUzvHoeUbg63+PEqPRg61X6vJi44MllBzyQx9e
8ZjTFiEvdLE2pZJpPA8rZDJZ4O2rovH+oZjIcFjQQA2mEneFNd6m2cb4U0vOR5sg
bfGQVfJyIWqrOk1aTUoWboSpMdihM7BuS5JftgeL/HmIcrxJwzxk5CGPTDvWlXMN
heg1jQANI2RvffchJk9Ens2M0Jbp1fGLdlFQPTyLU8exjjUOAqKVppNjywaVuF+O
jDT1FA3egLAQg7XE2swe1JzzTBfP4vO2gBbQNPOcTZGbsNb0dzNvnCRGZiRKqsNc
mZbs4ql1A3DYYK8QBKsTqWoIhBAyapACMD9aQnu2HzuRjfMcyzCIGgF2i7dHq4zl
317WSNVcpuPazqkjgxhy3AZjhmKOeI3Cb09Q71NY2czR3eQnQds+k21HjvatG7pX
GMOLXVkc3pVONkgR+DeyH8/jtSF7GWSErqhZbkN5nq5M3FsCr0z8NgXPds0yPyGD
qL2sAErhA8SHeX5NIHKcibQmFQ1QrkSYhhuwHGUw1fbNCpwB/hgR45HgGZBMx6kd
g/lNQ5EhVp/BTjve3Vb4vlS2TYc/bgvvUqPRAPiaCOwm9DJYkYSdSgNqPtb6ychW
Wn5mAdU8xn8ASWA4utA4TQ4gd/MGMRNXfQJJrj7CSQ1ZA0RV5ZOOUj8qclU/5MGY
Y+zXNvDOwItBcbc/LtwaOCntxcMQWHjJ/LsYpzg6dQ9mngYcT2jti/fZuFgTLrdx
2YL5vlf2XAsRXxjg4QPKZ4y0CefD7tqOOFf8YwN9O2GYhImyPPHXMtuOEb+uyHxz
cfQZnyjjbu4C7mOg1XdEFMw54NTUuVlxbVfoK+HYg/gBHiqJT5rJ6MnIBZkID9UT
kIZbOocTkbj3+itnyzSR5k2qqt60uK3Cuj9vA7SYE+R3ifCgFq4V3rIg9qqfDvw2
QDz3F9/Nm3j6cpgwc2h8/1UrLdqNldtgn6/fs1ELMniSrICOYLP+q0vIM+jthHzv
oacT4+dwm2ojig0IN5Wrf8bGP27p62LM+41y8+T1ulLjako05ErtEiOg8ky/Ubq3
F1c0VW5cbA1I9t1TVNTvwzIsb1vLLgNAQXq3HKyV03xsV94kPC818VfRzJj3b56y
ka5X6G7EWn9qPOOfcfaex4VkfPX5VSJfJgo05Owmn71f06ONSsoRmUI/gvqf44h8
e0HoMfUie3EWXanxEA/G8j94SdpicVCQsNO4vbYMdHD4KBwvfu9CwtI9pO70mkBP
9nlqKfpNXYMVylFsIIHtDiQGtesOj4jm52llqYGX4CIWKKVGm95i4fCufKLH0H+t
BctxXFGhvjR5u5e/5JmOixTG8qrSmy2JkhIQUzTH3rG0UoNPSFVG91f8+kU1TqDx
uxeGnhhUogw5t4CvPwdgafY1bXrX4c2KDTF0gtHpmRjDipek/ouGh57Vu3hiWVK7
/x5zGvJae7bZjbTV5MggxmKJ9/qSoez/kHdIcpxNUswammZ/xMZlngTcB/NjvWnz
ooTZOy+82pDu5c58Cj6j3Zh34Q0RoyeEJraAKHkVEFRfqQsbZShvhWd+q163YkDu
mMRpCS4usrl2xaD1prpaukadBw+rTKeOS/JR7vm7dVxCF9M7UPD2oiT+jFL76A6S
lU+cxDXv5CT1xLNkhBO3xMoAvrrZ3akqGe71hFjKBvQR0szxGroMCYY8mp98esVO
czv1Kloi/RBgJP2Awd2xk5wi0mXr8Z30CFDwqFAVpcUQXAEMoDxDVG71WHNeGxDl
F2NAS3rsTUEpTWlArRlaGOhqZBUzifxL0oV9IGG6VYF8aDL+HVcys3tum/TtbC+h
0TfcQz0IGWkRnCIBIC/XTvD6YKbabaHRWuXzaqu4sPubJtaWVapRKkWBH5QMMzmp
K9xlsvz67WNZrNkrB4q097FhhgmDfg3NOpdXZD09ZLSlnvVMwufWoYLFiQHmFMfT
KRmdydOjNaA6+WeZQyaLUMXnmhnRHcsCYKVL/Th1ZYF3YCpA5qQQV/Cka+fSbKOI
qYOfgafZV3P/81dCdyb69yBUuh/CSr2AYSWCa0I7iSedivTHKtHgBHICvL+q+GH6
eJpNsEsL5a6zxSoJ6PI7cfMIwwsWQGDcbeQKiNw7exSTdUIEdfhIEWvkmPNuTAho
NOtWj1JGHTr9i9Z9ymAGbqgT8W2Rc2c8EcyXOySETp1pUoPLzZB6pPGCbVlu7HfK
wS0j0tw50StQbwPyGxKA1PDLmKpfW9jwY48o/Easb05LgyDYDkN8Er2U6Nwrg6Q6
qCWXdFT1ur069WsblaiAEgqilvDT3ScOBT7S/X9V7ghp06vhS01SmCb72YqPB49r
Ko3xtIicQeBVbRt0fmPl2SMoizJVDEshtO9Vxzj2NAp0GRWrLutWuyC5IIe0y6X2
rzf8iD8avCjTmUM9/7B/AQW1tQZ6oCBYKsnupRj4zs1mZSH+CZMhJuX1pfB8cTP9
+hNFsTEEgrPWn7Gs8bO/mV4XKsJCPMSGTn06jPOP88XPHjgZYaIF8DP3lC0ZfbXA
N1TXFj2ZRZ39ZvEO6p07TAiJQpZWF91UqosCsdtMgVtUr31pkK4Qys0NnTKr/C9v
JWasYBGp3bu61Foz5PbYRl6wpyJxnp8kFyCwHQ2MdufK8+701RH3xuxHgbZsH4Tl
brkfC5WgXtCSOe1Y65fNMmRbIFXMLT0LvAJvv9V/woC39cQUhQfyeCXO7Hwo2m8D
mVTOVZQGI9eslDlxQM8X9i3y/95Wg0QfzaANDL8lWEHP0QGXULjiHNb6dAh3X7bM
G9zZRJ4zQLXbI/SjLYFjz/NH9VAnyiKKkynIAYCpfxbRbLFsHOxKkiiuVhbRBXNy
SZoTXf0ntzZvHxMr7EKILPhexohm+9KMTexdltgpYkacr5Aj1J6H8hpBdN9uBaMi
Qm/qINLbaqLe87jovF7PLzWIs36ZVdvuvE3UMWpwjCazj20RNWEDL5ujuJ7/kRgL
AikqBqzuBvoXmO4wwCijPfMqTtsNT7iSh9qLaL8EIVFjF8KzQTyy5oQQEdzgOLl3
eHdv1gKmsp7HYCDi/3tDKqwTOmfWLIPfU0HMc9ZPA8rwwCpQAsOrxIjx22su2GCZ
ZSJzOdiO9OVLcjWi8bg4A52Ub+QzOWXDu9I3+14QyFX5J/1I3IkKd/UK95AcWfQd
UBEPB3zJRhfCZcLnRab4eNqHrCFX1PwJgiEDsWTlgPnRGlVy6RKzQPJzUWCoZ8f/
xLOFbn00OYpTXjBYOS2hU7ydEl7hSJKf/69k8vYTwMb3EkBkIg5w2msXRadYs0N2
hxXJ32LjxVoHX06Mp7ZUywg980xWtYbDjDnL/ldcEZ5BVR46g0nlRVQZm21PPX8X
wnculRGboFrKbmQJu/sC/uQ9h7vCejRRBP8Ua7Zt5YqYBt+FZKHiy7T58O+dY2Tk
0M4Pe3Pw1ImsfB1nBcV9aypIAAuvwmT1u7BX0kWblv/VjhIvBWQyp516UbPzx8QG
e1SepGl2nvL0YjGIyZ6YutId929/5EjLILaKpPnzZwzxyU/p/clzLKj1Ynwf/1iX
mwzq4rxsV4xLmM+lEGHVUubOGFV5IBBYbsRdgsHjFHn6CBpSegOrTXXGdcEALtuI
yWEvi2gpkqaPLpwY7yHJFdg5kuQ8xlwGipYAqUr5gmMh06lWojtZMrjNG3DPdmo8
zeqbjN06GCujVMoA4Ie/wcNdgdA3wWtyuLo22PdaUq0lVaH24a8K0Cx6fOr64RLc
DiYI7elWwlc+dN293fOQbLPrgWZyQRQ+ILnxoEHAk8TuOcQjuTZUAK68goMLGU7u
EhnX3beWGXpXkGPoOaR2cb+meuzpi3Dd2+lmUYunk4NL71E06sxv23fHJk3bx5cZ
nNd/GZH+so5rUFxNFhUfvIZxZNChxhnCK1+/eB24Si35nhLJKw8HyFHWUArt1rXi
30BKeAGvF/atMRt1VPS7Wzc2qmpwWtoCcdOtnGp8f//wEoo6+azzjQ2QX8nWsDiH
YgnihrUrTpYYN5wD8+yALW0OnUfd3/J2Zozp505c2cyU1pejWISSslwlQqrbMw7/
qACmpvKYJNFrcY9C//1xx92SXmOZq7/YecNSusAHY25h0XOuTuwwogD0WYKe1lXU
Vaq7QVj5BEx1xsl+8UuhBnWIwT7dyfpd4OtiSLhGKfdw9FsHKVGKLMMSBPojUg5j
8o4s1LsyErSUZ7mcmifMwT0eU0whNch5Nv/PU4FeADEHRO1O8qecNESG5OjmT4a0
jVS2kF9H3PYG1wnKCDtRX61tIaniV5EY/mRed2uX+gWJZugpASgEXiLb85pr+RT3
EwLutdhK098KsUsvKH9sKsqHxCvDb+5jvljl9taqRP5h4lu86BCF5rLXYDd/aqgx
lXWOv4l1PN9GJwRYlxZi71bSrw3G8hao+IKxwwCvpgF7HqLshbjeIRC+uAPK/Sl7
a/xem4YE6uWMvRIX5R86Y9jHnqTZB2dS8zUOZ9D4pU/wTJEj22uhtDpRAS5YFqv8
NeMFusn6B0nMykfZhie+T6GqM7UXMmU7oFWAisVokjSc4OaVVv7n1IhKuSFu7JQ+
xAdLiu/FqYAg8d4p4e2+ZDE2+1JSCqJIkgAwB5EHS2Y+L7zBflhpoImZ/EvUEv+t
WeYrKVctvktQ6au1gR+OsU8nYWd0ijjei/iWSEh48FHtNJfuaoOLIe20lFZDEEGd
hcFlFmTsbd9+JbGZ9BZB76FaNqjA2xX/G7yFNpB5YT+ohZPshwXqO8ixJ4QpsGxH
ZWlAaRxfhRZg8Xe+/Gq07ycBId6HGhaZFkUR+5n+BYh1c0DmSqvxY3Sl5KZpdCo8
bKD4FxC/lEQx9Zt1OiCPvh7vcxy+tJa1wKiBUpJy5i3ry1XoilXONMqjHXIktgzP
7OzdXqhwJfCiqxW0GHaxiqNqNbLdshEGOnggfMYX85pzHkTmsdnaS3/vB20PZGFx
3x+Ef3/UMaRASFWQ6rZmnkEGBrZrBQ6QNreix86edmf+JWNrpqpKfBWplkZSwRcJ
n+E7QGdhR5T1MlP2++22BvoxiLcxY8whi6dllofm5TnE9OB3KskQLiD9fibr5LXo
vzJhf7OnRICmdJung3B3mkbEypRLYMnnIHx+OmHkoFoEOpvjEPTYp/6dX13voRnD
7+fy7bvJbZPPpzMXIoVJzCG0Pm5YJYHxxzQeMPNOn1eeprK7MqRqf+av84C75T9/
ufhNk/0WZq+jaraX8dCAmVKhokwmXX82BAvx3tTRIuaP6wxEPOoJkcmoVj5hOqhp
QoemM+S0FcGvyFlMYcSSYXOKydvB4pe1fuonw0pWaO88266HrP9gcLauWocjI1cp
rW+i3adhEh58uqWr4/wF8XX9YtBhc+uTdKe/NibL77R0gXPJRzgxk5f2c+EQRRwO
NqSDX6lHB+lnfKXeuVomckVSvGGTKTtbZpZ5UcC4p19HKKvejRZz8fzVxdy7bRa1
Qtv5EcLhSTYLyAdUngoIPvI33Gm9Z2e9KKxMqRd6HoMt7REqMCClcCsfbK9Tm6Mf
ZLYuMO3j6E2XBNSsgroUxR0ujfN+skv7BdMhPmn/yhiLIlytaVzYvsYQRWUP4B9l
ZRoRdQFQXLV9bkRqSl3MedSfGaeSOkXhzowU//NbJnRnF4foqvV+DIs1WoUAtzSs
yatIZB/YJL2pmYxzJwfBTnoRZL9zR+Mkx35WKMBsylNY2ftc0Cmp8PqwQYyNebXn
/gdFB0OX2uyic4azG+l1SDyZd19Xl8UBcSIRYp6SOLTNvPyRWmfK8wG0BiiuS1yG
VzNcOCiCKI1cGcAM7vdrfd+dug17ULBuBc+CmWV4qLEEfw6cWm1aP354jKs8A3Bs
tpqjC7GRmRLgdBEtIU8vNBqlbK2R2pQZbtgQvFcv+JvcQOP6Oo8Tpy3YM7ZlmhFf
2U7orDHt67YQ+kZ0Zxc9sSfs40Bk3FxtjgoOvVKOIyg0w0CwXPotihRDiVcVr0b7
ivoS8ilxb2yxQBTBEPl3spjPdquKUilo0IhTdnhRMewNm5R5mdldzFlPfwndPSi6
0k4LW4deVExynEh24i6hwqoGgb23o+l4FcQJS+LlBEq1X/GpiQPcAm96+TfA25QS
hz7OFq76gwexZhi1azJCC0f1glV9OVZdEkqp6HkTLctsVdMBQsvqA7yj24xpG1mB
GQq770cxjiHqU8DxYjj5/l62DvFPHCrnapGybRmCtP1IbciN9Izk6z2CKM8uDfnO
1Gmd+NxuMX0O2CxWy+f5DLywAwzotIAhjKn3KxnkyZX6UPpE6UFH/4JNP0yT/MmG
Di0k2TU3aRqXauC63lT9niUMYTw/Q5hKGCv5NqDDbAr//kjIQSXaAoLhkirxgEPN
PVAKxsKCWRivNiAxXywrhJ1DGqFGheH5A1KuObdvti+e408ax8BphKElEmG1wh/U
7R41sD9nGQ5NLK/tDz97q1YPI8nMQntxRFHZ4K7NL7ppJPVx90zU5Rmr/dCtFAks
ByeS23dlJlDr3fvdnhvxWwpB0slyovSHKQbjZgxGB2CAprMle4zcqpVo8bX5nkC6
XrmSqlZWr/8Ohz8FA0yVgEpxc84hcWwAnJvlLwzRYXlCpZVJ4YBx7VY2k64S9XYx
T/6pBTTgZcvycmvWR9f6NjNMkFQkqDSExqvGvUzTrK0a60DTUjv6MzYmZwWuujhn
2KlXha9tf9tmGdZRfdhPEiRb3IdwEq5zZTsaHATlKXs7V1Kuunl05kCetSHukrUK
YUU/hbdrI0n03j9Lotpg8lOaJ8HjRgbP0CxWIAqkS+El9P06khwOlvdv2Dn1Tlee
p4jPQw+6KsFksS1UrgrYcK7BXflcEeOXhB8EG1bOn7QpQjM1yeembSNJEYnNNOpz
ZFTtRJaOpfkpLUPUSoNisPVCQP74cdZGHxT/UyT9Vncr0zhxXKadK79XlAyNL34T
6ZD931qMoM6hBIg19XvwXZd/VQKVZK+s68DaGavmjawH0I3AUHOMo1yv3U2MMPVL
WqXHGOK42zbweVImlMj9wF6/nDdLnTF1zTZtQiI8nKrUK2awUgOyRUDoZ5qOsc2I
fT6IKOtBAl3BQt8bLyS5ZPDYEj/pnkddREi3GrEr2K5wWzAxjUs4SlaXTICS6ZQV
7Pt3/EnZtGMBtcws/v+7jsJ0sIP4g56p43zUA7KzWz5I/zpO2kDMz7y2RXH32OTU
YytecSmmj+z3SpZHIXnC1GsHQDuwkki4cHURI36GNDSOihrC+xM6M6UEkYApaW+u
nKvWaISsaMcuKVBk+1WDNSzFOL7ms4vfguodN0UFIbVTEon1v6WAFWlmYZzWDgr/
kz45pNCjasF0AT2EC4+iCHjgj0eNEshe0vd1FfRbmPOuq71vXw1dQRfgSHWcYFmQ
o/Yhux+F+8ImQdBQfRedd2TwexB5ICA2rAum0entjVEkzLouMElF80NEa+bvw7No
xAUaarBy06d3a5hwyvGufF33VukKewrhlfIN1Y905rQN+FR7tLelDozuKRZEAqH4
3camZrlRa/lBZdlCt0gJ9ndJBiyZ+cE5NW9ogXvmP+vEL/8BaFYVHho3G44Mo7wL
z0gxpSMDjg9VHthOtPkgCjN1cVZB6uvKtoCqFg652x1t+jkj66I3WCYO1vJcZKyX
Ho67nNPNf3N9WmvugFGCz03nXpDcVS0ptt90T8Ph3xn0EYgiJa2LtptWGM5BTELP
G/lqQnnibzg5THtHy9ODH01HehxiBcym9x1E+Y4eomw1gAe9DY47xgLnoxh1p4iy
XfZOLCyAI4smIfw0XBwVmvw6xjxP/gC95OwismseWvYVcXRjRghB0RAOD5Wy0A84
+rKaO6AJxcwY+fgYqe8wB1QyLK9zJBLkFSv6OOjer590RLPrbs0q6W81Ei7uLsf2
ecYcGuN6NKJhLos69qtUF9WHXtLqSPINfKuWI+5Y1HTzmsV1crwdSSGF8ugFUMiX
I/vXW2oJrrUMN+Z9N8SAuD4M0e+/poM2IizAglp2DrMZbk6AnbYCyCkasdsZRAyJ
vn/4wxa/b7PMQdg8LBM6IAxS9kLRUNP6NiDnamXJva9cwRlPmHXgODjpz8y+Rs8c
jT+cEgH5uhh3yJISSoI1uloiT8zdpAuypFFgnoA7AEHn0s0LHQMqsAnpY2MQKQ/k
IdUTf30b8dl5lWJRyTDf6RkLWQYJ5sEOYfRd9aC4epOPJjeawTDCQ8UhoM3QEUPS
HyphKNCrK2cGT3YfrMppyacZRD5/hpTN8FJkpILkM2V5zFrIFOJg5NqHQ01YSGjV
/PRRplNZ4ZSwh/GER+nLoeEqML5rXY3z5kYqn+A5NQ7VDymlrFq6vTupEAWz+vJx
nUNewIyww+a+dDHfHzIrgUucUTErSxyPyS+qu13DjcF5qLdnfau75oJ5FePR4vb/
pF3YfVwkguKHErtb1rqceoRpQuYrlTUrLxzmVMtdN56wIuYXiCeGQumvbX7WNEHN
BtG+yG2M8diKlfUwD5waMPyDGG7Ut4zhH0xXeKrD2Bgw2M9ID/61COOC/yq+hlaE
nz4bqL54F2nj/QQyNjO5HJyq/4DrWUuxU9cZGxM577+Ajbs9iHC416UU5WxSuZ9g
dhP+RaiPfk5acCuAMX1bLCShKHTtRbj5CytBTvtFKXEjdQhtDM6oguvx2uyM0LvN
S6t9xEigwC+FraScW2orEM3s1PIzGUi7vjaa+FOUXmylFcXi+0TuBEtd0J2JoYEc
vDTIYRmFBcc+M+8+vqR841M1I3SvDRl1OeNeC2VSV65Qme8qbipgH3TOQo5r6OFK
XDYwM9UIrGqi2p06/C3NGm3KaokKVR5A7ALEzgULvTPgZq34YKlGWILHEd57sUkH
2ObuPy5+HtoyrxzHtR/DGpKD59ZbXHzMbIpuSoM6Xvmwdr+KNhRT2zxsKOIg1sfA
S2Nyo7qY1ZIO/YnmYMN7Nn/VuzQ9GyfbmC6drPySzM+W9TSJyDylkF4nklBV4T7q
+B4aTPwuCbNsHbqwFeMZfTPWuQ0OdEgP3rav61gL2gwDJMg4nsBHBif1hsL6dSsg
8H4AZwB3shgC2Bb5jFCN7Mq01iiyDjoP6J0na0/1eqgPNHvHqbwPVA68F7XZn0/G
l4sprmXMnSknnCkzsJgpwdqZIVt8QoLoNk2uVZeF+L4MnZWmhRmUpij8tiPnW3K7
USG4RgwYD0fC6H+5YHpHkEueLCIqHRVkQfhEO7PClzSTQaCig9yq3XiMT67k5BJq
4OGlLDJRhsedFeUuxszqNWbiPEINtMTsPUB/rSlJTZiKRC6REfehSm3IPWsULQOx
VT9HSQPKChWRsef/bV2Esm0nDPqwtaNjYvqoqwGb5ZxVPlmnHCZ3EprYEWPWnH8E
+4ax9DbdI57Wa8ZyAsGszy7vAqa60w37Y8WtAxPSi9K6aPQaBalBEbT8SKHnvyl2
+88aGPo6iohO/eW/Cvgo8y5wfQoZLzTe7PIQsLcKVXN92MUvYPOWcdkN0DFEBSD4
A/128KHrP2k1lIeTe8JaC9Un+loADnE8Og+OEJokHHkIBQ1KtT1/TSys1orG7uhj
10YsAv6hjnELLT8af2k2F51rWlhAkZ3yEU33XiZO1e/+FMWFgkOtjMpSoxrxjd9x
lqkQ8HUr7IgtyHBNBulmFVskF/3SVO2bzT13fJriPq5N2H9CUr8j6WqeWiwqTCgv
o678f0S6bXW5ErJDIHbuAJRcpXAXd29euFoKdzxBtZQijp3O8NvYVgF/FzJbIi6a
QyxqVLdZHYcMi7j3TMNmY66aA6OcmnYnC8/2g36nOJDfetsoEbBGaIrpp6zm2igg
2zJuusKlZlZifDoRMpJImzrk0lLMPZppUVwGtNUNxzVZzSfB956kI76BauGckPgc
i0rVD5hUShmvnu6CUjZas9hbIo8hfJfSuVSqNu+B6E3/zE3jnufKXbZg5+tHMjKz
QsgA69js08zz/P1Dy5i92P15IwAS6zbG/key/k2QB6KZn34hHeotgigwXK3I9U9V
OGeaFlm3E9ppBaWKxqkFXoiOm3Rpg30L5ynJiHSq2eaRfpaGRnjFHg2uwUBYWJBh
W+BsopMgRtUYmF/EjPfgQBLq541AU2Z2/fxuM48H3svOO4Z/tb8OYyoAyxouHxMQ
DLCDu6MCcMn+x+F+BwAfuhOwUJFb+4Q7eILSt5CBBM2tUfgQvlanxJXHilzgFYor
xCwB939zv19yiE4BRJGXNb+12EIufjR+ZH+/gLzMRepoZnaQkMgEpMYLT5mk63sM
MIf7c1H++WcMD8yV7frDFDTFDlteG0p+69NdfFqlzTWUG9Vh4fa5OS42fNEqle0/
NOH4d7XfnLy/7mdwlyTpzhOQHqKIjMzGVD42lxZFbKD+e45g2LUKyRSAoDnXQQVR
FUNr8sNom4HeRHaPfLW6LQ5K2wFKq2wJSjdVr978ZHtL5/S82JqT4bihVSyiy5Ud
ICtlR2SwG/1/5sx4ZkaKREHVejaPWlhi+u3LiENHKTpnxXoKi7KQB7y/VhWguxgx
dZBWs22nTqZ83QiOtK9pJwcXTjzHQ5TCNc43YxoRN+xz30aaF4PuW3tWOYadU6iU
Fapy5DzPJpehjrTtbHj//0yjfzr0tvxm5WggYng5nY+tCc9b0tSJi4D5GnO0rerb
GNTT1PRPi5QVnfTKKeSOh80druaVvv9Gjx2Dy/iGpIQhjIllzs7wF8JyWJFHx8OD
z7NouNTdfZFMQhkeP1BFWXXHqbfzvnw2jwUUIZLn976T68CNkA+Ip5rb0j8XYPhR
MXO1aV1Bfs6KyQkp+tbl7yXjePc85rO+AYYCT+sfHxwtR84nL9+/EEHtErl1kPcV
c1HlcOQ2sSJkCzG0dR4KGD/mpX6/NoxUJz6fcdZ78+5QLQlsq1jY+Ows+6rSjo67
/iQDKgK/8uvlEP7v1EEVWLxqkNIKWto3Q1m1sF/0cKgHG9C1bsLI932+KUeS2ESQ
UnGpqINHr8YnVXJ5Lum4uqiFUcB/rvNFC4FZDkjnjLbh/mn6fjL5UcRxQqeyhuYh
/GB98JyPw9ZonOMNxmUVH7iz+6TuMSPFznjY/UgcJ0PxMtL3azZG5kdnBibbdX7o
WZXJtOgClPFP9huFWJzdY1WCRMS4fbFHIxTeilqXsV81aXCiPPFfLRmi2PJHCSTN
8OlsC1KkI9a9x2F5FX1sTY9XtK8X/0uJGXO5awI4VO+k76Ifa8dzAypBePItIt/W
OccON5CWPaSpYjidpU7l+3NnG4CW7xR584bA2biJDkscT2tcdVh72+FWIrmZasyi
cxLu88kTU6mkTkxouO5lTxFw+FPPcjWLIpQ/1KwkKmTiSzxNEg81jzwqpbagAZpN
HzVO5esnLqUYBYI+jCe9kVZ+6MgkkC3tz4ygWCZUCIWmUMsXm+4TDvZDb07UgQLx
gykjtE3Pcv9G5kznwWIjEWbkbQiSsm97V7ar4xe0ZBtMhbaC6wsDeEaPeRfbYACR
elRUxWraA/0P2e4M0msMydDAPJ782ZrDO3S1k7nD+BPkEIQTuo9Z3MQ6C2yclZNF
0nPPiottO/jfNzDpyJRrHldDSADfWWK9ZfqeeaWYeBCcLcAT5EwiQcXB1e4LLYw5
gTPGnEougO85BYM2j9WT8l73csIU8I3AbQmCvgdiDz0WAv2y3JDLyC4diOfDrCL6
dCZM92e9HBkWy7DwoMwuxjiUvisuSsh/owSN/4JlSL2G2gt8horBcjM8KnyA/CYs
YH3ZQdXMchd6qgcKN8DujeRa23cnk2tNJf41b9VLYnMisVeqExjN7sETTLIoDJ6D
w8QshjplriTnr7n6Dg63gH2ItojE/8pt9SwOli394BSEnSc7dl6okiWEZQirJBB0
gK8XApLd2XVcwyAiwmgKphIhwVqGbL+CeYr3wNwnWvVF2ZVoaPLH0xDHU/w8XQ3/
t5H/2dmF9oKmyb1bCW8V70IjBFZHToaAA7sTmnr52y+nGmLZXxh2b5LduuV6uKfC
fhGPmf3a3X8Je8awExKlOlIEjeUMOUsdoE/Q13xVsBiXs21jF5DVME82WAjJMoKb
Zmn2SuQ+EcUGhJ5HPd0IibsP6G26Yrqbr2e0R0aVOIjRw7JQo5MRGTlhsPm/3RfK
qfDO0IQM7psT2rmZFSFNZWwO94W/odxwObVxhG72PUNGuRegj5fn/mjCGgetrtIk
xMdlHPYIBCBdCm/6saPMmwWB/+gvN+o2zu5kKdfRxvEg5siEOVKbqT7HOaP5eJJL
9TqBUOZYmBvBjvdItxLpuBF3pjC+hcbtUdLxqvZYL7G4zvcjnkdGXDeO0a9f6gfz
wnz0MiQvwnNjLmSKRWVYxcAV3cQyxdH5QOFaRM0nG7p4sj6adBhgUSdZb166rBla
vSd/K66uHwCFwaQZ1+9nRmS+HNf/GjEzCRypJOcr4gmKvAbLm7e/owA73RbWMRCk
h8f64yQMfPw1sq5Xq8jQ+VBiRHstU6FKPQ2L2GOQ42T681z1SszKSZsZfayM/zoz
hL46dMkC9hhmhQ0R7f4HsVr+xPfKWKzmezsk9r9DxTCIT5eu8PDpTfqPyZJcLlpb
a4Zc5X5e9XuJvjOf/cfP1X50Ob8ljHd4yr1lEv2KvlvV+C3UTcTdbZ5YIu6mKxhF
/vxidRz/aBU8i+ECf77slLhdpLUtgqjXf6bsCDWj2lNY7ubPqT4dFgJwakRO3qsw
qGX0YVWGlWAqg1wJPV3b8dA8yQtFPscrUZFVr/or1+jXoKID07WXgzs76fRUgxJx
ExIpG7LQ9Vf9EKtciPIxTxJo5sfimj6L+I0XNTT2jiJNApKTcOE7Xs/dkcOsZVnV
ofvkWCVcpztxov8gmOkdIXpSN2GzXNMW6ZT2VE8jtg5NNQMTYTCqfUo6eojelHly
EjrZB2w/oPBVMKWRVna6p+qktCMiyyDp03JHO8Vl1a4Xxerc7RPWPyuW/DBZZL3O
eKzj9QYynanfwEWDpt3nPHn5Z+QH8QKOTu4qB2yobYwf6mWmCx+2paK0l4adxQWQ
l9uoeSZHkf9ISEgJorFeP2/F5aY6d3z1plursBWZu167TeFc2MwdyebWZN+gkk90
kny7gtEiek37bnizCjHP/2R2z0qulSlZfC57EV+DpuWuufHxt/KmFJyzc6sG4SsP
pOzwsU3VaRJXF8w/mH0ujZbLf+txYGyYIlNtkBBhnrvFdVFFGg4EUNFQ++H0ZBge
La/BFcPkIFCUoO9KYlKAnvT+9lCkzRKqTp64/+8RnKMlv/DY/ZvqESDsUXP6UUkC
DXgcClngDL1QjN7UrsP7t9DiyFvYV3d090qp8vbwg4CeE4fF+Ital5HeuM7YGyDC
MMWUi4EKe/zzXqkDE0YPs0D5tJj4GwmluDyxXgcaODiZ2dbovPwNISRN4n37uKOo
IhUPUD4CJ3jrIHyQytDL+6OKVt3IO3m+pUHipuKqW2m7xRfazjfm8qFWg+pk7IsZ
gqtCM2cUzxblqdb7Lva17F/xpyq8HJ5GvLkB5fIX5gQmtj2EaxtP0OPyZImFngq9
in/O5/Ye9U//Kjr6P1DGzCMrYpyAdAZD+9XTZu2q6Mw1Mg2sy0g5T+L6bzuwplQ6
n8XYgsWWzRewGA5TTSwCcaPulVj5o/kJ6H5LbbCDVk4ZQgQc8KLpaRTz4XQ6fIlB
V5K1Ug982ZJTjV2TACgVZHZVZzMsySMOSpzYcTztcnuuwK3Tu9nEZiHp76Kwv0en
40DicZ0z19/kRyVy0Lt9ta3nB1CSUT1EGlnFULJ+Pz3LWLpU+iGK7eLUUMy81x9A
QyUSu9bOQjAkt0yT0kRLNSe2w1qswI3DDcKnOLUYp1G//JLs+89JzMUYp2cCVMr2
bm/092Q2ASnRUHoKghE40PEmOv4jpxHFmHBOqZRIp7niiutMQLMQ01C5buFdL9o4
pmsmQSqh7IlyG71KY5HLzGdQnMAYg4AweMtBnymine7YP7iNDBpPch72wCf2f9C9
VoXr6KKcY0hQX1eCl1nygpFu7SiR+StM51vQxh9O5OwBep4QutttRikjcJ3AZPKb
X8UtVMjBHwIzLy454tHSbq05AdQuXyWLefJqAdcBHRab35n54nrK2Hj4itnEM7rp
RATwdMXGhcsHXR8VFC3kPMGX+q6M3MVCzATUIfhd57xlKnpxKMbW1g/XpDIvMUNS
1/RBEvrv26SUFDraWKi6B9bES5hpVgjob5DXG4k9BmeRmHYxZ1ZyQr/gD8HtMsBR
vH3Ko7EbliJuS9FKjq153e4D9fNvIXMutv4KUXh1OSoENDgHH6I/fogBn5zrwIVt
QTk/gJlnUNnsIwiddc+3U73RbQl6iDnJxYoYBjc5hY0b4BZVCrC/LE6RujHCB9vB
WzorzbF38jHf2EcUERuwJ4GuOkncAHuGIPKXCZdZTF9HN3T7YTrbrqZJELK88kIW
zWGrZrvaDLPZ22Rm0DcEV2KE5KjGOkhUp2PctQVrsSUfBo2VK1RB1Mxdxhjwnbpe
EcWln4oEWDTF1eMXkHSUj4H47k4FhSZfr2LpWfSfWYDR6mA0czyf4f8g5KUPfqEh
D2NMVJ20WI+xNdrQcfVzuPWAy15Y9aJ6zhSOdJtfrzxX5mYF5kpT7K4ERQUV4CPn
QDpqPu95zRRVsu2PljuuteO72pg98PzyPfF25D9ePQBfya6r3PzhZFJYbaZVljOp
U1Ze3LlyGNLld52hpnlZuo7mhfqkmmoAiCrvLL6MzcGe5GeRID0hpPNWMLPqjKR4
CHjlBa723vMWgSvCHCi4QjSdf9xDdvrhQkYtkyg3w86cYHmhhY7wSbABS9FvlBgw
vf3mljP9lbA2mSBGC66G3RX2TrBaRNAis+HnVv6rqEG4uUgPhoSrdflvt2ApsOr3
7VSIlGa28PQAeqaynyWWQ/TG2LG8gK3+iZgXQLCbrAFEDPT4M7nPNVopU1G2G9ou
Awc9EvYnkdjzAR9z5tJc0fEmk7ZdYVZLZLThyKqlKS1dr9qCHthOvxO7sTS8t/N8
Ls0fGeQ7XHTodLunwMaMSrUQXsHpvrVOqXSAkEQeekICJuBGr7zGRqpVeHOLigXY
R+S2PdexA9XhD3iLAn6QOxKcdO6N5VodpNhRZtYs1gZLZ9nHLJDSmqTlYoBqoixg
Du9PTkxTP7Ykrf+/zbC/aqD37uwS0cPKxurxQmLIG1h3sxApKDoI1ims3DYDHNWN
31fwNUc4eS6l71lPNOakvMv5Dgj5TScZqKtc4berBsxiSutuC4Ui2FaXZfOWu3xR
Csp6yl9qBTAlG4vH8ygoR5S1lBO2DZn6ijmQRhsXKId3s81BS1LBohzv8GdQMpt6
YUU8R/RyopzU5J9ivxqzUZK3+wI68U8DSD6WeP4nyryM38SJC+CpkzT5e2rtcQpW
D9P6xSp92nfRbX0hfcLLGSOv560YqXt3MDrVEkoiF8QkpHpGI5j4XAv2f9YqXF25
inE4X/7wZdfSwrudbmue7bF7f8xGXDE0iNUGrx96ZARBsAdKjWStB/oQDOZS4HqU
ZBSPtohgOolj8bfEGbSeIhyJRvEAKAAExDGNLCo08pKK5Vn/i3emTYjMDJIKdiGv
b8jvXyoVLghL1rA7xp6dBK9dnVAqA45qoRHANYe1KevawtUCCah37BPIKjneyX/b
6jZajWFXhre6Bcbb/TVLXksv/TpdILuOXFJyneW5x4tz3VhTcYdP1shSu4yRUhI+
3WVco3URWNCcm6uVuQNYyyaCwLz2UqIMSKMqGaV5H25VCn1BUiTxzT5li5r6USGi
HgNMf4u6xNcHVKxHd8pQxMS06Bhj/54iST74LqbJl5+xQNbGnBGMM+MdGhqWcHoh
zzoK314RQ3CCzfPZHmaQjhvZ5yC7gdsMhR1eRdWQRGkoroYAIppZbAhKhxTcAXYc
TMXjfNBt6O0U3SwPU1wyvDmtYNVtce2p6I6dMVrEstSBK6RPhqe7WT7Ke5OkwQGO
5IMnXpfmsZKz/EoGwKpVLJg3lYcpdef4wKtnsSTvbIDw+J6j3/eQY9t8zz09UWTY
ehJvjuld7lHEBCNPzPG4oykJ8rmfJ1aVuSnCTCuySvJK544L2Qe9MXrvRrayIWjd
SA/xh/K8eiTXi0yoWY7qauocqmNMyDfdnS6ETQWiWV9GvPY5K+T7AysKVv2ebQfv
x5Whxm/hSdanrYMzIB8pG+rS+isVWHsAYyi9UN6u9aHIS/dIDKJIRmmaCMXKcZC/
Gge8a9x9krXNx0xpy68NZMuLNm+5JMNyngwnNbRaRkpKG89G2qWQhaluARbFK7A9
LgDpVAPQjZLuJ9h5soL+0MDT1VZna7N0ZNk+XJjWqjjNrkRg9CkPNbBFAFWh6gII
dYbRFhz9HFvQKq+uBSeA1MjMrnb+mJCjiPG2vB+WWni8fVBDGDvPT8rezpqbSVAz
+h+jDzJJqCPFqhgTWu1WnBU9TnC3BhcQ6X3wX7ad9RJl4n3o+QdwBs132dka24A9
1FXdFx3PM0Bzh7s1WxsUTsBsjJ4EUBWKuNwA+d6c4bniEFYJRx8rTM6uvqeZn2QZ
54V5LLuB8m48Uag+4O0Az1olSrc5qq99lbttXIjuzspqgTxqdqlqBxvguPf8lxpp
aCPJ2H6bEaOmsPKZdIxkBR6Ulb4PWOocp8h6TT8v4ERMBDgs0kMSFyOVg4O1wF2f
0tAJtpXqvTbHXpZCbReCRI+VCYMmbmckAoQSseErDV9LQ3YH2XceBrWzuFx0Amfo
RtGVZx31yEwrBhodKNI5SQIfEW7I2YzATqw0xb41i0y0kQpw1b/9+HgeHJ0s4kSL
e9SoG2izHskRktAkhZiChZ8rjylFN3pJMfxvus30mYgBvH2dBb7P/BQgh5ct56vA
OYE9tnwe6pX7uccEB8ZcqQYu7s/VyDiWqdaTqkAB3AJPl5XT9Lo6d1WJIMu79q7k
6QbWdgnCsElLDBYIsqRLJnqP7d+U+WLjD73rOT4wxZA5vNIIEfIbxe7ODDvvsBu7
Jz5B3eoi/LCJHfQjvfS1blEtaVG7GdpLoLGEGA8fsC8bITEoWPeKxRsQKiQvB0bd
Ji9mIU4iZR/o7H+zfpBY5LgcOdCREwtkes4fUxUUfXNr6ukYgccyn6QMh2IMvqgr
1y6voiZoiGhoQQx7ajOMs6nfMJg02D0FjQheWATGKiB1Yx/a4WsxiwEsKtAA9CJ5
+iQV+g6ESC5Q0MEfE0W3CN3cR0OEW2unPmqhc8S4EKfTVHaFBJKiGyTMhoje7vWT
otlP30p+UqPGX32pIzZ3NYgB8iTwDeG7SQXoMLZIanhQP8N2DlsJgFUIwi0x4KsI
+g8CWuPPjOmCmijfd/54v0hOcmVr2FOuK8+hVAlwUimh52k7LRRIdEtYN6ytlFwe
f6vgYdKDC6/9ArXlxNLumP09rAX2T2xeAuRaSduHAawRlyfdAUFA8pCOf4HqzyWG
EouG3QqeJ6t0bygpSddOBQKcjtmIHVu3bea2ipf6RsxD4S0Ic+bxBH1jGEb3x3dm
2ooE3ouLQv1S2CR0mQa3MSg2IYQhBkJ3l63HaTaab5N5/8GUiOEvaCoPdL9FFvXk
vT4fj6miDVLso/WngZwd1oLS6puTPJNLptWKzpTOuqHuXQi6JAf1CGG/9EZ2tul2
8Xzm4JVJJC6OHA+gr5oOEV0CCd/YOptlu0E7NYilvTV7v83uhKrKvZKm0aLxyEUw
luIOCT9eXB0fUGr8HjrnNAbXBMctXIi+YaidkX/cHh3sKlF0vkICS5jAjnjLnVZe
OWrbrJI+4nBP6GupxhA7XlOdPr2OWR8E0SiDMU0bCeHqjeklMWgSWN3FkIaK4pqz
elxiH+d6tTMlZmtA6dmnOteaXFSn7NnSL8Yl3F06ynGmapMXdcu0D9KBdnJSKsaI
1NLPmXshcBc5BOdEiMSwIyNGiRLydKPNhsABe6r1isscq1G+V5TLPHeQ1yIm+9Dn
5JFovokf0WRfqz7+HW8vj6v7L+5a+LKWnoTYKwwOle0oizBrM152qvoyXVMshh4a
1mNEDyzB/oIjOczzUL3QFEFikmQ+lCocNgzAL2Hb4XgRYk6rWE8i0x8RmQIwS+p6
Q1H4VdVoohQiLh08ytlTq4iv0qsbjdd+puSuP8590/7wdnYemszEFrToDw8yI3H9
8ohN4Sz1BftbS8C9IWNOABcCORuefotfeATdaSw6WrAwMjoptRjjbFMMudqYulGQ
jl9rX27EgxjLyHGszhjUaIgjqqknRbgfPbJBcSoIFgEnXQFYoQP1R9IuY8KFgOEA
kd1KeFGIgg82C1RYm7Emnv5LpGWfrH1OTCQ8gD9dlGPi/RQvgWGusDPsipU/RwZp
FagDYEOEZediw4wxsdUBbuHVW1vh9Zz0b2FmSIsThD46DyOfgFiu1t4P1YNyG2oX
2NONiU8Cjh3P6EC+ZCk9lmlWO9mlIR3dmbQKzpdECKnO+oqI2U8gIqmnWVi9fKd/
kXe5Hw/y+rWCHTwtQmkcHhJZZcGsm31Xh0jR8U7krEi425bfC5ofs43d0jlvtHOl
5YNi+0XANnDFt3ZRYOhwE8PAa95GOaJvDI9wJnpnNNcgD7jzeK3t5O9z8dAVNt8Q
15o55NPO8rBv2+ZKtw6S8ynGsGSqzSLZJtpsYkXPxGNXWbZe3df244Ch4x32Q17k
Z91qpLx5//J5fQ0eM1r2akr/PZe0/zhugy2HBMHI226DVMsmjlJPwIRxn69ZHctS
8rAbp0pZViPNFRIaZ/vNhmlbExUd5Hq8eP0yD/ojnGW0rHOLTwPnE68n9bzyr+oj
XbjZJEQsWRrJLrT9DE1chNbGtZ96bcWPSxzNdiYol2Z86IL+T/2iDqVRBPIm3D9W
4l5iL6j1HZuZbSqtChKMNjDWMZt5FVJEbjmN5L4Oim52SjgOIP+cesXMO1oQ+uTu
EONHq9CtKVA+xCm5XHDSihWiodKPaa/g+8QK+2jQJK6br1HdMRkbQsdxdcM+thvb
01pX60Bm2oVIBPYOd/0pCzlFvn39RCMbx37R+3caaWr2ec4USBXE05n8qlDnwbEL
S2UkBsjxJzBYWYzFE3y2PFVtQLnF+9ri1do1trPeOJewa1Ej/IHTEa+D5vwNg0em
8bZ/b5TZ+zr6DbS8GcS2HKwIIig/RmLHF3h/rLhoYwakD5hiqAGz48rX68BeenKQ
D2HkjokBEaoOA8UE4tCNpA15JXgfzwPXN5fjOhPAw7KB4zaq95zaDTR+f8fQhrF2
GJXrgdqMmAYxpMFWc8SGBxngkWccvOY4kjNx+Nl1VuqU8BNucoB5031+++n7Vxvj
FhaqkhNQjBwjfk8vMgLzKZvkocrFQ2ZQFuWGF30ikvqeuSqVhmB+ed6ukGiZy6vg
zY6JEPCgqmQ/6biR0hZhfIPVV3p6AKvK7EeWj5OhJbrx95SAubwqbpEPFGZOXnMW
FvlSjH0ZVwH1qFy7FZlGgfmfsJzbGrCCnWEsMuIW984E/8yi/2OvhwlHzQZlr/rk
H0nC1QeLaWWi/7/ZiOft3C64FG4M8IwK/ohJ6hmrfZDzPDk70jGZIhg7y7Mr8flB
bYrYDz8HW4srYa1z8u0wxATsbs3Cbu/IcSxhp0DtUekioe6mMyWxjNiF6JAuM7Mm
UtSqRPrRcvX1nFmZOWwegbArEY5WX4OBZNnKu9DMwKuebztCDIQG14t0iIWwiFYN
gzwCMZps5800/WksFHJZUEwh3rAwx4Mdr6DmlWTXbftsuyQi3u0815cpsrZBK0+V
5k/1cAbxRSDVjLJIi7bcV4PpugboH5N4uxz60byxzrv5PV2YugjID9ME7Kwoyz6r
MkaeAiAq0VS6/Wne6HVc3snSZu3HOaDXNoBlelDyY4ZTN54JJvpUgRJdH7PlOeyH
frJfRvA1KC7rjSKI27lOcrdeaV57+Foe3eX/w4bfTX/Rb4TobDS/hzUDZTLCp0pe
nGAXVwWdQtcmt4tlTfdzY16VTKnFUTCQ+S3r1DD4hvPq+vdBN2lxYMMmTZXjNkTm
X7eqRo4ikJiraCbK3tlU0cZGsaGM6cR48kzgvC1HTNhBNbfQYoHZF+VGS5pRvfMX
x6vIaxoFZUAwXg3BJD/j0tLpbovzMDfV1VLORDWdip+ndTFFTIV+zYSA0dYsDTdy
rTvTOgskICE26x/k9eni/gJXnD70Ktimc5JobAptWm1ow3qvGBpTEIqitgBX1BKe
2FhdlcXotTdj3U/kQ11RtNALj8vxTCf26SugyggRfqfOgnC2qAKeMhEmEX10KNQa
uAQg8cKgufYyPQSoIWCDL1LHcgZ7RB7NYpaZCZm7Pr5WyAza5wg2qKSkAP/ITChJ
C7cxXh1d8SQLB9IRmZq/KUqgsDU10kBA9rB/2wZwt3ndlpUlXaIH1WZpczZYledP
maAn1fE2ncB1mveEiLyo8kvThOPOHNUkXqOYJpdTzIq4YOZtT0lq62WQ8dYJdM8V
oQ5bo7SGDyomI97Vs3Q06Nq/t4unevyh6Sr71722YoqbKhgzYI5m6yfghcYuoMXB
AkIPttgkficxG69HSWSSab2o5563xpNAldQX6V7NQ/ADVMHaycHnNiJULSN98UwX
FGchtAxoD3I+td6/ea0EaDZ80E/xGHFyRk/CEtwL1yKJNBketU1P8+7tPUnydYJK
QXanLTu1FqeBRv3pgHuCe5x2mil46dYtHyUbB1YqOjho5SI3u0MT9HiwR15hBH2x
i5A/81GXhexoU0Qjw2EvxfgBp87rtty52qayOmQ+EXphDa2uvNPdnWmwctt8uNjL
TjbYFDbln/nmKDCHr9T9oYFMbWFrCpxmPfQzrOYhCqsTW7iiLueA+qUjyGxgTget
1fU1GWst/OuHSzWngksXvKAOzzJmb1r3/1C9LeerBYeoddUb5hFjhXT7HgMizFfm
HtfM1PwXRbRM+MVg5y516aTUYnzuxKGYGJFT34bjj0VxFfpw0aI+L/2vLaeTb1b7
lWCovZIEm/4XfWvvoRjjypadpaJFqJi0u70H+T4QwJfrE1Vj7RR8vj0rLhORcA/F
8OPMlaobmiTi6JaUpGVgsLiJcUq4AVUfi2YlptTvdDegd1kH/VQqfocs2HY/HyFQ
yoNSB8sFDhoKZq5ssk9mkpuI2rCLSWMEYR17ryuQhSx2zV7DXPKqoG6SViy5BH15
TRlj1gIlRYmW7nRiadOvRiaNdSs1bfWgdAytqbzWfdcKdO0GbWAbBZ8u5LBY4OaV
qBLQHL3ZE28wz1QoAFHIB+TZBxHhnEPGOl4pQ0MVRlwuyFiKiNCxV4mWueQ5tDns
F/8WoN7NHemHeNHagYh9FWyzdqGtaOabs5RFUlxKct4RfX+fY7oJ0Mx4tasTSJzJ
+tApXYOlN3DPhbtBZUx8GEIYjcBu75PY7JSstRksSo7JsHibvwAq+DkvLIli+SeG
krqpoPllIGXjE5lXxrEXsS4+4ZR3XnZpC0e1cKD7DJDU0HlVvjnQNtT4EM42kSkW
LwSJ9RSQagvtvYkH6QWgZoDQSPeSwZjigGavnme5oAHhSGJiiUB5OItsB3afuEy7
Ljkp4pRPYdRVGUKOZnucv+/vH3mh2rTN7sR0YVpu/H3HBWpk9esgbmGjHsDaNeLq
j+wQHAarQXHFbHMxPzjvqirkKlhIDoTuPO0raZdmwL2Wfadzwgg3A6qhQGJulMKO
SzhQsy8QyyA7hPzZnelDUwb90tYJN46tZIPOKp7FkzI/lpS2pFPk5UvikhgCQI+U
HYIK+OArp+zJsUb9JMsqq54Gw/4ki/hdwb4xBXfIHxMZq2mlwnWkH56oYHVJ3j6H
QLIdPofpWyLwKxEYJfHVYW4Lge/uQb/yL1aiGaAqoA5yfsrUV02o9jD3thvSIX8c
6DsW4dDaNWmu8c1vNpnisrFJ3H+c1l0q610CNhLgI1/68KsJLmJn1UnpwHiZbM06
Rx0LidXS55KzDCeIFGvn+sZOF3TPLa0tkc3C5pySctnLh4T4dURNAFF93m3GEHdJ
u6Ng9lbypFZj0u4LMVtSE2YIaXyVR+wxCNl40u4Gd8kGKXzJOFOP+HhWsiQ12RV+
puvGQCBX0XvSsoGcnoRy0oGDwRNZjIr5DOcUOHcFLt8ZeOpQzsaCbXa5LhWvuowB
CCLZ5zPccs7BQRWqp/t7AY478JZHirPOLnVA1YcSR038ISZjhnblIJZG2e/PV3Sy
oW4STBaWu/cBC78k3RLcsOtrioaGwbjTeAAj8qsOqKd/YsUErV8KUALH+j2qKE5Q
n/Uz5FFr60OsFMVffRRnzgBgCZdnMepAzrjjjEORGfwp62ej6rDhPpxqIRJ/i6OS
mLoFqE5a3vWxFZXKsWwNaFQttqerBnwTwTt5GMUl1SOHFeR5oLwp/+uPmJ1Heq/y
eFB4qHoOwuxFdwhptvM0EThVpFo+zbW/ZaemZC+UQ9XWV2vvZzkOC4hd6Md3XxT6
iTXxTgveN6fSMe9s/SpIY9osxWcioEPS+f8ocgDjuSQLHo1dMcicxyViaLcb6Vt2
poxxzccGTtlohwDFCWCW4BsV9/ZMyhsNXBB2Re5Jc7MtiXfCZSVo/G5lxu1STSLM
kIjZ9nCc/FdS5ofW9WhXZL032FCbsEhhPLYUq0SuXlYhzy35h2JSm7xVy/hDwq8J
A8Y82qvaqk20ey7SULlsfIG2mEzTIY9qAImpAGkiwMAUFmf7uUdXP/Pt65G/jIzk
WOV7wxBO9nySo1oU0NfSAVN8G26kuRKU5+bVDd8NQ7ZsNtCuaWkzOvS8TVqlTGa7
XQfX7pHq4ZVSCcnNz/M41poBqfh58XesH2Q6uKjv22NaDUg93aBrBxK356J0HYB0
0QSBwETZKK9KR/t52Q0w2WSjPosUmXYIeYRkPno9qXvsD3F+S7LSws6tByOxFMr7
8Y8kPLybGaL7w01NPMdQVlwWpd6CAC9koWVkXo3Iha3Fca16d6uNltKgnCJ+dna2
bhz5rDA8B6qphI3IMFA27y6kPu701hsY1Mo/nZVewy4vIFzc1HvDvOh0HeTMxs7B
uuJuosaQmGcAvYhjtEXTpxWLN0wWh+3T0EGVyKIZbyXgobxJwAzMZXrkdQZjKwTM
x0DxPNowuxWZl9YtSnD+dKsClyt/6ZGwVVsvgWU+jQl5sFCFF6EPNS+eIqE6arF2
crU6k40/b9b7RuiDw9Oh0HYwA0hHnuT6QgLS3qTg0KBSptqDu9cJoG9K4yjVAUvC
JLV0/IoqJupN+4Q8Va7linakjm/fpH2/HE61AvOjnsk73j74gpBhCGZC3JdVVTGj
EiDFJ8meF08GJgESQVl32kf6L4vk+qel4qhjDtgJ9pXDicIKV9PWLcTcLBiK/B0r
7PoN7qWCNyJuobhpkPtrfakN6AU5y81WaVBH9iDaR5sUrBwLwEhVwTrUX1w6D3v2
1mxrlBldnLwgIUz5gGzQbJKbRDc93tfak7O0D07hpuvbab19XnJ4vY30dleo5kwT
FRS+bGCOnHuwUnUTaSZkl73SlNbjP9Dp7EMlMc7U8EIKuaHvk+iixeQm5pe3NXd8
ncUXlk9hVFb5fzdmVV4wkDw20fUxnt1b7VjTKKlBCneZdShrEm1KIMZcavj2xtiz
/b2RDndz87V+OaVG6eu4pX1BCTi5SEucZA/3QWiwQS3ts9QJr7T7KCZehhowxaB3
hKuBDaXTbaSy0RYqf1hkO8ClqczisjnW4OJRhEEpwePEuAqT3bni42Hd1+Gz3/sY
68286qs7/uYKb89UeV9ZnX7X01QxCLXjvJkyWmT7PB6Q5012pV93HseLSd9oIlkd
qZa7nptyZM2YflFdu12hsUoCSwzbnceUNN+eEnf/7vwmlKu4sXMBs6ha+osSYI+Z
a02wEx1aAIpKAwHr8HNBXaWaQgYCZEFUF/DSv483Rg12jCX81uDvXku8qKHSZSq5
JY74NoVjIKIu6XKMBmhUwBMErugs29CbcPj4mdnKu0VeEOdBxr86Uj0+/C8zSAZy
TtN9paO8DfM7/gJ+LOpwd9ZH4jQYagaVa2XVDpWj3UCOllSW8cZSsdhf6IizM7TF
WWeZKSJyRs5+FwwCE1OYGWLUxOBsVjUpGu5FRDBksen3JZ17cf8dszc5vFKLp+bO
mDgmeEGWuJgMxl3S6iTWGB8dMtaX/7UdF3rJW6IMe5JnB/txyog+a8lNK9aiGVvK
xnoyjCQBprd4jAPhQO12sOZZGxDgYilFe+ornZZLy6INzz9FP1hH5e492VXBdkZn
9WJPmDZd3G7kSZSJY+iLg7JyWuUqL6/3N3aYud5uCTpuculQFSiiJVWg8ZVJkJoc
+KogRsh06nWBaTY6Taq2UO0FAA9sED1C2de4s/F0/cpOp9iFFa8PlSU01gpbVx/J
4Jl8OAQ2iffqKpE2/kr9o6CmOO1FiOCxzrs81Uo9c1bubmSJbvOnLC+5oltbr30A
5e50zePS0YtcT3rDuXimGdthCj5XDHomsu3yh1VpxEOII+bXajZ24qVtqknJw5Dx
yMrSFWFYSbzzE9JMPH3IU9hoTmnsI++pHBP9VwbfFGcFiKMCWsi1EVC93z5KN6cP
zPAIfHzT+4QE34ypgrpLo/gYxsyPQSk3o6eH69MsqnNOLsBh08ZQtRA6XPCEn0qk
bxR2FEZwEp7TQogGbA9MNWQRSteBFUu5Uss4U5qZrCIv1vy4bsVZl7n5BzNrxXyT
0/Y+sTm6wmdXKD5y/fBhr0MVD/DhH3k48agPn9kAOM2+rgvyzmscvwiOpLdX5Vnd
ZsSqKu6XiCLugzVodng/YMuH+3kqAD41fOIykG3ASMPseze7TgBEEa8EutEwcKIe
tOEnsYW+4lEX+Gqv3eJJkBdmfHSEDH7KLYVEg+vk6zB0leCiwNJFfKP7uzEecbtV
o1NYfTlehfcT0ZMC9RrZW/JuICOeB0iRFsiXNaZ48DFjgLq4KnEnEFhUJTshnd80
+og7+8mozSu8QWP43UHQXXGtklrt5PdEBnka2rOXgJo5lr3slUVR5Nkkmuw+9mXi
IdXM/GGJ1H7j5rznVJ1hY+/6a+icKqdTKyUKfejrBpy5miY7NfRExD1scukDyhcC
jS8a8bNLog8w9utpPOj/i18cIzc43rfkLlW04qH2d+VaYnSstLxD9YFY4EWvuyHk
G7oXG5skKeugOwdCf1ywySjRRrUmHVR7gfITdIq3fB2KYtoIhOZjUCHnIwSgsoz/
fvQTaWMF59h1bZNCDme0BN5g5Kc8pgR25fXMUxtHJv9pcRJUCW37Cx/kfvJqDr7z
jokZ/Z5zUTiqeKhtQSWc3/kdKrhi+k9vXdHaq/M8HcZOVawgDhg3iI/+sMtCKfxE
NzitQ5G6/6o/FM537L+ZiKsZnGB6JYvBjLa+EpZaRuvteOW25DY1bCsErFu2GgiG
vP0yY1QpstGcCivlEWGwEq8yGd5aCV9UKf+bVvfALGRFYKCIY5WFf6ldTa+vY2EL
YDaIauQVn6AYx1yJ+wvJHVfsYw1/+TllRmeo985wfSoqYoXnl2+KZ30mwGO4Ih7c
jU7XCLeUK6DCJ6FfvNLjtkTpJBUBsLpAA5tESRaJXDeHWbepu7I9OXMwNZose2H3
W9ZGhhWaelwjeTnu9fEqEfxOqxyFP1utqMS3mPSf3BI3u+E20LeGxr+gcg2817og
CXb3jNv1E4cfq4PUaOyFAS8S0+tdMMISGHPjc8K1wspSFSJvn1whS31KcZZlUr2B
IeXrQ83KSb6aJ+73ZC5D1BiKm+NJqguqHLspR+Ku+PtOH5Y0Ng6NY8bpalB7RAbl
Rj2jNZ5ogNjDZWKPfZYsq21eJVPL1W2WtOQ8SU9AJCwn7flADmn69kYBcNtkDxzp
FNK46dlzdlxIqTOf59nrS9hdMYIzfxKefUDlr7uE1MdVC/EdirSRRTivIQ7ZiiMI
x/PJDvhLyFiUxQVIf8QVVbwEcOoGa0jifOu/nijDBwFN1rD8L14N475028v4CGKr
9X9aQGSIUonMhcAq97C23VTkK/24yqO977oNkhxgav2frDGcgJ01r8i76L7RzQ+R
Xfe6eqCZBYD0K/2ZSh6w0buifvCeeqDAa1HqhUWQErYJ61GLwD1s79jqATbIwn4h
Bg8gZdLBiKLNHAmOrkTFrJ+5hMX6hPF6NBRWfpgMqbGA8shyo/ejZA9YBowXZKr6
17v0IHL80M2xLgQwkvUXxdt2tGg6SWBYRUHFPEQw5E68O+NfkkM0BBvJtnAWBgws
cRSkwhTqKaw4GkUsvk954/ppVvF4jtvYIPefqHEScOGPwr45ZF5LkqDXrPWTI/IA
uk7Obrw1sHNO9xAyxtE2uk+DWol5khhk4ImfR8UGBaUF20vhmqlT9uOIuBaOeaIy
i4RzjN3CzF+SgOiCs9TPlH6bL9rVb4t8cg3T/tKGUwvCp4ZlnXLS5kJY08VsTVGn
DuAS1p8pQjJPQOBENk7arWuMwIORR4vpXQE4DMWlAkr6p77PO4dvd0irhr+SJqWY
RbPsM4ra2V3b7YJkr0BtXhQqPuwLPQUmgcPHe04aRDXsUJuMrd6ic9BxAbmFqrIp
e28guP8Couks/grddS+x2LfiCJnE5zpS0eCdwUDxWw/H/yIFDkUxUaQb94X1yMQl
FMNeZF9VItcjs5KwQp45N+k4i1XaXM+JKoQQmqxOp5uE3LQAn8ETAiDz/gTwmmdq
hkJ1hAqpvq8oKOIQFFdbL9Db8L/fGU0GSgNaefqVLVERjydeTXmTA1LrVmiBdGFn
0fPiR+ifpP6l1Cr81nA8UyaW0n8qXC2i3N/t55VeE6YLAQmyHm08dqGIgWz4Dhuh
NSkn5uCJkbaSU9xtwqJE1gnAPLYDsJ1/Sn/pvlXsRoZHuYngTAybSDFbPuq1SX+H
Ga6uRGeaBSz8IrQ122rew5x4jIweb/YRryX0ADU4vsFFlL6YRoxKH34l2O9/8h92
Wf7D7XCj08VWEbw2miBjqqo01VVJV8LhfiEbivSvYX2Ml/J4LchlmwA1ZVLnDRwZ
pmu3rlgPGJIjFqRuD9nLCRazp/UgU8Aj838+kovtakcaJ35s56VH4ektoiYjIDno
T0lx996r0eB+nRVvxZU6YF5wLInXGwJsawHgka0zmBLjG5ue2IFjI0FFdWPRg0od
hVeND2QGlaHALwHlq0pjASOnxrmZeg5t3kmUKajcG3yyXLMDSLcTKVW4tGsE60GG
9zv3TMNEbNE1c0CewzhpUG+dvKoZgHdupoCAR7B6mHuu+vyTaeTT1sM7nAq09V6B
zMOPiu8C1tLpZyP2DgrIzIPnkNnebtrScC067iVazitcDSQSx4lkxS4g6NqMhpRH
ierPfS5J0qlMQbU5zb5vUSTCLIZLEfTZJf7sbS4tc7vXg6trIuvsaK14DU8q6e3I
ICzWxRndwemaAhglWjkYsMZTWCccv+RCeV5WUAFN0vfiMWLERr1S+j9J8gJLn6+4
fm5mpAiTc6vzLEi61gUFlF5zxW5NkhcQqiHO/g0WrKUDEf6QxUA9Sb0J7/jl3KYo
ppsIRnjfs4eTyC562pkCuR32KIbLZ71kjxcLa25LRyLSXFjXCiS5eJkvPKLiILEY
vqy6LzLZS+xXXz6r6wCgW1/xcxfe9X7u1idIn937/DqYdG0gutSsTyB+KwjeXQtt
pcgAsxT7s54DFRY4cm3kIWOQrsZFNjjMOPaTcu+SwY0UQbmRmkNkfL+4EP4Kza0K
RCtJXD6zrU3SLAzv9svt527y+BJT+7EBMFLlmeLYj971vdG+Oka1HlKaUewxnzo5
WrsAVwAiGGoHKVuFeSg5h4UjhmpAlerSEBtlQ16T5pWT1lRZQ8/MxuY88rg8IShw
vlf4ReL44oxiNCp7RoZthm/q5AZWYo0pQ/hBhU2Ih4wM2nBkpJGIylIxAX9wcA80
10u/iSe0K9ZR+fXrVkC/0tTnrGzQF7jCxe1Hubjpftv1whJa0lmlr7cqOgGA4KMx
NH6XbG1Im+whOgIxUCa4PfWhbhHpXsxZzlzmVogdxaxByIUv9bXoTPw7lWNB+Mta
kiY0KkTo8ol9CixHv7rjMq+vbvwD3RsLBqVy4pf3AKeEPhVPyPjS7FWtMj1OPSOX
P3ciVEVPELHKdSVYwWDE9LmGUXG041iZ+Iz9vdZd3pSUETya5vaMdvkkrfuc6KZD
/QbCjjX/X6eP/qRpWsXPuRwiA1jguaZwMqq0rBKdA+8GU3Q27StV20w+VIh8i85n
w6OP2oSgh3cmTL9yvM4b511VjCk//ESG/qfrilDSmygWBzHVmqish2KaZv4igEtC
BfYxJ6jAXQaECvklfoGt9l5LqZvFALgbPrKvjwmtoYPZaYbh84kF/YGyrvM9DSZy
sTxkcbf2LOzgELZNO7yPeNHsaaq2id1sh5HhQh4cIJ5qo563+4V8cZkZVQIeyVfJ
oz3q+49btvCL+36OUP7fWLIKZk7kpUsBJw+0ESnXHEClTI4tOl7jxB9QMAjKVKZF
P+svieCCcCEJ5WYbBrBy2N8/OYzPlHvINCdH9wFCbgtfQXYo+2Ix5WX0HFXas4hg
NRjzkiH48V4hIuxYQA4niX2fyuqXcQFf/sJljPowUJUFjNvCRTcTCzIs/7IxL6iS
zzp+Y+H6yU1fTh1k0WCb+YtT/urhKF766mwiN+1oXJFJKc/DHjdeTaG2NdNkLDF1
+gJyf1IlUQnVvXjQ9o4CYDad6tvU+c+xxu7DIBrFRT3CG5aRdg71QgylZAmMvAr7
iKe3vKXJfj/hwT6LVMfcSgZ2o5RFYZoxJ1og7kGS9/4kGRth31n9DLtAia3tFAmc
bHlfSQawyUftrMFbZzAX4+CFz64er8E41uoiCU7mxInVRrKmFrL3VyKpKVX3QAJ3
0YebYV8lFg740G5yTNpcH+jXnqOo4ayVfm6F4LBw5hAAtKHnLq4cBPxbMtC8hZex
RmuW8ZaVgVDLcIeIuB9ZGLtOoQyYnXy5Y9rIUNqky9gbf3sq+H0UdGwGfBYlKEmZ
gpRDNElvaxc7gQ71/4Z55/dxAIz5LYUzivQjWKtXkSNhc7vTZ3HFiCVHITBwm0S9
q1qcLWmhRdu4VWQC8PNGNCEk7pC4n/6R2aJeyyNGLsUcU9HzTaTqpV5EBWVZCbJQ
yRxnTJdL3w7hV5G6GFByZ8xatPbinY3oV5D+b+B5qIdRsohhVAFBssBrdEeCelvx
vcv+1DpezHWUH1KQMNPO9RjafEfjVGKtHo3tI/N6YdkK1R00RSx8WIUv+kBvgo+E
kUvWZykLnRcZjBI9ADVZFzhJvu6R/LmMWKXhTAnsX5kRz7/PgHpeloeT1YRSAgtf
r33PBLkO4j+v2CjGazl6+NxNbOk2QfDCtOrN2Fz4Yai/Sd9jtNFMW/avITX1N4ht
XIm7NeuOZNOvw+foaGrT9Yi6A135m21V+Ou0RIAd0zmYHOkhHA7O+rDObbkIKOix
5ywLnNdW2lQaDOGQ+oGEexYajZFDyern1u+7mnDt4Zx8/+SY8kUg19DwDuDX+sLS
HzT69ZY7TmgR4KksEpwksrexK/J/aanGSsNSEKYtbHHCtVjKr3CQ+N44U/JEpPva
Q8fiKjY2iwTWHQE1DJF1xWRbe/AC1dFVkQuHrm1MWao7y3VSHkzmvSeSI6FizXZQ
fKAXGHnYGGpKFe1AZX4tacny+oEFB1pByT7FSEq5eltiGa/RcK+Nxvfpr0Vs5t0H
Hfx2ZZLrTFysF04T5aENJva4geNutnNmcif3pekqfeBMArHiV+KOG+DImyT8bzxn
oWNwmy4hw5Rb10H0GEKL0TXDOVNsemPfASPTC6pyT5bcQS0xet+I73Q9xd+TNO28
KgmQEn02oDdG3RMHdR6IvKThFJsKTeAy1TGg+iy1NChzWdFGUjPLQi/ZvHDriS+X
zCNw4qOM/D35d1TQNOpvye7RsZcaVibPifaBfJMyUDhLMEWyQzrRYJUKXHVkGIym
uG/kXj75fiGpDnlAWS1LJEkCNDe3Iw4Q88zmQmuGwyj00gADBuq5h+Bb+1R/9mul
a09OL0oeEEKN2sRsr23LVYEFbBd9Vy+JcJvJtD9fF3HMm3ApIA3uL+2KuqyitYhr
+C/Gc5HQUJniidQWXGnGKfjFBNf6h0qEw/+NdtCWf3+93RXKEJN3FH55WS3rhV7R
0UTjzimOLInj7BTNOcK6H+ZOs1rdD+7yQ4MHsXp7Xi/geukbrvjPbtOyMs0uagbk
1z7lF9UeE/vYMnMkDi69p3fu9QIV4sUn0gX2XDVStDS+RYVG5LYAsotLbLzyrC4T
B2/nazHZyXNweTp42zog2GSQ3AziH5Q0IX8JH0BBVkliRbBEcDkkH4vvTLRnxWc9
8IEvhg7pY88gdFXHYYMFRto9UizqtQfvS+/l9uiyIAdnGr8QYNR9E3VIxjC2uVgb
eQ2q/x5ufwW6oik9bnoWT1NMnLeXvgkrsXQpunHbcVpdKODDbmPxEltOfR9jQA3s
BfcMznk7a5JZIkzg8zY9vaIduCLzK2FS+XYGS3V//xz2fufQti/mGUVErO5mYA3x
XjRgPHi1wxgVyGAS/Z2rlC7PZkqUWqfKWbXk2eMQHxlkmNDN4fXxWRExTMjz+u4w
CzshXpZN1Xs5NjS1AoXJnORJjaduZExUwSu7kfeteJ3YtvNhnpJJvBHmD7an9rg6
7oKgzSPrpJ6p5hnPhFdduZkpLf907c8XByTKdRL0ELAFb/sxPrX2zZv7ZanzNR6A
jidrKnKn2Gh09jwMvKe7qmOwJIVyY2zekVtV4IcPjC/+hqiT50AXfxFFj6a2OHMT
8Xb2vN3qwPyGilzHTC1OxeZSvoAw54utgBHv4FH/BTtVqLl613e/SS257ZpKjEZt
Bjhr1nXMsvYfrxiwSO+SiY+AzYzYcmc8W/N4A91Nakl7s9ZmNdvfnmZoHp9xRJ4o
RXWUh1/eaCLLtqvQZz/vjLArlOGgGsv+QnhGLuHQVuSNE7jYS0tru2SxcqHcJli9
Ml34Rwu1XQFGrvmTQpEDncQeKvLdlJ3OPNIWqBulhqYiY64fUA3ZrSMQINydKC7K
sxkv4SkHH/ZxPZFKd9xfW8cjF3Zq+1/5P3VnSlLzv4cymAp0aoLqxrV4gctlccbl
DFmPjIroPy99FkVl+SwpTDOq3pFLUTntzmxr/ybxoMF74Z5XM5HNjYK4jFwHrptH
18Oq4lv9HZDnluAkinFS5YAF4Y12yGVUQJC9pTfyb07dbAKtS7JcFdQbjX2W5qpV
jx+H/Gy7TaiBUSqyJ0/KG6HGU1N0l0zOl3gQlEsASO8NY4LTvwt8rj6nRUAi0dqh
g7gKnz1wu+di68oKgwuSJnYtBqsXYfj73ppfYN3WSOvDM7Q2Ekp+BDVnC0hDWQ8T
kM4f0qQD3skCDAlA0uuLt+QeaB/3jlPFfRfqJkUOSRMSq3xM10+kQ0+VFFISgCqq
gmHEpzBJu2068W00IZjy5JtV7UeHW6CIjLMMQwaju8Qdlt3G20jDi1F3WV/dCk2x
6bsMa2CRZwNh6fILPDSkh9ev/Vv/X96TF3fAH6ElF7En3UkXuQUz3+VfOwv9QvPd
3vguTATkzoNux1E47iZN03pGkv5FAMC+KDWF96rEsVVcYY7K3ge8uJosuwUaW02i
PFEPWuVTR0HWUFjkVMShnNbMpz+mVjZ5LYZXi6Gtr1pjT4Rff2Egr81ANdnp/06s
3ErNgh5Y4A0iV0/qxzQZ0OMPerXSekAx+OPzdaeoVajqeguePWdMYhn8prU0hpa+
4XgHlaEZGWQzIoXobAR8rXTNYAL5nUimE/iN/YVkPKBg6ge78Kl8t7G10+Yfehdb
oMjpUBObFY5ScOKcbOqc5nDzFswow1fNqq5d9TKU59HpgtsROK0GJIC6e9Ar//EE
ApItXz5j4/mIx8yz6eoQS0PRM+HteEISpBSrcTJkKfGRqUFbWzndOV2HB75yudTi
/FZbpGY+qUwGO2kBzYxELFWOI0RAg4s0dTcznfgWSXkGL49ij+BWkJPjP3koYLIv
eAUQXbfpu5k2t33MF1DA1hZPyx6+u8npE0zzmgNuxIN1wQW6zK3dLjR8jS8ivhbn
l2YRKa3xyCFG6B+b7WVzp3vqrzOjb6UkRRhHECoQ6AZ++GqooKEsKFTtpO1O7+58
XynXvMQNO9B4QoEiAVB6iBvFD28NtzDoykheHe1j11TGBEQGfGwTjSAfFwnUSdn8
OW4RhEGujUEysbFdgY18v1erX9UHg5Cb7xM518tbWXqK/pO63CuNkUiip6diHjb5
25wMmNaNm7t6T4whwE0QfPVSdGp350UGVSpgX7ozNZanmPCM9FlmppcoNj8X0Ayd
6QH9bVtmVbUECKysxEHt0EojErPOLXHp0b15oXieUizEe3jW49qK14IQ0ZtA0rN1
jahI3RR+YLumQamTPzkqxO1nAJbFfkuQxqBNkILyx4prRDz6/1kFMmEatHsNTsN7
GMPo1BSGBtj//zTgzmzq6945bAMRt0RuMZIppBz1L3M4hltY1nENvbz9+oH6l8D+
xky5siHdFw1oauEPb8MI3a8BbSJtRURULcPWJzKF6DoO14toKghLrn188tjHX2Q9
3GYq9dNbM9qmY2ARedHI97olgoxJdO456CvDJ+WVRdazPZN44vJb/V/E4q7dBQiq
4Hm8KDolDjoQj6MLgodv7EZ/L6/rMso4oDzXLuLYsLK146wFAXY7WJa+jH0uB8hB
15zePyR1GjKuTd1cPUbgFvJak383ZGW6//Hbci0uyTMoCMXepYXnupeYP9A0O8jO
P5zqXXeZeM6nQ80YX8hsoLCYEz8LyMGpuz3b2ejHc+9ZZtEXPwqVgbQJU9cR4QY8
Fl/ej4NtGedq8LwYrr7e0RoG9B+62c6P9jUnprueDgx8uAPQk1CaSKOljGoMTs+n
1167Bg3g4+TA2MVuMlH5Rv7iz2x35cHcZB3aihhZjJUFL1Qcdy/t1vGf7DTbJkKG
uPVw2OEFi8r+iZNGwWfwKgeWUYc4ZhMiaz5j3pmsMezichDmVlMaGd+TTFOGeMM7
/JhBsLAyXBXYsT7/7pLLXbx4H4gF9ZUhesEwIREzNuwpiA1XdvZ32HU3NdY3sxx7
LEAQXWsyLMuOBLWhq8M7huYzV8LQh6Judfn8iL+ZrqhzdWjPAWnZbnoR/LMqQjp6
vrk0qAW2gx4k3RcE+mwbKE66e2rmC+6b+8qDkOrvSQ345j4QiZY2bjToyYB1hQVf
9QNu2s6nAM6LhAc76e4n6J9eKkJt4kwUzT6SsMSA6JqcHwPadCq19vrfouGV5sSf
BleizXLsRcpN/NJ2dDbsC/wUe8Uu5kdH+fTNEUlXrDJi2FhfKUjm4J6RricWs4uM
5UCIAurnkPt4Uz0ZMiyQ7W4K5XZA7BBNF+ymY8a26njGhYc076FYu1b/L4JJ4UIR
SqWA/yvfxrbrdRsjnWWNafKxlwJUC/n7SHYk4fp3DChLG60YYuS13IbC1NcvEoym
iJ6R1gueexfvANP3Tu+BafxCLppesX+p7lPqVEYdC+dD+w+XoMmO1eGnQAiR2cOj
DT7UknhuexUzZisNsce3AqanTmtdr7PSK1E3XO0g10HJdk1lI9N0CZ5MXi2FqXlI
9cA52Rm9TVvswzSVFsP9lPZc7g1UX7mLiwjYKDxUt+fjVDek8I9iEgQvjBZi9SKd
jMIzz8bzegiluyw2O9cPIGuP9ua+BjM8rVRN+gscw6C36DO0sauZNZc5d4a5yRVI
tQicjMR0dAQC0dPe1cyNnKPBFJV1MAl8FMOJ7sr9BILMNvgD0PQFunrxNFQVZ5kx
IVdYS2GaJqUNFv/ZAJJdqShpO/XwGkumK876VJQ4OtZDKS4Bl5UDt5dwwrKXr3zn
QbaJUKN2mUdtF1X6Mg6fjE8XITw8LkfGesKDOtp3VoPqVSibUgPSVbbwBTrqJ2Er
KQRWO9GUTcyqBgQxgMGjLZSIvOUBKO0WxLHv0R5tq2Ng+oCbBwv8wpC9J4BA1fym
VD/suEcAdvq1tzDCOJ9ofT24dymBvnq7qa6ahO0hrDT2S5znB98i8NdHx3vwfjY5
Z4F1exg0u5AotBaOZpszru6Jxdy6FgbKNB/oufVUMWc3yQY0pK82+Nc5xKvaUJH6
jx2TcXJMnvfZYIxlpCtDhd0FMPBjitcgs79u6BLKbBSoC9lNUWVn6NuF2S+jEjqc
Gn8T2VOOmbHoedur9+m/QPQiA8JqQ8t5BUOCYNAXvbRrhn9UYTF0Kw1kuz/0AqC4
7i8pLwxawiVC+dhflYO1UfbD9fRzomprU/MXJVW6Gr9dd5vPMa8+Ve5zARnhnENR
FA1T265l6sKjKpo/xGAgD3ksNRHNuBTLIMJ0ExJ39Gj2/oZ1vqwHZ4emBE6pHC8x
/TJWH2rJH3HKOt6cdYGchtUOusFv2Pd3IrQrd0WHrl1XODwJ9lKsrT/UYC18Rt1n
Ro1XDcH2QmTEgVldGwzVNfrYE0OyKjLl01cqGhXFx8tZzyr8jJCSsMX2tCoVTD1S
wCrDXT1qyqyVRctVT1s9Q3XtUXfkQA9TrTCCFCXsCtBMbaIA+htGFZaFTOjisoCq
S7gY5QVRJprpJ8jdMCxB5lcA4tVYAHgkTvw+dD/017inQ1UjxS/LgbsIfooGwyTz
ZNSgihVXJmBWbY+IdFNFH5ftEo8DD5XF9NTQTIy/C6EAC0C7PE0GNDDrBbkp+hHf
0AuUBRkB85fKubiR/bD5VjtAx6FNTKD1BMj61yaccOibJN+8LPWDAmb/hZTR7tHM
hDJRSGvVpztnHCJ1Q7BN3aKiN8AkXGW+2tA6bfh1ojRleSOPkdrc95nBPY8Ht3bd
RV8pctrYK724nXc2LbewMDt4+TKLM7TtUcRQo6/5ykTLZyud3zRE4fjRKUmDKvtu
Fnj3M0uuXQ7A4BnaESVJUxJFGgUOW6NjMYLuSlUv/FkpOXAQdC6qN+df3snnHdiQ
cA2OrahUnpaNC5IGi+PVQIr0oZ+bfFzcd7dzNFg7v1UYub1734js9O2daB8090xY
vhr11yTIc4/XxA1Y7Mzd8qdtImcDDAgpn64XXU044JJ1hQX6JmKXZap5vis/E9W3
oaWuYuqagzWkUCn5/yARTHn35utuej09xjX3VH9DhLjmvb3y60MJgSd2d4dePmU1
1yCXrttUOF6/SRmO08RCBCGXeuqa+q7H+JeFeXLdUvRCq54UyYnCPPHtC2n3C5BF
/Lm6iGJNNdMJW+x9Rw8TwATsUvqPNX0E8c1Xo2mZg+vF9WmdzlU4z+kLmHghXlD4
QIAykab+YZOpb/Tpl7Z+bv4sy5pD4/8vSz1OCLgVVHTMmVkEiCfYMM6VwOJFQU9v
zZ4+f2ydCGosMzpGaMnUJa++E7j/8EIdEB9f6GRSBYBTJC1V/K+LC6hOXPgN340k
VltKHSdMej2g5JsNbui33Yf9uXH0uFfUnlQ6xJeUb62wjPhok1jRfgbasUDnC0I4
HKMDlm5U+CL4MJxX9VlCJqR2bYokn7F+ylwXPbroDUvzw1vABcPmyD1sSLtAinHv
LyLhs2Yj3RvSv69Q7QkCFTadDylMniurrjzsr/B3f1haYR7irKJJr/C17hU+VI6V
+Rj18oWzfrU3yZmlXQe/Q0feZn8HX4Ce11a5G2nzAlYe4zM3L/M5Dhb/ZoKxmX8a
wITPDxctBJezK8GXlByPvWvC8tLamwfpuyLpuf1kXk+hwnVWcXjm65OfTZnGf+Cz
G1DIRXpUxyCcLnD6eTtqjZJxkUYcCwhSbQ5nlEzNy1PqQpKOPfrX/zQzZSkRcncL
0hpVtVq0pG7x1C/OjU/VaPNdIxeelialYQ7gg4aV7YybM9jGIqaysS2SeRzmlUt1
nLVNEzeN6p8meuTeAWjK8cutGfN06OyYBjeEPWS7NksHtTSrNtP4KkozFFfRT3rP
ml/JFUsPNTnAEuvF/P2EqzN4PTaXnYgNgTBkZd5SH/zn0YWUMCTTHZOx/Iem3eZK
3ArsYPA+0hi6X+WleMve7ADT/XXfQtT2ZLekkaLamghuFqEFKzWNLrbHBvC+Kopw
N3mkmIcuSUooH3yMTCKpEuuyIarzlKp905pO1GIsOebaBweDVERvWWJePoVVxATS
qQxQG0PBhfpbO50lHNQ51LZCsEHziEZ7pcvYU0Yu1BT7aE6HUW1GWVKR54bCORjb
zXUKq+SDGkCwDYuCHmJ9TZtzalU94bdbac1CW+zYU/v4ARjhSEXQkv5AF0qCqURP
ILLHUzcqp0R+YQTFkGD4eepvlKuRlxI25kSbFuT9BakkTiVMUbjVLSXGL4xrQkD9
gyenp+3dIjDux420RxUgIQ9Mq7BE4nukrovHnUuL6yMkXL2m02JmwTLGSvrg+XQE
m+Ntbrop9FjhvDFGEQJ7tA7v6P0sUp8eJ5iscHx3hAttMOJCm3YeJKOjvwDgE2il
YQAnz4MaSZd/mCV/R7M0y2bz+RMR8uQN80Z7h0QfnLO4V/gmQN6ic4AI+OeesK5o
T/a7cREIpiIMyubIBPgJfJCsmKzobjqatZ31tSk2hytZ5jM1jGPi9Yj5IR9JfRG8
pbwc7pb2FUPi8jSHaNFKXmJF55qCbTh3+kpkucGe8YDPiH5nbQ+umFhGLXf+QxHn
9dt9U5BS3Uq8y7f/YFQh4tNAwXw/5VHGVvzc2b1ridkQbkjW1y53FQ/A6owbNFeL
+LHzkX/kXajKD14gxEzC0R2rVYOKfVPphLI55O6s6Z8mQYJoMHhkJjWN/mTFVhHQ
8fY7xehSMCunF9jHZ831glLbrmKus0vJ/w9VyUvvyHafwyoGE01S4aPMtRFJfjp/
3VXZdPCnORYNmqWpfPqSLIdtcCJg7ni8zF4Elw/Ppe9EwLqCDJHB+cMK01vLcbSW
V+fDvkzwn8GQ+yWikZU5jIE1wWqeMsp3UsIr4iTPiOy7kiI4Q5sq/U06hqyyGbFz
MXgE/awNJYJSOKum2i/PsRJRwjs3fyk7xtpFkibqzcRiyoE0chI6KrSfOJ6F1Ng4
s8eD9lFPhAMZ5M7AwhPf/azPKSpqFOtwKHmLWHDLLeYWfk4z2bIXmM0/48gzeZFi
XK91JPB6V6A77KuiMZePtsmu4cxH2PEpIEW4bakBhF1zGk5hDn+Yu43xJ0+i44os
AcZTl8Fc3MBYIsQVFK/eBf6d+/weWyRjrsgLY7onmm5SctJyk82uwcwJLfZMktye
JMckk5F/ZY5i1vLw4LbjS6q3HjoaAd2fBhtQ6Bc6ByA4GnBgMMpKeZbDyEmn14YX
XQ4Jq2JqfI+A5Oh642YRPD95zQ54v//hBHdyJNSTGgOfXfGXFoBvux7pLTU4LRKL
mYC9iWpFfy7+lGOUiVAVTNgAFe9K9X1JRS5KlFoxBqYsv6xukuqzJ6dCe2kDQdLt
bBm0+y9p15mh15Lm899fMdG00t6ZNsAsAqYG+7Z5FGYJxyyyUzlLQuktxTpEDj4V
ejCD+2G3yVIsQHIiaz5j9RVzDuqOp6kBGCrKrejugEjRL2ybSFUinKLjuUnD9jL/
pAC6P9WeFvj+igKJZc5r3Cwth1qZ4FIRJReuHuPali/nWkY47f1Y3Vy7Xzoi+n/2
DvhsBUvDFlezEfnXbNxjjQzLFueKttacZuOXwUu+OKmb4DX2edhqpbxf4vNIkmmC
BdTDVATDysXhHbM2F+DTx9SEeXr1t3h0wngAUY8oa5U0f4sgEqfjgy6lCa0e4ygR
cWWAfpBx1SmXHmUgUV8nf6zsIKy7WZZcjHiA47R1mkx/TZ2yXNJcik/aAZLC1cRL
Rr39xesUuc+w74XehLcYSp+9+Ct7kMgBEZG0dwl39MyviavC0uxzMTfyUUoYIXW7
/neUg1SEqjKLW0Z1kDacRq0FUH9UuLeGvcTPlXlXs2ChlIJzzes9ZPT48ORFpJXa
mFs/Zo4AhBUQ9sZUX0zZ21Kcuf658wH9O15WdwJ6FGpJEpIAW3Cc59V/+VfXnamh
prTO53V5nwUCFT3mRajHw8yK5Gk0MRbmSWwlFPxxFb69EXz/xKupr8KtWYm3DtZ4
WxuqZMRijAEtfyfKeATTlmYeiOwA40RE4g5YdGIhhnXdN9oOMXX2SaXH6SC0e56i
vFzr5+mpNaskP6oZSAsj6JdAKpRCfom7380UjyFCX5SVQx19S3yU2Rc2xuxjRf8c
PNopAiGYRY/q384B3aFZCi48UTXvDHhVEraqbdA8/34XF9DMjA9BSaNJ0uAHCcYr
ahhF9AFNmVy42o5IEXyaNgHN593L/wzxv2xKRKALXl4tOP2WQ0wOww2ZJ8KJC3PG
jFRcKHHJdUNwLrkK4/q3F0uokg0jdx+LTpcB6lEtoy8cSlFsfbjMDGwonoZMqNli
FH84T6xsi+5U9wgRXjvNHsThf7orsG/u9aPs1zB1awXO9yxFW8bOpsfBUSjCxWil
sytGwBInw0gv+DS7b7FIDvGBxhySMXUBcFMOK8NPq2pan77qgPMsHCWI2zcS+vue
o2MkM9mPqH70tShSAdsFTuRUWrMLP6+0HxaB+IrN4DuhVcwyynGw167rBg0ap1AM
l34NzhdTqs7pSP76NtV3VyuskTfm76EwSDFqXuMSb0cDiejnFv8Lr5xehHFuSsTH
fwnOouRit+QUTbiw1kQB/wu67lCT80ybCH7BWqSlEPwK+ehaEshI4r87iPEiJOeA
SJrFxmUh32MBL8sNJle+dEjBlbZ2r7TcncSh+Mqm98x5+AXnytys9OyGB/vOh5wN
s8QXJcb1p6iq2p5usN1Kk+3DTzwxLbn/B2hoxMaLRzIkr+WoufhtVx3FF4zW8nrz
BKJja+SyNvU1BamkREto7Ep5CPQclBdfNtf0kyzsr9VyYX/11ugETVEPhssHBLsU
d9BquCF6pvOfNjizgdZw1N46Vht74sw5xpNzD6gjPcVdYnIpb9CFu6odBAPmcmM8
Cj8GIMNVVyvWc11T6ahMxg+K7chnej6lXxwYZiGZTwz3J1289EoCsp6k5UMf7jvP
Ha/e2e5Od98BBDfN8xPCu9BGs9GjwgxnUxyBuNwRiVgvFB4NP6BD/huub+q6ysQb
gzlnsv2/EDDiTWvf5PW82iStTcgvUQXxd4p9zNlchJqCrKDGqqyxp8nslS3i10Nk
tiqQVFJAe6lUmfnxByXnZBHPf48zut135ucVWfRZZh8xkwKcb1dO2dYb51SJFDZ0
GB2tdIfTc0fkPB0BjqNLIXJIg6vpxqnhZCctaglVu7KUQSHrtP3asDTPoJratUuC
BbxeM6ajAD/EbwusJ6G5ZZxWvY58xMe2+mF7Uur0wg7koTp+qFczylR5XTJ9HH8G
klmcNdABsYp28VhZyiH67XqF1RkNYQstIgtQRh2MPue8bGONT2qzgbXXSL0TwZUp
wxxNP+/W0iB4XTI+odPels/MInBBv0zTKYYhK6/gQDnmGvDNtNSwVerE8ls8akY9
u/0CJSIEmZ+euYFva6bWQaPU4s0RwsjASeEZUBbPcPR2iVo8uWbQuAIifM97dBnU
aEsYPJd0g/NKbve5RVQS8SrYRwZ7jPcxtyJ/xxnCfISHBTLKtt1nUhnvZ67Y816x
H/mYist+ys8VIkNLkreoFDCqcH6xWb+pXSPdF/z2R7YjpNzlZY9DpuS47JEZXfZO
mMuLJ7mi7IlbreOrws6ZuzImzJArygBQ0fjsi8xxwrd2s7cU6/FDNZn4sZnPPk4H
B0GGeJ2akJfHuZzzd84k0pbLCFRPlHn+qyVyha0qPrwdsfmw4gKxHDsIjkkgRRtv
ZpT4rMcEsLr6LsvpCESqTgEWXK8eIVMKJVukjd85YUNJit2Y/8m/xyL1+8GHsBO+
zrWcc636mJVWsIlPT+CB7PErcKnA+AVMdIFhQPHs6+6nf/KVi9cXe5FfsWwN1J4v
us+z8LEVF3rv+A2HzyXSGv5VuxbGH9bSpkBkFEqvhFajAVW8riFdqTSLLPP8kdqy
3TIi+gA35+YrSj7QBReD5QP+bqzukS2za1pLZO8K+pGcOo7Gtlma7dOq5Y9Oc/k6
E7x0gf9jrW40cP6L/uTMp9592ZVbHz1x4p7kA87hn7WgkG7LmraLVfXrthlgFjzo
/ZqtZ1dayf64E8wldoAisoy0uHbnhlmfK2TjLHFj08EbZLOIJhbiAR+ZZ9Hz+DnK
dT6ofk9K87Aqn6bb2LbeiIiJQkJnIuRpmbQfCoLX83BZR5N8f0NJlTDikT79u3jF
TGRhEjnpBt2ZxUSzRT/00G1q6TfB5+ucp+MWmW01T9DbKoAASNnAZvwCW/X1kh7B
5bbXXFuBPd+1x2WrI7XWQ0Z6k7rtXXEKfdDUVlC246U022x7tGaSRFdKu60dF4vQ
qXcEl5SiqHk5oSDBpGuC58zBgyCTfCy65xhXOl/COvojKo3xsBONWnIenV3c8+0F
PoiYzrgScGnC4TJFGWoZm/dtbQd2KWjTq/iOvsXDjEiGr7gviIcVyOoFyz6m5ScC
W7c39+xPw0Lw+AUIS89SsbHdASjSPL10lTsZhhaNQOoXi7ysKQUId4DJ2oMmZAzo
h1GA4DMBIjC153sjQFU7QHR0PCRNa+tvGAzAnqVqtwMS5RZGOuzwHyDIgdDSmKjf
/WuPdKLA11YBt17MiX/gGpvoApkdmiPP10YojHBWnPiCEnexUsXpfvRqptT4EBEi
DzsxJmsGN9vLodObmRGNe7l6piPxMggfmgGsOxbXD9rpMrPlieysSLuBivA6iGML
wv9RKJghS7Ed1jLOH7hHGATXkeBHrr9npNLzElZADXqsU07sktRUp+M+JTXprnzT
pa4S0+PrVQMYlo4miFH1lAfaH2qLVgn59j4eKjMLVYF2ug/4fHN/kRSJj04/nE1s
j94a5YOuSs3EpZ2q44pzl8m2Xz3QsFSFBIUg79XmbXM857UZ+lk2wnSgZ3mztCnq
EqyJ2Im5HcX5Cb/qYM3k4D1XBl1ewotOCJqJw6xBRzVDDXbgjQ8ebkxKI2ouJuQY
Ka8WOSdHLCwzdNEFwEr519WaOchUz2e3z3bAhduAgADhl0tcGA6I3J6S9pednMY6
hg7P6/Kp6AW2dZgshZC+ASanZSO72ozQOCaBikj1eAi9rJpCI/wbjPcz94h9+AVR
lNMZv+CPzEwtQciGkGktcNoygr/bAv8cbZyeS6grEUPvvNRP7GlJCxHem+9oOiTd
kHC4nofoP2LT3N7+Dlwev2/A4y+JuYliramxHJPtWoTWIfOKhsvP7eE1eObbyN/y
qm9gbuSKPcCRo7KxH28kI8RjdNzfK7aeQ4wGa8czYt5lAWoPbORMzCmYLXPilZrw
hZ7KgEsTWrVs2kr1RMiHNSeff5kDlagNx/w64rVhx9kQlZHIgTwgWGtIdRm1Gxb9
N0dkqjtz0QiY3agt27Y49XauUUB3adAQje48tPKmnXbc5Ty9yqTttIUAzpBsVYNu
WS4ZmRQvC6RgNHGuyDI3tK0ety9lvu19255/bOf5TmuG8porQnRO7UBAdzp3Nrvb
RyOmg+PRxCSxJhdeOlliDCw40sMVlzd+BgpC74F0hfluPP351QbYj7ufIi7vR+Zt
NNbGwHgOQ/6yMqC82Qx1d/RZJMHc5VDaRGsfPN5WozT3NkSdhuvPgLGCnJwxBmQt
5Ql4CrWju6+Gv9TN9zg9Xr/2CD6tF0IZobJXlRQ5UmAxLM11RdFaRqBgLT7noJ19
jxno6OdfarSmC6NboY486CqqYsEDx2tJgu6ZdwHHWHIDEoA8fEokxHttzzzdGacx
CNliYf84pqDlgXsL/8Ga24AxSQ4avINiJBQ3+BemFu/1gCqcdmLxv02a4VtsU+w6
VgKBfdMkJaiAynQq1ziXP3gU6QMNyEkwNwZrq9ol0l3WBYVog3JH+a9YNVo8HghG
Jfk7Gi2C/UX4XRsqGn+lBAqURoEC0rypKj4CHSh2gZahMvNqMXPsiRlk/0UZFCV0
w4mD5wbDUIt1/12UPhgJYLYBi12MH8cJUTyun3aJPFQ75wyGoKbZw1+f5AGzCB6A
C7Cddz2JHLTojvcLSbZhKkijr1qDLQv1pgrgMybAIqQiUYnqSKvuE/QnwdqGYWw7
fgrfuyJ8b0gNg3BdscxLnTRSZbGIiFzAqJtYEIPLOxW/ss716ddRfpmY5TMgYdff
emF4Oso6F+e5XGbsHFeBjs7kY+HKh+yK+ftR+pgMdlGsevMezihF+kmDZTIyKOoc
ZOXt/Jir2Ih5Zrc8gDjnHwQt2bBPYFtgjk50XZgloI7zK3oQrazKt5LugcGnOsTc
QzGi6k/pEUOU10W6u8GsgHNSAt03ZS0khhGVPPEJDpxWvOq0tW06u+4X7eKuBS2j
OchxWhbmfPcuMHGas/+YQc9j+dY+y2ezJncteva8ewuxh9PBBKDhKsVm+tmUpL4h
3v5KclFcnuBDPqJF9298V90ZVKI2g5c9qbS0sPGdjT0toaifqQVITynVTVj6d3j/
63K4zbS1cqVJhtN2CrRmUXJZJK2z21B4ml+C78mZncApd5cXVmJQORswHvBfNRSQ
AH7qCm41rJV8+EfWtZTU3Do2gHo7z4Oze9oOaMVEcIsSrp2NCm/PVY5k5Fb/MBIU
D1ZwwhqKzO7Zi3SAKICwuacphokupBw1lIEXc1OXQTBmc7uK+8GfGcToEiWQWiOm
RRXRqYaIjZP0Hf5q0jS+8sAEjW3uRDDAti6QEVEaLEs+muXg0Hj6Zjo/cKECdzLd
8CKeO7ep7ccdrjmzr13bZDEck3eFZbuPDpFc0mTEHqTg2QfRcW2ASHy/eHO26q28
X/wsvAmF+X2IEg4J7P8f5JLMWyWTOPupaCALYJAkuF4Ggv3SS45W1T6c18E+Mt7W
rYn3DVls6ZFjyPNyiqyToQvJJd2wPUKOUdW77fBoKF11zqpszWPNcFF9OLFF2UJg
SANhcLB1KsgI0Rxy9/Es6y3B6Qy1esIhTfKpqZEvgu8irF2LQUN4x84WYJn/HE1c
lzDW0JYh4YEiHiNUJXkQBsmnGD8LvTCB9yUP9P1s+c6eiBfNYf1lHeOpmRzDezSy
4WPOdcDsBwDFWFGa43L12gsaBT+bMrOKmhJ2kiX+VhvP9rwVyy8KAWz05Yh9xca+
wKQfC/qO0X2AJDrYUfXc/xi1AfQTYiuQFZBiGSd3OexT7FYzxiKte03LEaeiKQiX
TZqkBHzVxYt6K7NisvzfrAHbmGHglLTvteYnMotuowVW6aco39+EQENVkywFdo4n
/ccrUndHVGjglR4ZP+OPEZA5qkcewf+guC0DRSE1QGJFDZUckykU1W/2E+sCF07A
9pco52oWRKGZIDtyYPtj23aGGk6nbTUR/QROMGjZYcPIOSV9SJ6g1sC22GGFEV/y
R4+D8SJk+ph8Qvhk7qjK4QorkoICTWGrA/BPLYyVz7kZlrOb/T/wxQ+6EiyD19sK
PxdgoTrKSE19aKoeNnUCe7kJD27dKwbi3P6u6qLIiU902z4KEx3YdvG1GSMy8Kl6
mFKSMryQHmDIRz1kjL9S8jN1z2iFCEU9frc1XQV8FE6qwzO+HVV4WL4VplJGRycE
KpBSCYAnH3LPMsz41LU0JuYqvc8HnvJQG2GlrvPq7IG8BrSF+voh9anhkHX5wfqY
E1gpDqNZXrBYalg4b5+LhKAD0il3DawwlYIwGsUYP2y5zBm1hyyb4LA39K1GLc5D
PV8J2pp5DyHvEjCVPVrc+zuC1/zbwmkyPvpvfHX/9MRgBi1PizvnqG5y+MTr0w6V
iaXOj1o8h4yiw3+IWkf92N6eHgCIjAteUuqDPVb/d6AX5Zyc+8nW3+4FAuWxrRhY
0WJFVUh/FfUoAXXHYfYNA017TP91rXs4ac7p0BgZgFShetfZaSjD3AurXTOh4wNm
81cUHiz+6ISauavHSrMOtUFFcASSON0RVx+NMVnWex6SgygU5rBx5gOiTvEHD/JV
YFAyka7q0eEjDyLYgXxbKFDWGHIsOUCxYjlRwZVRAjFpToTjP0Yvks5wGmsPAmz/
JhFPKdcmDas5Z0FFm7upDtIaSBa9MNMOc0fE2Nyjy1cxsl9dD2iQLNTymcvH3vtY
paxhgRmRigE42P24Pq0tJTML+D8z6YA7i4/kFrR31dym+rSZCrQhF/X4jzyXmTAY
R5rX6GmqBhg3HHWOCFk07iDYWPDhWF4zVi84NUFrL1NnrsRJVJkyRV/jY642UFX5
NkeFTmGuqQj9jR1NMEIOJSiLzKw0aJgrkaaZBVtNKmLgbvuE8W3TkZJCunrRS+UI
95LFlnPNMQ3/pCTAuj4WVzRRwbh0E7M9Xm1mPq1NBqL2wbbduM6ZkpaRDSFvMy8L
QJYe3Iijj1jDXJSKPNPD8RdQM9k1vmKVY/A3/G7lgBJxW7G4AAGR/KM54x1T/etL
aPWkvFpdmp59D4wIS3xinJGd8MN9mqxyumETIWDyzmNFkKHi7PGnokf52ugs/qVV
8bTHbzqqn/x5UIv//vIogU5ZLVZqlmGrCOJifxVMKUndLzh+UlCG2qhNGNeIhb+G
a7qrCMduGKyNOic8APNYOQNEibqZ+Hx4WRJaze14M++vfT+46mnIXdx027cTgUIM
ZueuDbmjbm1PI5PFCg2Xd2F488eRSzndTxh1vpcYsSy9tx110OtNu36rifaECUBM
qBpfASQQjfIhLmRahJb6nwpq0etpzAm2tOoYXc2B+73JzN8FpVnyswgN69/98kPn
RLQG7Dc3kjtpnokBC1agLXN5QnAGoaQbw3QQ74kT58B3oOREmp1TBGRCHhizYZm2
OC469nH20qSQt/11WG0eu4xdQ5mK9PO4tRg4ULo6KBrooMxfPsZWJ9KqpNXxXjiE
4RPKLrlX4ZAV6u6XS+YlsSxHUQ2GX+MLk4+GyWNiKPX1Yw7HEc2e4CunS4XPZ0jw
tA5TXrfB757TrX/4w1iLSvSSqpm15SV65l92Lin6062PeSF7bPCzDxYkTQ2FB1Sc
nAHizpzRNb4ATVpWFRnD54fRiOZaVwWrcyPuqIfaE4bUrVpN9bso7hRVCpka7V5e
IH3j+WgbXxuW5TrGvMHxPshMQTfRAj0dFHDhrZywzRE6agaIAIyS/fOSqCBOXFnd
YDxbaMLmSrQOHy+nE3nCSrnFxyC2m9pT0s3hfNUF9zWs4wKnmSXrlAYqt8EIydE9
SKrLZxuoHpeorYj5ZH71E25KjbVladObmsGMeO77McQDzlRZk/VIpvOv43u865H+
6CwfTPE0K95c+vZmgphH7Too689DbgPjELb+S9msYzXWKcQkVmuwSoa+aJS4T60B
t3vrdevUF9/QfvGL4c0llnJU9TwEBx8Aqlu7pvWQPxaVppRxNAosUnANAjbDhcEX
oeI2x1hUH2gLDIOBwLxhtRlkkatLww2LRaDZlbMuNwAtH1fRxTUzJH3xVVj/VQSp
J/oKm5erWsnxs16ldyipbLvFwwYDbMhLEDcrH2gHUpiRvdyfXhC9RRZOoju1YsIE
q/s0Ith58d0MJ7rToaLIY62nhek1y7LwghEBnRbBBaTIVUDjC1vBsdJSpY9pXxnS
5mlLAJcCifOb5lvyrOEAsUXrMW3U2tiLKmA5O8N4lmzXds49CD547M64qN/10Y2J
g2fMtLXBb+RnvxOjIilUfbnLIYrBOrtgYraewxExMi6+AbwoOBylI28UTCFP8OvJ
YL6C3XU/YXyzrm8fUPUKxJl+V1/CYDfzw4yed+RpH2XhAU9zCeVCsSZl39mpoeDH
FXCUA7uhqm/u1TxNdk5fakc1fYtrw16bVi+84qMQxjr2J2pX2l+A0+xEea4qeEkj
VKnOThuDib1Z04xx4Z4ladSZp3hW5MLihlc57elSvdKxiLj3W8zyEKu9vfifxw5/
QsL8Wf9Tf53rRIygmrJWKPDxb3ndDOhrCD0Cx4dIIyv3NWo21UGlD07r0uy9QM/P
/x7V0Wv7F1PBHsKLq6mJFGYjrc6e/U4gQyUOW5Cb+KZaZRPtnYrHjIPjr8qAPFpw
zwzrpRypCxNkC+WKiCMevXf3bOzwC+32IaqzleTwLE3xmr/K07c/8KFgjeTIuevb
LiqlxyjN4WOHsB09BKuVml1StQQPSV1pF7DWanVqZadzs4xWKoIvZNokleOWalXu
l6e4mJmbqb7RNosj+sIKa2IiYTn0q7J+Vtyv1weCU679rzxTbpAqbLiDTCjg2zaz
ys6v7NnM9hemvBC8ZT7L8rRHnKXCYYGIeQJjwIgrMiflDgA1o3I+aPgKjxONGCoq
heZ9pEp8pTg0F43MGGgcDl12FYJvL2sHbxjqkulwtXJyU+k4GAlHfxn93DhtoX5M
MryfhD3lxlFfaHTfH5LX+MjspOJnH/Yonc4Dy7Yzv/ANqzygDm1I+cD9YT/+rcGw
kXrb3R4mV+eCiYwjmRnvJCy4zKOb+UoakVzsG4H6aLWZ7pn396HJcoZFNkWr1jFH
LmGowX1zARFf+qY8TYiqDM1S9NypJg9mwpjQx/SYNvDyUJRiL763veHIppvpUuSj
A4OflT+0crrX5Fqy5S4jr9hzhXZBQNXRMhEsJUVnywwqgaYMKh2FJoduUvecvjiB
3N/wXDvAWy/zDo8PFc/pDuib7VFiG6qaf5a3jPQLVmGkibcLS5wKQh4OD/30sZT6
8Dy3yyQDwDm3oqmWO2YxrgIYBtIzwjsSXaICERuJS3NITIhFS8rNNKU7J746z+SI
HzwQ/6A4qeVFZjIdevS36yz+nWTaeVWtV1xYxtchbEw2qzEzuAo2PG7IUfse3qAW
2XMW4NhBv+M0rbO0I+dBJAlvTSH6/DT4YIzW1r5wWxFibDNoa/ji/T8OWm36gBrQ
70zFy0YuZFaD8JgvepAtF1JGyKvrTvqyz3aw8Rb0xEYCaeuA5PJGCz/NOcsn/n0G
AGymg7dNU5R74AHo6WRY6fLRN2r4WoyofGwuvFF1Ly3DaG3RUxLHhzj4Al/S613P
3SfH33DGjU71JUQSyFqtA45rAQ7caMtc737yT5kBs8V34e0dBRXBOpQU3vMFLiYY
x+5V3Q4yqkT5OzQGeOGZRmJLZy+C4bF5kcpd3NDRYoqbD41pWl2PCNdXVZeovXw0
uDh3K/thhu6uOFWcQMeg5dkAOevCH1K2jIzFplivaSj0ZtHbUc48naw5VLzqN54F
dFZjfCn+9MguIZ30DKJi+bkt9FTR0FH7O416O42yaGgxwh/531qjY8dZwzYVQSVh
p6OL6IvP0xxDOEHBUQuYA3Y/zZY8YrNBv2rUsYfcqRu0/A/keFpqgrMBgYoDnqAx
AQPSGCEKSbSGtlPocq1gMAaKcBBrkQVb2Zd+tRmXTduvy1tm8mjKvcgayu+/Pk0f
uXViuJTX6tiNjM/c8KhXxC59x7o+2LIvrpdvUuoVATPrTJA5P9nGezf1kRUDmfye
8AwRUQ5icSscP45fj8x9Xcpt1X8N+6b95VwJxBm/NqkW/ud1p7fszTtexBtDZay5
jSakg6LaJn3kw7as7ffO/599ZF6qXjYCorXvB+Oxxg63eWwcsrUs8EpmwIkv1Iaa
HgqSQC76Xm369TwreVp+QPHY1miwNadFHQv9lIqVZwqxKUYisfGs4kl+82thlgyp
AXm9w5L5tgjyaRmMsnrRYL2N2UPQqgoxLwodUshUJT1OZje3a5DUEMEqpoVX+owh
3VvJEd8bE+mlqJQyHpE+kxgWL2cRbKO75kWgcwfGV1OdgX5ZCsYoc+rAMsSHCyPF
xF26GLHYDuf0jCOr6T4Pnq2gdzkWMhZQJPe7FhqbRXLM0y5HboJjTUiEJi2rFxgu
atHrgmOtGHhbHaqSaGsvCFA8tf8n8PvCzk2r3XewQ6RwU4bokGQurUL6dgHbhkkU
xlLsoL4x6QWHt4gn5S96PkC+7PLzifKesX/pam914oyN8zrtgqjPwziTCWXmio4f
Vw5T/KiLBijWcvYPDSCS2A6+43YjjE6Oi9UoPeYAPV8IxOG6VCpShLoyfz5fastT
Z7+993GibUEdrLhm8SBlv1zb87Ep7Fc+3gF0bFiZx13AMCM7PrU0PptMeVZUsU0J
Ein3G2faa8HeMHgUhb6uXI0SS1VEHqYUFK6GKrFhXI4ZHnLjU5kcfvZzu44Beck2
MlqfiMJ1F2ktUgXcTj2w6ujPTfJrZpSL+yeRvx90EmLr8uO6NTiDuQHhxYGQoaBy
upcXZ/BKKJgnRg5mqIk1nnxNgNzpAUyezf5XkDpyMlfXu11kbrPzvM/U7M2EPKDZ
2tDzK96twwlwH+Roex+JI/CqKfnhTAkhY5K1tjROjtgWWjyHEP+O1G/bgVBCttms
qs9bd3xemzBdLgIk9sBudEpQYplk9RbgXuPp7vQczDSMXEB2OJGuH0N936O19NJY
s3tUTZ4fmxovnENle0dM+scuSALcfcg7fhu9PFaXtvppvN/ev9ax2CUsJMuVYN4/
8pXyJSsBhLAkh+fdZtiq88ya4FXROh/EqcB7nOiZcxtijWrv2Hjw/d3TL0FiGpAu
4x+R48vJjVm7SO4Uy6vuIM/LAH4Amf9X8IldPWis/2/Jcb2ec3fvj9Wc1dehDeWE
2OBH670U6hm30l5L4ros6VvaZUofTVDnpnHr6AIbH2Wt8zRkx8vKJZb9Bmeobw1E
wquc7H9Y9Q9+7F0aOWQC/8f2SCqZl2bssz/GaaN/QVKzx7RtDNADD9eJJ4/ZHRmU
kHdrdprlXl2ivtaRr0iXRcu1lIzvzEShMHbEZtMop9NFe+KCz5C08iztV7Gg/1UI
fmD0By4bbJklMo3JmWX0jnn57Cgj8Rjq+umheQaxv+8jVf24r/BVdm6vuR4vNxMn
yI9gff3rj0Td9bjINibDltQXpT6CcGUGzYuTwplo16Xcr3kCAyBXoLoD382ZWj84
nrPyHVtwx76sV92FBLRKO3vcXIB0JHOSh0trNmoLaHZ2IxEAlcdwWQJ3kFQindFt
NNhAWYQVeS1PtAwEget0fHqRuStcStI3eUcji2HZuRtZ1fM7GjT5gjDmc6TOqfMq
Nal247wf1kHrhLYMzED98i+Wz9xMzWgQb3qEym2BnrFCNWiJO9wT1Zy47YnNAl22
A6NFwQn1Xkh36xmxK9Ck4LoouBu3/D+jVOVKNvSeP0tpJ/MZQCNuYx1VcjIEFG+4
Bd6tW++nHrhw+FqpOKpL0Zpb2xLp6QL5KtNUJhL9WM2+IRRWtmO8NfzuvJO+9sNA
5IpB6v9BnGUhIdgZsQzs0m4Hih0ipa7j5wddCTKPV+TwDtJ0oAUMyFE/Pxlt99iQ
hCTDSHFeYX5rtTQOKU4c/eYBfysBWZpi8ws/ELEGbzt+6bDDzST/O2rmUlY88O3s
cDJpW/l+WIXfehyaO8UqU05zgQXhev98Cz6bo3k3K9+Ftjj7h77MtJY+nu5f3Z0o
1Xidcah1rcakzMhR39GvvpIRy6+lfx8p+vOBfRgWmv7h2F37slgbvUuSdC1xProb
JayNJGU3Fu2ptkHinf5QNjTJFHyH1oVyboRSDe9cCmuHajnjkVU6449LJ+bBjBGs
mMcbNnyrl/aeX5u5le0hdcMqqA8XY4gad4xgb/i1V9TrMUZlfYRqNs8Hqddsbc8n
hYyH2OvZUUg0JuRSP0r+15lGty+lIrCbQB1nAos5p1rKMtifn2fP9rmK/TwLluOu
5LpAQTg4xNYY0K/0m1EhobRfJXvzk912FgdyZFF/iFs3Pf4MxDn/oSByC9V6X/pE
4g7SDLYQeTa9Vespn/RU/e9DD7/Rd5c4kyvM6kZOiRS5+dW95EGi7TmLiDJ3aTYn
aFPL6gb1GWiQ6d5RaWjs3T4xHukqT7qMOxPlU16X+CsW7ABYrMYD+breVVat24fA
JKz1dgx5otlJXkuGsUsQw6K//MLSbzLl68SI0EZ2dOXsihBRikwFFXAlfV7NVPjT
/i6N1MP5h/distYTCxG6dBJkyRrTBhxOJIX8pvcz89WaST349wEYysjdxj7o57Ia
BKipEa7EkBE3bzJtNsNPOta5sOIBTB5xfk0d9I/xeIQTdJ9/eniAAxUWNXzGXnu4
xD07t2GrIIEgEIG2dlZOpkP7ToyQjV4jXx4GBD+R5uesfIONGB3R3oYN84Puxvo/
K++VlbnpjeytxJJta0NpyDsZ7bSJV4+I8xIEGDX7ZqWecYmIzOdSDT4mBDHD3sxn
coXH1Y2UYuMqasBfaFbm6LJ7UiVfAQcE9GYpffgsD8EIb5FqJqXD6yrK86CN1x90
JIzzIGHViDcTYcAY7Ek/4/5Jh70W6wghX++pLGHH4WmHomaPq2yL6BHH0XGbAjS6
B9CSsbXRXgDcH9Wo2lKEeiT7f4xNku42FfJFFuyiUxAXwvEwDbgQI5gjJsW0OxL0
WwTP/9R049SmJZCDFlj1KMpJEq9mw8F4+mYIh5Lz/AKQfVX2ubNIjqN9CfhM+Bkb
49E/c0yrYNwgDptD2EDkr5VfXvMm6aQHjAh56asAfhn5Q+KKOtzJIREl4xfzuU0j
oX1dLQ5CQ5VwqcpSZ8OTVqf+Aq5TAh2QBVL0W41XutC0waH/y9L7qtvtyIxRVYQm
FmRsWxlUg44vcGHbNwKe6qIYopWZ2Fm+6KCj8hDtjJU7fFY+q7dkFXU+VFAGNwMz
qC9GgArylIoSfTgdwKEAuKloiM259IaQPogf7OQslZn4gdyeUROAJgueiWx8XjMl
kF1+Ndnui7yG7WpZNGI0ESMsrPzofWISg9hHnRUwteKKeSEp1zO4QZugtju38wCT
sOiW9Si6+n52KZrIaMtqwKZzthHr4tmES7aB6VUVkRbnxSQ68+SotjLsy07w4OGs
7VH+1/pTnfeHDjuGZtFv9CHHWtNutcDotQwelG6aYJyHmNEcG7rF02kv3/hLonTR
cQ6HIj1GJ86VHR3DlU2Z+OTnjOnZzNHSx7wLJLJH9xg71Pwq5NRc9tDXjbDrjbcE
2i57ZYCxLszqROR9BKnp4AFcetiF/WEqF/xStPfCu6QytVszZIU9BEZJXu4dODU8
/SaURLCsGeUhZ1JzgFZAU/j2JzXKSuqA1Ls8vLH42EawVG4kTYx2mHYn0Y5cl1vi
BV6bJZqcXfl90S2YBjbBrLWuVEB5+TMkB8EhiDkRTGAH/jMN34eZe1nl9DaO3bNU
GHG9XP5T8efz3ZldxghQM59E4jJZ7i/kgQT5SKnyt29BvtAn6AgTlfod76Tnot2y
sVRngxStDN4vCSHuhrgmHqYuBtQJuan9SQVCHTJaBKXqosuMKEAS9dwtKXjZMKMR
BLhNodAj/g4ZsDWcNy9IbK1dIUmiKUf2XCJWi3ZmzLdDqWx5+1GJCOBGo0sIeDt4
veQBbYrxkWPCz5aJNvy5qZ7U4ey+4IshMuwig7KY8V0gqMuXXPA6GmfrLPueYX6K
+3Opr3W2SZEyvDUowTNluxVqeQYuQxvWhqc6XpSs/HkpN7yDLv66K84WW0k9qXvt
qTiCrQIVmc13SBXn87AjtpaTAoYtN/43KzmAAgJxT7M/UvSiG7lSRbP8XY3xVl1A
fsZ+z2Rw5wNkkg1FUrKrTDbg6ebBoWv1iip88Kxo7zD8JWsB/RqMJk6pjTbHOXdm
XXgFplAQfFlnluGVV3+D2JQkbUGfB5vNU2hcot1c5f/XS1S1RIHPsAyvoTBg8bOR
r760UpelCLVow83AuLDXBnLfs3E5KJlTyfAzzlGt11uRJiTooNMJ6k/vm+qfodzq
3Xmt0QEDSvX/qqHjDwQsFAiiAh77SX0qGJ4N9qPco44v2McwuUxrjaTcJvertSQz
lfGEQQNDepMlR303aakDwhm122lJktPUwUm6Zt0Dvp//fKaqQezn7jdRszJ47bP1
jM65NncWNQ/wuLjEU7septoR4K2TD6XZbiFxw3ISWKr13LoMmkQrrhtKQHdN25MS
FmQF8lbMRTw4aCiDbm923GPCBmkQa0x318tKbwBjhPtj7FYMvjfK9CHunLOP+WT2
iI88yurt/8PRoUPrcCJ4YJvaOWt6vDj32lJeRKctbVFsZb35k5zBgEq9lbGm5LsN
0qjqcdguH1hTGWNMHx09FNAPQU+zAbaVxfVIoRnTumLoKyOeyQDYAdNgSSSfYP0h
KwCJJMlLIgPWIw1cm7+5N6r2fsI+NSFNxXeXjkNTXVQnfm/wusieL0wNUVpRFrLK
q19njgXJSvw2qGi5leQlj2WyKMs0x5O5gZAH+gUI46NRt6VB08y+FPgHM8i9I3S9
ZV4KL4hRhWUJUodHowNtsxuC4PLBv9ag3G7+rMXergx4rpEDIzbfYnUuHvjy0bSf
KC7A8urr+aubTxnt3mCGOwzTmFunoSG4XBGVBcgfddd3DLQYS+Pw+RrRxukfgyS8
pzjDKIL97QdJ/nX6P4fvX9+C15H6sg39doFzYXG6mCwASrQsIpnnVxhu79xVjzrE
NUdI+WSZhcgD7hYvN4Ufxr5AFFXiXL2zJZkdH7/vU/sbkLlLDsefxUBIzz4sWxDO
lBDYUhx375fnEZqaIHIK5PHSKbPNMuMF7JD4n4quP1QQHxhP/JIXC8v1kV11nLuI
jEakLv16FxRoxzOK3pqE+TkIlUAoEiz6BbB8kgr6QZwAcReI2eJS2lhDlycSTgj5
6inVkQxWOma6KmFFfx/Kwf+A+dpRIqW5JisPu4f5HdnLRetoi1KP9JlV+3gBzjJj
MqvK4yiOxp5PU7g3cXom5QNnDYItFrm60SZpzd0ucKnxv+Dib/s1bJic59EBerkr
BNN0JUWpcVkEIj9DLl3H7917q7ynczVnFK9bDIhkZ+vhp3XDpdWYYEKOQ/SdPdd5
TYfIhEwCr8x/KDUt0xWGGkXgQjMilwG2nr+BFDfzfaC1w3MATXxbXcKHKd9le+Zq
gSov46MKdLnKSM1IssayeClxqOryvjZ7Sxt20Ya4pEU5RVgwRrF/xjsuHF+5KDbG
e10LdHPoyqUmbGVjYj4q3diKxhjd5rzVnNail4ffrpIXwNbx5hyxteldPi7+Gf7a
A81NwBLGpysesHW+RWhbhKnN6x+BYa9Djba5ENyx3WSsD9728RNHwZauMKe8DpLB
kWVsSgeKBSC1NFigaWMZ+2pu3ZAjoSTujp91tJRNQ2bW2f8wVC7VmPN4D9wjGpBb
kDKeHmZ191yeonQsnAAhnEL1TD5IHm0FE+lIhamCmYfKu/Hx9SUguUMGR8VBt2Ys
dFO4hBcWEaOHtukctoJ/afI7L1Vd5ldd1kKVH8tXTx1//2x2jIKX2mq2TzLkleCU
FMeILu2yE3OGErOGVKfylq8y9UCe8DC4YYUtEAb6pnBGeIQ1HencpzFDEDBuBrjc
Lb0uvvt/ow3Yqsq8jlfpgp6neT2HD68/lob+m4q+Vu6g9joITWE6oABehpsrUpCT
T0D3qJNQL89vdnd061cgW2NhpqcNoU7al1YU4+iv5acJesdGxFarFixBMSX62yQJ
CoUTylcARcxDt5FkEy9kq9+Fm7md2RrmV9E3NWpGYSuQkOcVp2vxcr2ML6z2uvgS
vS99lsqYNX1hBv0piLvDskv1SIs0ZYKYbgsw/SYhvua6Dwi6WSfddsWBrUwQ1HZi
hDBd/qCqyU7SGJ13vOPuwoGbRZVDyLZBG2sNvourTbkippRSPha1d/fH3MrC+gTL
jR1wHYXE2LHYYhrvy0gJqQkY3NwoO3vtMfRpXf2U+I0Fer8scrlh655UP+xuPMVO
6wiSu5CdlAsblH1eBKwRmCx60mOhir5BTCF3Lp4f/mnX+vg4Nb5dOCq1rY7uHa4E
EGjZCnR7NJCDoAhzKyJshJb9kQKZxDNl9kocWtYRtCqYCZB0V9ABK6sFGcjZzHxc
2oCHwADpJI/LhAPCYYtg856PQ5KnUo81i5xukeqlL2oeQ7Z64gPtHSl2+RtHwS5h
OD00pQb/AzvattdAbybXjEzeqz9PFB38xRTc56ygmixmN1Zj+PMckA4VT/fpIuZB
iqj2d9lh8pgYi4uYK0SyhTnyeAGza3j+OB+A4DEg+2VwPB8hbXfy0Zj99T74z4KN
hB5gCgckRvXkiyYdsx8eDvG46pGZpyX8CjQoojxvJM8+BIbwhRZwvPsaPB1XIxCi
VaFjDuNSw5sVpxskdinDAJelXBMTJRfNyyvY7t2/OU6WQXkGzMQg1gQVrenLoLOH
BVQOH3zagTxujLVx7+tMdiJzvAhGn7el4sZu/VnKAM7nMvtaS/9AEPsGUqdKZd4Z
1utFjtsxHq+55+9ttMDM69Z4BZWeZO+/XaVoBO0RMmyhdESRYAdX7JYNFEdsbltK
kSmLLGmkXiCZrJHs7I4YBAbQY8L/uKO4hxx98T8mQCFK3nzycJ0ruelj6ZNaOWLM
uDCEgMnBacevSlcPle5pZ2JO/cYgAfYWj3UsKCoQaNW+dOqWfteySED2ptdwDXj1
JNEi4LZOn0z3STIG1hi8ZSCCkYi2ZMhswST0t/fttQ9y3nN664cwEwybjGpGC9Tk
YWC9vf7/+XSc9iUO1/2++nfgXpccKvDgtV19m8k+MEo6lTiZtrcCnU9IfmU3hawW
yeD0mCNLFhGm2AsdzvnY3ChW3WQqVo8PxSYaLRBp4H2IHDYAcTUe8WYuq+6Mb3+r
sDYbNSxGHGJSG/L5wNq+ixo53etHgZIbMBzxjSX60MZfh7W+jUq7sPyhmdeEZ2Wc
moxGorOz+nN0Sny7+4wRCjJyuh3ezdsda3fWiWq87/jJTg9yPCSB6BvUHUym4UYn
SahpzrJg+njLCtGTqbPeLQCmbd8FUiqyPHwFhh+G+1m8nwnnfLlAQtTj0z+KwkyF
dDcWj9JNRUy5xWNmBSk9khzFgjy9W8ZIYpL/OqC3/nxrq6P02g0+V+dweJoKAnR9
3OW+FziiUBFg+LGT5ag+bO3I71BfQ3W6D86+cZd3pYo=
`protect end_protected