`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 22976 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/9huKRhRMtvnNqb3Z+UU7TahEoHV+T8U3P3ufru7l1O
3DlgtZzb9QxCbOjthp9+wDkjygH0eUfDrEl1ovhZG62izgEqnHXKLdtFnyVZB+jx
VceOjCBB9PgPO61WM/V3EoFvPrL1BjDWwYxDHyluEr91+yTemnFpV+jebwE5L3pD
F9pV7yMSyxgjzlzKg3Ex0hZw9dI7hXQlAHsuBe9UpsutntmRuza60x9Fqf/ldP/F
JDmGlDOiTyU6wQM/fPZjz+7jiDqw7Z2vOMp/OBHJCSJ37QY2hrGVk78JJaF/tWFb
UOCrKvWczNi9LnUI5HIqusdR1SFA4YnXHvGX3XsMepGfqZ+kYztDB6tyk7YaZW7R
2OH05cfeiVTJaEC5sL0T4sjy+Pip56GiJFoG63sWtO1JJcBIPw3TeToSpGvz0zJ9
YcejfqzlLiFfj0f+sJcJMvcI5GiBjXDlf+TrtexOsPK3Tnb0hzIYozUJy237qBUH
/DRLDAiwXPhBWEh8QzmSKMK2EM+F6skVAQrn40F90OlvJD1/tmB9sDdaVKN+E0cA
zqzqZAt9Z2fEh8WBsEoexaIyCzR1ZoniZeAsoQFbxY0jUig/ywJlJOg/FWM+Josf
kpWnzJBhK/gi1Hv7m+veWg7gH/hG6xw3GV63vxsn1Y30NODyHevL6bFv84Oh7433
4Cdws5in0khd4qqdsrIpxv4LEFp9MEdde+9yJfud2JdHJjrbS2PsvfLCXHtJgp8B
xfz00Gom8E0cY7rnc+9DWkIj2XpmQQI7w2KtUD2tQAevzI+6TT6kd+Vm2ILDfh68
R4bcQLlCda2dmicJ+gQCX4DzWg1O9zKXMlcPExOvHXRJE5A0eR+isfbs9Z+eSuvx
/PziFcqmxcCWZBDSNlDomfTTkruydg6seH0ZdMac/0V0q75sqWKoGzwhmXILKkN5
trC007e0T5hi08rKn72/CK//06qV6w2cDw22esSmJe7HvRrt4jM7kA/6QfIGEqpK
PDgfO87/Q6OkzQKvwEoAS0hkQiNat30X440HFtQR7gzTneRFiaKVktwYf0gITy6K
u6NdILYwCK+rpBZhgLwu8qJduIFxZnl2Omt2/ojDiFk0NmuGaRvwS8lEb73xI+4I
yx/2e8LTzKELP2l1bAXDs/V2GHP6/vF2DoyHNZW1gRrW9cy7p1hvLzEYG8PiKJE+
spqSr88hkcioP8NhWDaLilNid7/GLIv6dE7IyF1B33djkTgBaiUE4Qt6k6J2HWQD
SzQRFy9ICQQtmXBwvR1FRaevTNnRX3+zskW1RMVlg+sLnpRFg78yOwdY0QFfoHya
Zq1a2uW7/nmOQAsoD4GK2tjVfxqlg3F97CVy6drtlnGPs0GS+8Yn6kLX0sw4Dmwa
SADnkvslH7e7PNHBn92xz2kclBazMhOrsciJjRGXl1rI0R0wSQx3RuPSOstdS9qn
+FXDM6NBC4VS52lJjkLLOTuMjjBJLIyZfL0yAJc7VhAWdWsdeLG3l8Szo1DPWt7O
4+9zS4skEk/1D+8Ocyc4t4SR1WEpZwW0l4OmNFr+mGy2h+fpt6crhKERwVA14kEu
rdywyFIQ8mg57QD6NH1EC4YZdxiFPxn+DfReNvucUpks0gO/IvHsXLjNQXb/cI5s
PGNFff/lj9MJd7xpLmAWn9XsFdS0aTxzVe+NCGIHrXf88MKNfhitp0XYRhOhITGG
VrzmPlkB8/0t77rbPHWV8KIuFjGWH5jLnZ+65ybdxsqZ1KFt3lYs6PBsMyczlkab
DOT9xbt/eNfSSMrxlzYySUd1RGxirwVFZ9M/d4zWc5MQW2+0wraGY8NZBRBOOUoP
ZWdxoSh6BjCgFi6Xg0Z5lM7BScDTKk2N50M0/m75DbnbS7mp3Ze44zhqzWGvSkwS
GOc02Ao3eFyFPAFqTdoBXOwacVj5tbPZB6ILFpNQ4izlA22QcdwigKfm1HiPwK7G
iKAP33e9ObPf9A/k0GOGWKMsa5/lFAIBnPotAZCHiSOVoqs7czohfVZdvi+TkXL7
uaYG0URS/7+L0MgYaAIJoTvMVtYr0Xb4mhkoWsBWjhSGWJO/MWYeBslFqaHCcj3U
T/xyWydyAjVUqHBe1PxBAfuP+lIsTayxfrJG4qwojqNPhdA3cCRLYU+Rx+vWgHAW
hMElkk8bv9r3C7qIy8YmjzKMFV7O8lq0jRd1Luu1RDNKfiUIjThQue0PwvDtxQ4W
+uU4tf67DVJ6ynNDR8AGY4pax3FZTAIPNhuJ8lsNUsNdvdf2eVIV3pyghCUcC99X
KzXStAB7fWS3VfrrSsK398aeM9iAYodqIWQYxYsUT9+K6RWAKfEuh06MAD69hQcc
DausaICEZaUAeTkZS2rpIQUd2hyXUi1fYGGQ6F++SpsT+nCmUf0oJFKSjTPck6gp
JbNPD+mbpiIdJMVoUaEsCo5G4QmHSDUPrf4jYk43ivZH05ptbeAvdi5sXoBGOp9d
JMerLedpfLxgT5t/k1ylFWHPCazus2rspY1wFZEOZqI3Uxa58CQ+0RDbUZywq7cj
KgJ9nTm34I9W/oLsmN6MIWPxsMhLpPgb947oy0iXv94FTmH3Grg7NlNTPvwaM9b/
Bz69IrQOOWvbu6saerj7xYPK+uavJW7lZaG8svCNI1L+99Rh2wiPBWF/d8WuBRbD
GUTGiy5N3DyJ0Qqms0eAxVTjSZXkraWL1F2D47W+TDpA8zp6rLjVjgWQ+mjP5THo
P+ZCZMXL1Z6lhMgFJyUedXkftzIijjzDVJxH4oMusWvsCxoSnU/66JSDsTQmlGjE
wku2o2FNUWs56tSbdvAZ0j/5PwBK9px2empRKijj6fGyq6faED9v+6mnMzk6xzS/
/s/r4t5k9PP7DHJ3othZN6PFpjCg0vGxbDAxorSJY8X7+FbY7FSDjdG+tOjBt30c
cd5YKSgesC/chzToz6aLY68AKZjkfG2+fZ5V+xGcT/7HD6KYZw+TBBU9vPiC/t77
fESPoLlt4zyFuU5KjqALSNDNz4TavNns4PvjG1tQGqBYbVYROzhrz9/DKx0N8kxW
N4PcLwsRt5EXPanHBpU4m3Qa3dTePOvQZbXEBPy4IOQdNBSAE4yu5D61jRj4ciZ7
H38rLSwRWClh46qCUk9U3yFYIJI7fxcK3sg5fuCU2XqbrJaniz4yWWxqu3qOSTvD
GLzlXwrv9LYlVVjvH0vfYrpUtpuW6sNYnTk7x6jYLu7Z9X0/oe5gOfTkVZrMuHDm
VIlm7KZG6BlkRcb6hAacAiAp5D4EQ0edkm71BUijBbMvaySgkWsOdpt6pa18R9M+
NzzGyYkFTaQxb7RBLxCRcViOgtdFuPzJ4SX0k+y0ZpI13JYsN6CLAHx7VlNnDrv+
34/MWGbbnlUjlLCXARnCwCIafwjWobsXDIIrFvSUQbk9pvh8xPVm8CbKE65m5BVa
ueJpFZ2kv7PMrf6BsX35AEwuppgpk7myoUoE+uH3reDBCTKdOOb/l7PrHb7iyYIi
wRMox4qffoxc82UQVSK2JVNnAV7AUbpH0KbU7BVJkVawE//89UP+hzBBBXFqn9fq
VT4lqiU1TedIKCst+UVdl4ETf2FbrChJ50JllDyyvGBJovlaTyv5OUi0XoMMPruQ
01lQyB6nrsWM2S6USXk4SOPzG7cIHG5hE3xIbrwAVqGtOsfBjvG1XjgMHpfrycJY
ywJfhmj8gCppXeiWX7TOhut/5zkzgnEEsJlCtejSC37LC6uc80FmVIIdrvwzBNxp
dHMQDd29uFn6+pQjkr4nqbZARFOti6JISlR+Y1roMVcNNMiQUZCjY9uQ97zmJH+V
btLtjrVAQVg0QGY8c4yeqUyqqoGgAEAZ657tjdNEa2BqsXZDGnYj7yr1wcOiAArm
Z5zskA5iAs0O+FvVo9E1/NGGqEzAzI67qfedBHyj84EVg6+xYPxfy2Xf+fGlfZU7
etBp+3GuIzLKSYjFxoGR92iwMBzAtin/yg0E/9n1HKeteF3RgFYon9X/3pjTTvsz
I8W2mOqbpw28TIO6bhrXcy833C6kYLBsrpXfVKcoCzsz83OaTDCVxRdPxCZB2biL
182KfUkNc+DTRZKY6v6mgb0J48JNnwl1ladzaILPAigFgiYzgPknb830mIChFgpK
RspAhtGsN169TO8nQCOxq94IHZ9xxa7Kkhzr9ctWE0nmcYt73vt6FBRAnNO0OC7W
SfXj6ZayE9XHnZSYrEXPwRdZIXbhR3rawGWuPPIJAigambreXUiLuxAbKHX0nutz
sTjzfpoHziqoeVpnK4+LH67FJIkWVkCM+kCihT+ZTY6iLeuit5xTIvoLwLzJQ/x2
JZoFy5OEELePpnNAx7oTFG23Ih2oNnBHIcVb2kaE51p48Ww+dY4qDcYTl7aglWRI
u9w7pttQgdoVbFjxtLPWwGWidQ85Q5MaSK7fAW53qfCYO6zYF6w4v46w7+aR0fHQ
Cw132jS9hom4yzIRbceSa3zyKEnhqY3buS1dsGm5oEv0T2TgJQJXlMxY9lt7EjVH
KBYWsxYk2z0TFX2AyJk2+y1yXpq2ik99Yo9zBurTOjY/I15J1uWUKuYyhsorxZWe
B084abCYDO1sJjFKPKb4GRildCpMLcuDZLe34cxVP3tQkRqEP+yt2m2Pd5U+aGKw
7nyTT9LLvwHWRZ+KxtLEc1i+HW0bEw88gX153I+ynYNIolkgUZKMtS5D9OM/nOlN
BkgKNQZVCV2HTiQeb7GUJePYK6LngmagZK7IBR0q8COh1Fv7g6FrpHwfW/Bxa2Kz
XvjA/mULQYzYsaevnQ389j97r4+lDq5N7SA6sUHNOTH7qZAICUppbi6lHD44HIWW
Uwf6HeOA9SWBGy3+HU2QjGi5gegxv8DPek6XoK14k8GLXMrfj6Sk3xAhMR5dUTEU
z6eWJrPDPfpRu0ZYJ4aJP2LFKTuz35/K5iC/mk5U034v4fcLOvowMkFJ1HWWH/7x
qUQowGv5WDImgI4oA53hNs/iuqPprP5qoYph+4pPZKvmMmlgp7JwZPc2m9f5H0t2
ngCS6gsGqZ7YheDPRgESGasSQkq/CF3G0/7kM1p2SIJJut7qwgwAcdIfI7x03HZw
rQzAxNEHbXP8ypG58wcYp+VBXmbXmIB18O1+8Opbb99JRxkp5uGmnj4ONnBRwVAg
VuV/JLXW5UQlYW2COndxoY/MK1lADxnjwVaevg6z8w9WjHjx7GfuBWsnnQzbw54i
Y9nplXBXa5n63NKO0uqwMuxQMCtOYoacvzguAnM2Q9wfX8Me6nxXoOGD89d6FvkB
rUiXi4QnQI9wx95I+QjXoM6f/q8cAJ9TraTm4EHQzhMu5bbbE911xSfwtacWbD3g
9iCjWgTzlXzwjjPzFbSeNhsxexZl4MRlopdFHJO5eFRW1q5ADPZev7apSPQII3ur
cz2QiXDSDG7cnSXW+E01yeHVikZqwaDoGx8F/s/m7remD40mSNtisqAe57/PN5Fb
GCSpshlP5zBWxpUNnuw8Hfg64uJzOHqmBc7ahC0yB+rB/osrB7u1k8CsNIx7GcvE
oj1ulJpwqsHbj8mpWdM2cs0v16NxnIBfHOwQotGytGjlwjVFulOYTlmbznHtpZRs
v20pDLrLmY2mOchQyaRFPZpy9osMENP1puSrdjN/jIwOKvw65qwQEGsh+6S5aPKH
U0/p5FusNI40S/IX5jAmjSiTvhZfQ2BQmolpY1w8M091lmBs58+tm3WqkxpqZCqe
n0VXPnBOW8XqpHiqP37g172tZOn+KCr6GdEOzjhGTRV+f7pBK/rHD4tRm1jZ+/OU
oj3/LJGessWqhpEboI3YNnM+mQ6ML+L5Va+N2PgjMXDYeTCiu5Te4EhzxwG7SDRX
29py1KdgaOuFgVyY51uwnq4z5p3EObI7b7ekJRti6ZaBG52KOx5M1tp9Tz6lXzOZ
P+WPtsVGu4xl8j3NUayMnLAeprEGhYww8a7gw152wxYvfkS7Rd7qUC6oLY8gJuU1
J7O4CapXv5QdmtNZoGnOhrgh3QZ/e6dK4Ukrr0auXrtlDcwnnMLx/GdaxyDIxgO5
GhudN/8sQNRMg3kaRw24THcZ/lxA8RPfG/WixPnaDn3M0AL7uq6Nu/Vx/j7em4Df
vhr1+4K/DixA3UwSq7z+wkknbRFzgiIp/92TctX7Rm/RK+9HkVf5IGo1CVHH58F7
Q6JuKr9xgoSOKLS22LFkbTz7im1DIwy2N1/N2Zpz/UcwtO2S7DOV3ne48pmehSBu
72hHZ8KmttFZeDmUZx3szHKYEe8w1ThfElFxTErB2GEEMHOrDd7r37g73FXmAUuN
Bqbd7Fg8pOtbZybQr58nCo1Rb4xt5SB4cGjwLD7Fqpco9mSIZt6Y1SqVGpiJR7OY
Ir0+7Zk+uzeug5/+TtPKC28L13KT5kgPSvMp1CUZfChZPCs9FubcX0hmzjOj5x4n
rZnWeI4hLz3ZBbn5DJrC0CM8DWOnDfAfWBqVJ9ITClikX0sd934Z8GUIDO7OJUFM
993+3wdal9LD8V4OTUTB1PKpAHcDyC451kdOH5iCj3Ji5yO8meJhMMJpnDSysuyn
9QmH3sGUKNnDjXzGxGlvHZPHI31084fIKV/7kvfpF93peBS0OWpU34Etc7KBQ0Ef
R6ItPqnUxwa6m8zgtok0dpiCCD1R0rHldxg2Cm2LcsV4pmahMPwvVEZ7nkR9HPl/
xB+FA20tusfPRffKBNMKJ3mAEZiIpPBmEooE2SiNuYGza3OlqcYRbP7vE3kVGPGO
1Ox3dNgBEYvSc3A5psamilnCcSWy796UWRYizKjXOz33rBaNZK4K56jjJHKv5V2E
QNlir4tPZoKMFMJuasHIp+4r5IscmFKrrRsQgxi7a7uUTWQf1rPeLNk5FXHSL5qC
3QyZfTsDCYVXFRYLym1ondi0vPG2rHrlBDTBbXQMqHysh/VBJ/6IFUyVFdC2MyHI
eOiSnuVmMJPhBCa8ipqMUQw5SBkAPr4NvEnaXZbE0bUfU/NjhoSmpip/tgRQIqAu
NFwndlfahkxC93LMao2y+fpS/6lQ23kR/e8/XaLUGEnvp/M5GpfxAHxF+LPpbrhy
/aw1ZeiLi6gbW6P6TR8SIVfFPXhAUyk4CfHTdS3OvM3KW1TAJlgvGBxLsZ6cuYxs
JhnevSVaPFaJyjihVu6DF5eGr/NohAhVHeMy+qGeiKhp92ndxJCJAhBr6+cHQ5zY
z9SecHEo1p8A8U5y3NnhgoXsKjI7SRJm1PPALds/vOHl9babNYzMb4lJsXYkk0wG
QxKDMwq68Vg0bw7qJy7VuGC0wVebXdY0AuPglr75tuZgYZR/W32LM2VjgNNuRxEm
UVpIFqPuMrSlmMQousY50Gk+8YXGfk3uIvoYDUGdiFZMyPg9AhiM/G1v5Jf0n9CU
SMiym1QB/UIwpsDNMY+TsUfhlB/AYMAMygOPVXi7IupTwi3fwqqBJdLNiLs2xLDw
J1+W/nEN8SgElCDoZTa4E2ejYrWAanNxaHNcLyF/Lv6//nF7IP/rQDtuqzaO9+NX
/mnXldTduvzuy3nYkXNP0jW2MPXF8iyIO4B+Pa1I+apP31tghX6zQMP3skRjJ6JH
yjzTg/YJGmvvpvfCQphsKXCBYqPIHrCU6kQ9lFeWIx7Q/XY0R5fk1feYPzgw0Lxy
UBjszdjjoJwCq2GwrFoegze8PMZAUh9Ih5K905Of1pBzcwtyuPHs9k/bIdRcswEy
t689aOF4H41SrDoBPwQhbIOjpJm8/GGB0b6SWQGsFtA/XbqiOXqu3oxfQu1QiVL+
wOLpmGLKjmZ0MAgYy0lckArIsGzrCo6sL0FuitAkJ9SODYGQeTGEC9LbVc4X4sWi
CZE/c0uQ8zC0VViQFig9uAf8IGcvjDlrmSPdOPIHI04wI4ktPJgsw6DurmrJyB6q
79mjsFmzc6rBq+yt180stWW0Yk/V/FGuSRh54TA1SVdU/z93c27SpqbyiPFdWwqv
aMtf+xlE2zKi9kbsHxC+ur1vfiXEbOXJ7VS7p6qOkYQIrQLtb24RbjPP7ys2Lmn1
edjob04TYnp6OCH1doqGQ7DdKfar+kX1PA5Xw/594NSmPw6aKRZwZ9/AAH8a3L23
K5RbSfl128XmGk59TLPz7eRv+KfuhmMpeWaTBKL5EiEfDt6GDFaNMtfKDe0o7FV2
2VTC4aGN6Ex6n/7M9IUu/kYY54rnT8qdqi/vZ2ZZll3ZJ4zqbmy4PeMhL2ieXlIB
f6jru1lAk/gYR0Q9DAy7o5jMWgl+Y5oZlsZLzzbCwPiIAZhrEIymrPPtMIGvVeHa
URibj2tWdv5jZUGtheWIVKBDwZDyVU3/99by59jGEc6jNlZCR8ZJYw4i8/QrGjzX
evqzeiNTwJnG4X4ThaYISsG0rX0zPH7FnXVYimkb2g09Gq7FZNeLBwjCKnJ9+7Up
URX06nGnZWSCSQigrwrHgXXIRkgXOraJXbWc0B3vsOA7bF8U6Sm4OPu5PYJZCGrV
UAJMth1JBO43H4qoYAo+mZTVtQAbrsTvYRrtmXtdriM/BLdHHOXwzZ6UhrfN9Dq2
5QVezFFb7EX1//Ya4kJnnP1OctMxcge7k0WJZUXexL62NzVAkGGqr3r2SMa0c5wo
FwRJqGlq28rKmfaQeRCywKFVzii8dsMyCwZY50/vcTUa4QpW20usan8iiRmfyYt2
kEhXPILXtJEr9TV9nvZomrGE8MdR2XF0BeJmYbguuRY1DjSTSx57NCDxl0GryggT
+AOQhf7MJtTjbpLMYQr0Q7RAm2lfg6VxFgmpWun+tImgtaIbeXAOTbIRWt2hl+yG
dxowgU/O6RjMNVKZwzUIQ3iQI53rilpzSWsytutq9bhCLWWYViJ2TqvdOp2JJn8J
6z3H8t10UuXrp+NH50Dzs0JRozyCqtc0emR/B7Oew1Wp8S6W2dK9WLGFf/rdcqW0
pL8b7yr9dyK+o51KtNY9szGEbolyA8089xkr02giUPv59v1K4uxd2TecL5Bm2k9P
M+HMNjLdl3OrGmLGLgPEuaaWUxlI4jKtAUSpAw1t/QEadGG11+bh9cAiv5cTFcr7
ciecDHXxnOymViqXjxsSgnnynpSzeowNOrQZVuj/iitS6uUnaRx3qD6j7mpMwABW
9vXPzHzEa+Hgmeu3oFYFZfxE81feSd7k7CmUipa6FozUfY9BEpPgzN1e9ujd9Rc/
NfFUfwdaf5RgtPmPytg3LiYUkFxkzVRXtDMDj17TpWO3NGEGPdeyeeKmPFBQ42t0
fqSV/xSDlO8UaSaPH5r+GPypPlGMu4ssAiBLV0zPm+HuaFENX9Fm5XL4iF8locl5
TTY4jRtyISabv/ZDkKtn8wYpadx8X8XMRaHBC7rz7NXqFOtEJRCtVph/zv++Rzus
FnRt+ddP57TIUN7YOtMjpauk0GXJVGn57WiSD9XpMoPEHDtMoSXDbi98a/J5oBFK
d/5adQXltTxPFeeRJ4m7yYoS6jvDVQiBZf6WOHMTtoMPapXmKfrl5dckyWjuRxDl
wA5DdR7KUa5Og/fWCkOmQ2ZfVBOUCC2ta3dLHMR3PlNkO20wArOH/rJOSvv1nw7T
iiQudimWeo6X3H/jWQTAVwWClw0q8DIDWH+IerQE5OipafLcQJHVh+o/qb2wRUj+
fq50+F1SMXjCYsAvtoiMXAFpXclXmSRzF5WMBXYwrJdPFljaKWxVBtfeP9VJjpii
QZhxYM0LB1P+oUL2gibcNQn+23KCYoyuXmMBbO9IGgYItvB4PmL/WFGDxgqn7nS+
9zgkHAkuuO2B1O7JnGlRJvc+V8fi+9oMLXNNz1KlQuU0XgjiM1BLEXIVg3emVb6D
jxXZZG2YON3NA5hUoOyq8aS0EHafA1nr+7yePUeJvXRLmpxDaMPAfuZfYYZyCUp/
AU3VMSLLVpyryvYFs9nWGaSd4gVvVQx8Z8lHTut5cVO4dvaKwCk7sLGI3JcHSdhV
JNt0qv+/5RpiI8iLPLzGRAOWpIgrt2jFj+sl8pX/Owsukr8J414MfRUmwIct5PBK
rAeWQEOMIzWx7SN5YvbLrseAG2RCkB5W7Mu+V3pfBLVFl7kgzMiFu4Qt5gHe8uNM
hzA2gEhCZZ3HpTkk3WQohIVTp3a/A3eHEJj07w34tgvfmgKu7a7VBiXCuB8sNc1s
tJG73sNb8VNOBX8WqVSTIexAQzoIzgt8pzCqqZ/1UAVhKuGrqQGqdZUFWDUWiq6q
MfQbsZeU4g5Zog93eiweNK8RchzJbf9cQnlPnRiXBpQNGAXNpd3EHDs/DHfSlqvy
O2oK4cQ8cPjYoQVBEr4D6rpgLzRvWr960KoY3sOz2NqR1Enyxjg52paI65D1Juo9
NBslhEbPih2N22E3Id6vZsmNXxeHv2LQ/fuIci1voq3IPmn0J5sNts6KBzOk1tLb
JifXd9YN/7tue0M9BVzA3kJokiSKOtL+xbdfU4+n9g/N2fpegYA5iYqUYYJStJbQ
fG4D47Ni7ip0T09MUux5C4K0P+phVFoKEAMbPPAIJS6n8wEtqan5T6D0ZSRrUKCW
xTj8vCQ9Fp//6nnTCGwzHJoTWXX8pxfB2k343XaPAlTmTSxlpFxrV22nMwY28Q8U
t0Lc/xJVBpHSvm8jiv8jAazHsgpfk1b1Hi6H+5aSKNKBZNHxEIAcWGYcGAFUOdCl
VwYdfdgPl1VA7FaFh7KkeH6apuNoXw8FYFv+u9fg0UeAi0OR0GN8QKxD2ijmZTum
Dh7R958gTfuos9FuLHUjhjcBzuh4k42mOpYdEjBkDwU3x4NbyVY2bc4sUfkABzJD
36+L1PF8qsE7WJhDqAYwg4WweX/3VGVAZs7JK2mXBYFUI8v/wMhrVLA+R+uaXrvS
JGE9TZTBy9m+G+yfAnQCdzUvI7bEAC01lbeI82x81ATFjb2sszt0xtNqtDWl0AgT
YnrlVmEOnrkmCOpD/2oPCGz031CDoWN0m95kbeLL0M9ai3TcjlBy6bj52QDJgntd
vfo9zRKIdyLpXE3qD5aDespqLYOofeDHIbWC7VwJa0rUu1IqsrVzVYjSa5bjrDOi
EfUTCXySEVrSJIR7Ah8YzwdGx+2gkr6ibwbWEbT3lzYbGw+l1YI4LCiMXqLnnTOW
SfQf+7NXCy/eNzouItmNkEJ3gR9sfdZegN9C/TMhM0KP/miPYczVcAqKEjPXwN/n
Yq9Vh4hUCFEjqc7bTbM6f27qUAb9QgJeiHBawZHvAij6M6+zeLiNpcXX7xpNuVi9
WpDPyamIw0yGhA71T2Yyn+pz7AqSDt/KoARlLgAJ3dAlnEAQram+XKhG5pNBYAdC
iSYLT3kfjGF5YRkI1dxOa+dkwRFYgt4VBOEd4F1qsq8pPOe8Jhr818RO4IF+H4Ky
+acYFtaDxxtcEChM04MRJ0DLZDczaQ9/HafXCItGyjZo3VbhGIHPcNIUduZnsB9R
NC/FbrHPd3sDPrDVeuUjCvr9b7IyP+FUp0OL8Y8pqGu1YPsL0se/QkseVbH7SwE+
qdc62/23uaWIi7n/l0FmyL/eMzVhosgOhj+9E3v65PPBUf7jDzUkKp8jiqnjhcOJ
VhcGvl6PO8551OqpLsksTL/R8KsDCwVNJWGWw2FWbz9l7gMpubqnY+RgeNt1Sq9c
HSpqjFeQe2YQr4NpgcKqt+uaLgMYl42IIEBX5g+3DJR4m+gTIwJnE2107SXYZx10
G1NmJny+/CNHk0hqtgoBirdUVz7zo+ziJY0FWbp7z4n0ORhtNmKwg0ewp8R+8MTw
LQ4Sg1gU5oXovEi1rDPN1zASZatOESLwAKMorwtuGo/9i3y+W43oMrbh45kOPPBj
F8zKDd2blor8LDNyg7j3YCslRCfv3st51WhwRyWYedX3L/92XsZjh8iJAbbVk4Cq
uY7/po4yB5cksgzys04wrLIGyQmJXb/Q9TOo23oiOgVtIhJwOTA9p9ANBh9JGPs4
WNQVODn1pwT3xkB3B+0+12yRmDpb5LsZuRk1lGlBTrWZBil04mXLttjn36q0kwXz
fSZLxn8axactsEgrWUH5FXsbd1FcVpYYQvLolwCxr3OGgf3oMKx+rr8MzPNjXIfS
Tx9TYp5LR/cCgptAP7I90JIqU5FmltPTuauBGBbQeIz4GuXZbUPqIFlQnH90VXkZ
yesAeraUQN6VM08hEi2sA6Vc7AkGiLyAwUPjfzDcOxmTzD2EqJsVR2TIL1dQ8ote
EdPmP3GEILhwFgxSFwMzfyZjjk+a4nejusEE1yTAdP58gEGXRIn0qsaNFiZxspBo
E4nkQepGjGnuub1TSWI2B7OeTUIbgeSn6A8OY+eUbq8gV6r9m+NEBDIt5mN7C87p
V5evdjzLUjE9JvnlpjZuUbfpBOYG8jiLiAy6JfBGZaCRMX6w2/68uATS0t9qIEjx
1HpwZT4O3y9Ww1whH/ZlYohsmzLvCqD6NYwX2H0hG76Aa0D22AvczcgvNvDURbru
2zY5mLjMtpG5evikUbXo8uHHAxSmcApbnNtafE4D7Up/f26fZlo3b51y8hSHtE8e
vTKgRUlOsl8mr2VTHfAlPkE7U5AAgU6NZ38gc3Ju0tK9LyIIPrzBB9vnoNwUEp6U
lXYSGayLQoUo9iZT5rdRhOXsaKhvj6rTuOin01HwsX7MXSiprF656SV1J9lxNDFW
3BRzrSuE5xAbNOwJxpjff73ddbFnwJcrfTp/0vFxCNGYMeqi7RQN8+222CwqNyah
TgiE+dDHEdmNZCwKMbuslZSbcMiRi6Nv1M/c0sGpjuyxfaXdx51S3zIM1+93b+8Y
dn8qaaA+L0XtsdgVqHTOOZ4JxAm5ZjPd3Z7oGaY2uzo3tQef1mhfUgLcMPsm4Sw1
sqchJndE+wXHw6N/AraOPU9sDXGZ8CTEjI9bXeZIJ26EXRf4DDIFaGznnye8AgTx
/cx1kb1CvK0bJtLAkushF85BZ2r3Bg3f6Eiw5RfGkLUH2eydR5AIUZyo8+HIueA9
5PiyeOHYamaLJxeUIwc6XMjpxBl4E9RLre+lLXWpa/x/Q7nHhV372B2MZGDCIk/f
mHgOTKRScpTVFOeTmfkIGMNJnDglMhfKnE+jKjfTKf4x1AaD4HvNaCOz6/35Hzg8
q54XNOkQY/wivlhZXQTr7HcX8cvp+SZ3oTuvGBwox7IavGaKCyxTpq1EH0JkGVkX
Fr/RFW6O8jJtpyExfE8vFwJ4V18TsRr1R8oiAXcrxN2IvcwuyiOMt5QU/72qrRXB
wsNDW6HEzFi1ObJ+U6LH6Hk+oMLK9IMX9sknIKQUe/u4zXbD6IYAxMZpJ6MjrRrH
P5yLtXqnd2FRal62p/Xg5Z4acD3CriMRTKWiIToJWv58o1Vzb+HF4JwAkitp+M2f
fFYlZ8lF9Ul8Le+vC6/31fEDyJ1DjqRv/ebtOTOxlKloXduYXomlsk4NnaEsClQ/
SVG7+zwpoNGgP6262q5FBPGUH4a6+ZoZQq5nXGKetdjMU2Dju2ZVgxCkh2PTahM5
Zy/WZPuKUzSmfDZzAGBAWZQw3FoGHMoKxro2m3UaiJrnItVMZU1Q0vATvdXeKE/4
hLDJkEyHiPGTN2ljPRg6UlCMRrkddSvgm7SBi2WF24q+umkF3fYe9FSBZof1hxMl
lO/SmJZTTsL/khYdulihHXWGTXKj6cSyfR3+GcVONstnarbu3wf++szmp53DP4yP
b5iHjdgo+2yGslQZv5JIqd1anYF4QYuDzpnvdYsHmSZizeiFq2jZxijm9UfIbqy4
refGsctXVt4LRWAjU9J5r0PBM0vdPY0gmdPoPgnkoUsj8ympzO2B2ZPaSD9TOTyL
l+n3KyhnaCRV9LSw8eaVmHUylD4WE6maVTuM58uNqpTQ0tbO0DfnKxm6yOa7oCGM
0/V8VrIWsnBIV0iIQDb/udpGee679Rys1n77ZY/y4w5jCCkH1izT3g33PT3E3I5P
KtdGugaaMbxPgNtVad5+nDnl7MtpyjsFn6Rljvb7mK79jHJz8U0Ryp2MzmfpSL3e
zrE4fD0rnAi7LBx7p6G4IDNm8uzzbvd6x3tgv+ebi+9XsSTkOqJB+kvPt5wwy7bf
S13K9eGjc1MI8Loazop0uc5/7g0o2zcf7c/OVAyhYXSRSfp/7qdkvKX6SRSz7Fvp
xMtF1C4hPPPx1aOfTvS5EOhuzNWAl2C3uRP5+ucEFdT2/Mj9NJOZijj2qc6SN27c
c135D5dv99WgrAoPSZu/YkILF2Bbh5sPHu4jlN+aouPO2bL4ybJGxF8wyzTrJEyJ
NBFyISaO/AmUDssky9i0Q636usC2No11k7An7SDvLZBZ0loEFF0uQCVjgNpw012Y
dljdvZx1nca23ANyUmralP3YCiH9sPbNYF7++0sK33AsBAQwm+VMKUB/uwbwQLlJ
ZWUakgYCVu6E/nagKjcq9RYeqnYvtr/ObvktvNad33cJdY+0AWYP4uu//Dq5mZch
rRhdEJbY2pVoIqNkogcxjE/k/e1VE+TpY5lhcSg7wOa6epPN5SekZBi7KXkN9VQF
ipvnY2ZecWrqw+WB6Lq5Y14WEPNjEyct7bwdbt89XLPEC0fGDmFCEcFugMQuxwub
TW+VLOtPS77HyUnlwRfjWj5f+Kx0/PqE9HHT0D6JgqhEmMNofNQJDIoapCUodye0
COmyTB6f1BD1o/k+wxhUsEUjhdGz9ZSJbeOy6dZ4lMivZ/nPKNGGs6Xb386uLAhF
cPdNcuqOUh9rtKh6jJ/XvsAdvviwJLPvft65DncGD9zZsCttg96HQV6rQx0lWYk/
CKt1ftvbb/AfLP/q0zH6WS20PJMfUAT5eM1xA+sbj/tB/1B4ZTtX+wf/3ubm8bPP
Wo2Ia9fdjC4MalcWGptItzoNAsm7RN53y4xeqcFZiL8v2FOjB5LdYt2GI6DRpGzT
ZUlnWoXbVkH+6WSdUKbtc/YvFpUpepkKvWvfjVHzZCiEGYWXUi/qWJ6JKfNkVknh
7UBMtLKQvuFN+wmizUcJjE6LcIrF/u+3l79Q/3i8aQWND9s4al5RmzYHJHRRGTkE
3fKYggQwi4c95BUvXAnuqwZTNHcpWIeyGLY7aE1cT/vWpowFIx4/FzG/Loux6ocX
cr3rHGIGfmwVsCSXqw6kjkx5InVHOb/e/BdCKDyaxKMIzjgywUi0cOUlqKHXAwA9
sdxk+HpJO93l+cYu+AX0VoTU1ewRhHCUHDFy02eK0LHFbB5AYL3GAwYvE56qw0ol
rleF6GFfZ8KqUYnKs694JfM1+ACVZC6TLJ9IowW9MVZl2Pt1HDBbiZIAySMnmzAm
uaehh0wPCae0cVDsuc9Tt6O418cQyzkHvSWRMiEXxN+YLwL0oiFjccIkFeEGP+Xw
u7TGbplEmBEcw0fLZc+tirLI/1YArFF/sIo15DQXp4MgPypywiLmBBj7b5uX+rh4
gPZe921B6lHcJG0wf1oIWmJel+WQGmVat9ODj3lAj5H21mpdK7HrEAHfnPB1mm8w
BqEsPmQkilR8sNZS3w8aiuDG8couvCJmaBhnZSoGiw/nzmllerWdbLPHoy8b0iU0
N/rJETtEWCYJ2sAu3yJnbvynNeaWPhZqKBAygaWjI1oS7wOYwfxAKwKjlkRpGXIP
0EXRy4+yAkb5+VWYjw00pCoHg/HQGYNvR+H2zxOWPCyIgfl0IvLZLGx0VR+plYTJ
xvwFN/D3Wbt/Jb+JRPmzDvf6jflS7vEvb8IVpu8bPy7SFfWzsJiEbphWebbRPntw
bT/EGbHmyklEI9GXDhBfN9mPz/r0j8k6jfB/IPesKsvG21OmRGBWx4mCOGqUw3q/
Cb1uEL4BY1Rbsai+LwIn1Q8FxQz0kSS5vPfzaVzCVftC0OE3bc7hZ9iSINRj6UPe
pCfUYoggxGLNafO9Y+0UXg3pZFb7mwJYdueTy0/cdAogr6Q/NwlyGM2/JFkammfI
Gyke/kQlSPQx2xo/0Dqja+nIPoWhKoT/89chiaIqaI50trGOBodTr/wVg+/KCc3I
E8m1ocYMDrcvyyZB8oD1d07RfJhyZ7if+AFUgMktOqOJ37uzRLfVVtHJJzaOP3NS
4pR/zNpIW/yhWkXC0CIzbzqYdEgwQKVYMJs0cnpL6Hckoa+fczEJpdTY40QI/EPF
ZEOeISOaKaBb2b9G7oVfhVXvZooUpoVsUOUcJQzPRfq5Ezqm8ynmAK3KQpI/MXUx
2IghP3EzL7YhNKA7glXFg1DRDw4+cA4FAcPOCjCreca7qmbTz5NggY8do106XN6K
XQVkWKckrnObqnX/nCFiZaj2eQB5AkdYeJMgk3dtMbAXgMY+dVasVCZWdr5Xdgc8
j3SEMeC+54+iqxJJn6VUSzxOEXsh5CCZAeQ037Na1XlzuxMilXDqxSzuvwVoJiQs
Z5vLOAAaG6yXF3iJe9DsBqRmbbHM9xqQXuBqCk33PA73BDRAitnRJNNT4oVq/ZJE
F6eTAiwrzJIy4ivZH8vFJ2GXNAlpVvjwLrwlCLvHS2bg3GnfbgXOQxllA+n/NYry
gAQKZGI7WFFr4I1VvaYnG3Nq1GpT6rfu251ZFV7oqWN7aqOJ5ef22U1Chd7LiQ1g
eaS5A12qf6j89nk15ctPjnHZjE77iDuX9+sVCwwOU1GrwaK1TxWGgTIJCrGNv6x8
We02ml+w05ySyhJBdaG+Pf1ecaBvgjeHVH5p4dbJTTZQDcJUZpHq5lDO0w8EOhn7
yl1iRqLk0NGTGBVYFAjmgecCMgInwUX5AS6vUShgmWqKS4grrqhMyL7GYMrLHJ+n
Jo+rI3p6+2ryciXbXfM720cEP9PRVoCRicULniFM22xXUv075UuPS5unt0wxFe1A
y2dnd6jOyTbTGR1Jd3tAI64lvdtY0oxlgSHnqd/Ho5gc0DLz8EM8Pgw7jUMSQ+Ui
CiRJAf4+yTiedOzF3BxZBLpYWHEvdmocmkWEHhkRNsLgxdN5TQyMDYl33rFPhK4v
eORIDjpRn+xOoLpHzWhl5ZiFVQ8jH4fk806KRSVWVsdVdu3BQRVO6IwQ3MbAW9Y+
/fommpSLTxzqVjLcUgcKfqd4PQINn4PDicgJLkan+yYIE6Woj6AxQIzAqVBLCdTm
gjS+M9U3+4rYMOvf9DA3bh+LEoLcfCNi+zL0RlDPBnMBtNfTTqU88Ezb1nAPDBrT
eiexY5nOt/RkS1L7feWZOLCFA/3KpjZLtowwP+LSH/oPFYbOCDXK50MWCAEOAO12
IpxgRai1OTBpPoaYbAIT+dBI3x62VMvF9wXNbxPjDZlcLxyIG1tGELVPwFK1vKS0
e7QkCxpywL1UMLnPuEw+WhRgpnX26eVOFesxINwgJHT9osVU98mm9/ZrHaEamG5H
vvsZLDiPEXL657S3K0AH1bKYIqvrZJrr59bQwmuWXLfizgAhdyyw4UubLdxs9/i6
TvnRIIF5e/BsZH+bwjfB7i8rsWDLaazTn65CfHD/i6kgmVVj8rktrXyGcyaZ6Fp6
vMKc1E4p3yM2pw7QvXyZUqSfn4qLpmsoyPZ0E6SzlSVM33CVhYPWZiTg7UAozbiD
iUcPPj39PlwXDYCJGOQqIDcBsJJdFwS7jvWFkP1UPSUPF+ChkmI4tTaXJdNtiJHv
XO/ncih897zqvJD3R1kuHVyDvMQN3bEAdTcTnZcyJsWFYzgJGKeoMYicoVAvOtrk
kZkY8f5LXzn1NAlbxRS3r0I05Ug9zLz8GO5SDxSKHgiMBeQ7LE18SMsKdH1CXi5b
YP0FI9fHUpgk6cDlvYBYvbvZQLYUdbzKZc1Xb4JmlAO0E5R4DtsFIeJQuOGwlX/2
T/NQnLkQCk384Vp1cKQlOPlGeDVBmMU24X7zAIBQFl6s3I23Z09swq68Zn1t45ge
RdZjfo+/kGJx8M/RWQoE5YKi5UGRaMnhj2HPBmzzc5XVSEmmbbz80BgV+L2Zuqz3
E15ILxRTpY3bnQRPfVuq/fN7tpdwe91zxswfnLZBbJk96Q0dHO+1uncu2JTuNdoF
RbXlx9WDk8AAxlZ7OpHQ5nsvhnYSvmF4lFgsf9pgas8dg0SzPoQElJehOGM30+R2
wSHXoKZiy9DdTLUGaJMpaFCt4F3pErEq/Q+r9/ZjT005ZqoRjRQjzHrUwBpq56Jr
mG7vjkX+8F0KYAQk9CkXbjXrN4FDmngfv7PHaFKljWqaSQNNMh2yZkTINGGiFapP
+zFAywhbdddWPRRTWZ5XUdXzN41ch3i9wNxpXHHm8e3DIXmrwfWPiD4mMGG6yLrE
XZ88UDPeXHMAsMhrber69+a+4mOxMAElGFU0pPKa3D/ztVWITopzNHZ4HHK6X6tg
aKxAUoQMt/rVOmd9IZ+NFJ4r3Ph1CBClAw2vUS0RW5smrbyfSNlqTanx/axLRGEw
2RDT4d/+niCk381qIrODr7rVzcBcetlLjOS/inGdkgxUozdr7w0OGbdnCAOhEpV1
hv04RJ43Z0pY0D35IfbSK9LaS5FyeXQ4WGqNDZ9jAjq7P3u65D1YGUrt/J+aZezU
jEE/Xzu0KZdlQYDUeI9LzkRI58EPakkImzTms6MzkcMkuchM1iEoSb4BM+YBQgFt
eAWXUCzQR31ZazIki79/PDV5/CvINJfr4s3e3Tdh5KYeOeJMQWdH0qBpHFEmhFkx
85BHJ1wM7OdIN/hwJ4/VzuPMCXMdG52iA/BruQQPisYI90tRdNJ0VNAuUjiNfzRQ
djl49jb/rVIAENGyau80w/pVhqCDKPLeTnF0kyH9iD549IIGfD0GWctnlCWc35RU
e9OiDezuQ+pv/m+8sK00H2yXBEl3LSwBKVYRt8ZYhDPac7npgijeACOJ4f1ECJFD
TF3iQ7TBoM+UGGHNZUWxk4FJolAa+VyNPjoLcifxdMXI+jnzf28Z/6CFS75nhjdD
nby8gPjAgYZdaVsv7huI7A04v43oiPBM7vW/UkcvWL5TjmmuRcK8MTr+Z9AxWe3p
xqYW+SqwTF49P/eXNsRlp/WhQs9g3GKWUhM/oeD1FqLWGeBqVDk+4XN59eQVBLOx
Ztje081Lvm0eutIba0xZeQiqywcx2SSf5/P3yEiuPuUEcDXmPUW5eWYY02XQOIAD
0Iy4sDemk3qU7KjXoM4eMzJ401TZos8EQZyY+Hf9uqQQcn+gmJM9LYMfU6vT1CJc
QC4MR386sQ2eiOJUI1vje+67DsOW+puh2+mjGQFHFbihPZ6eyxsjWq3BYX9B+XQX
IQ38/xZDf8JynHwrVOUFbMe8ob3LKDEOcznTuR52pZWD7rZxlUG+eoe/1rvp0+r3
7oyNKYlv512+Bv4p95B7KnbdrnqYl7kR0icB0qSckSyIhR/B3AC2Y716xpadgLmX
68qgIPXKT54lq1pBPXZEisqEeMFYey4gVzwwkYMfcUO17WDlCtYIvShCN9Q/39u9
5Bi4hbCtSD6WLLgYjAJQiUPw/Dj67EXOBTw+yS71MbbKjqscfFXiNCGOhwhMNfXo
wZoqGQDCf8EHHwdvJD7QgzEnDI5XqtL4qVmjMfaHnPGw8bjZBan4N2pp8VHDaRPI
sS42rQ49LL8yyfd5EeXWFYvwLMzsdLcFlkxrS8eHkmKhK+btN7lrcYnv+Uc7yLnZ
Y3If6E7jQEWT/mpifHBaDoFLIs394snJUTBD1PPvEobnP82xkcBn1pg9cfM9AiYb
pzXOuxVh4ic41zNOHi2X7a2hH5NRqHfAYFX37Dy9yc7EavW1tFb4YO9QG29cZNQn
6dG6b7Hlac/vYDhtmjTSFXrALVXXd8dW9HQJaW227pSE9GZsGqTOFS3Gtk/70nz0
PYr2LhVq6FOMgpvJbaCDVe28OKOQavJtkUd7VSxr6M0a8F6P2ESvDei2lYHIhn+a
MChgBikg1FIeF96w2hUCSIqFzC0imivrOZ6fKpRMPJPNV7fJ8ZO/LYuvMQV+1Xm6
I0BC2sxfReUvtEXWQCUsEXAhxCEpGVOaqImBOFBzutySOoIPltoUFFkwN0289Dct
lXojAkB0WUCEqzLzWQQATzoQw8qmpYTqJipeI0kR2FnYFbLgVyx6hBuR6xC/RQO6
4jXXoeSHLgawdPtvFq1g2NKzlgnzn1WDrm8BV2E+Uxjwsl5bwC/CzaHhgrbOFsvp
pIhnYeEcm4XDVgCiPRISP3WZYPMxdlQn+zkdHPxaa3WvBzci07/4s6d2/wcru1gl
2ODLTu441XYMIjtJe75G2zaNAfGsF0p2NrXO1pIejTE5lcBCdT8TbBFpmt6V+CxH
69QNDTQ3+Pw/xB4RYww/4cgPxNOVA1Gwj1bHkWYljrzbjcy1E+OquiuW8K4NySp1
opZhKDkxtK9ODD+MXuaFgHRLtxCQDC/TzDuRsPeOjB4xWdmc3H7641VSnu8+3F78
yvzjnVs2X549azixAoVh54aUXa0T1+XujQwFzeAP3Zv2XeJQVioz53on+LWXCcau
C+04Law271nLYqxLnjA4uopMsrbRSOoGp6YlB1dJWcKYNtU3mXuHKXXquE1jiY7Z
dXBDlGiOxhyEzhPu+Ys3cqvUO+pm4A+OneMXCcbKVWu39/F6b1Xj3Fm/1iJbPqNB
6uZ164XuJRIa447u3kA63o0wIz/RCMJ3b1TkgAI7PcgxN1/09g1XYgeUcfJpzCX5
5/ddbMfkLOLg/8IeVC6OcqeWqwRr71fcuD6BWvY+BOMcHtDqMZDpSkpjLHIQD5fi
enCNx/CmZlOkfohT7hBUxoSnJy29Kh0ust/qGqxzTuybv4VznL/efWwztSJKe1Kx
Ijq2CriG1dszWWnhe8QlXLecI949DWcT/rOko5nbePk0nPXkZBYNj+cOm2BUOugg
TiD7dEOs1bn1qfsjB6LWUKnLyQioYjwCIctOPf41+bMx1XXGQIDzX93zmW1Q/lZ2
USsH2uXNoDqJixeuvxCC3MtwjAEG8SNs3PyCUIoncbEoiWtiWIKV9COQ8+LjXEFl
Hi9p8B8udA1qEALKT1fYNGk3cmLdrVveNbr1PWcMdLNl/bmpA0auDCR/28gjeGyp
nDohRZKDenAyn7a8fC7pNBNPVH7QhZ0CHH1sA+jHs8JNjVBMva/irJ2b0t5stBs3
tlrF0yVEIqlOq8d+EHq+te240DLerD7HZBqV07FgFeODyFCAqSERQnMSN0gt1dkJ
6vsCJ8sf2nvE+qUnZJhCp2WEuuW/Yg2iuXR4XPgeV82xYdLmw/B3W/lJ8xHrQuXe
Eg9kyf2BjGz78UxJBwlpAMXL9Dimyk4agp+brJhYvReBiPSWH9Ztt1HHj1cikd3f
/FNtAxivO2vHP3gK674MM3d97IsgGalGCfPNxhNOELLQUxTiXuOdsiJUpzI9iJNY
WgBRbZkAz1Q7SupF2JGKY4Lc1sFfTk/Jx/5D9XsyMx2L2/sUPlKN0UI+n0fN7KZM
IDhCcvlj9ITfqAjq00GxZJRi4GeFrdWudLT7wS5ZVydWq/nXX2kERIlILW/wWwFq
2Bk6DZ8BsoUwHzSOgu30ju81HhXBBk7VgJaox+Y/RmN5A9kHarXDj7aAktX8AfLR
3hjkGro1wOj4rUvjWe2uFhd4vdFS2U1jNJ+kqiDbOrsFnqK4n/Z1tE1cVu+4mD3Y
n4UeDxd/q6S6BowclfeGYNZtQRwAbX/WspYifqbrlJhH2WBAT4B5Y5EdlQzHhOsR
MPIDdGi/SgUXIgDXp9gapfW5lqY8msw3KTLrE12o+fTGeeY8FxW8f3tQrvt1OE9p
ckErA53BGP0DSQOrWtxJOJvejU2lsXtEsyuQv1RsQHdiCI+OOIehvVT2g56FmMUw
lO6v8cnzkrLnYBeioo3D9bBbys2zXKTRzofdE7mMS9b2+xOUfzcjCEQ11NsF9dVi
Fcy/0WZ9swgpUI6RYVNyPVZRmto/1jq8LsIeZuMogxQm2EmYOBL0VxK+AjicIZe8
Wp6bueArfyoFy+Rc7IODnNv1aCy6UmS921bQeiYXsmJlfeKKRmBBiYvxa7lsbzeG
k24R3tr5Fom89YBGWXtv+Ok9T+jnVhSqG4nPOu4a7UeXox4GmcsTCDOv6uRY/IQl
v69BTZM5Yyp0w2CqVD5e1gw0rVi45cLvzKTGUx3i4XTHwi5MkAM2tlXaCE8DQlL+
qpN+EcsEb8/SRIG8/kV53BECy1qZgdwlPWjFCrplZGYJqNBlH+fBs+/rzXxm2/HX
DydCYp6BBppbCQODioeTn+zl9eDrenIjRHEHGRXhATdRY+o4ieNUHuic0OEFJ6g5
d3U+yC3Ht34jyNzABApifdzsW/PGYQyBEKseHXKkKu0CcaERh7oklGRw3tuFFp29
Id/Hn2Nnyf1rcUrWd50vU7PWh+2f4HRWPcKN2czqQwyrjIQf+FHyQgIZPFxUuTZr
4q2E2+AHNnXs4vzl9yyK/aChQtAlx8qAUSfnr5ufrUhIznoBbTyybsdlYh0SlDQK
Urfi8DnZbmvYDkFX8A9FY0M2G6+vIAXdKE/uZR21ulAm/5n6VJLRk/358XgOeWkU
F0lWsGdIOddR2IdishG4Esuw3DPO9hKy97kQmZBndVChBIf0HJtqfq2sNnWHrLEq
6d3e2/WREGZOVhj+gxC3gmK//ja46GguFgqQ4W8Zxqa9Bh+eNkXrljUIUapRlTOv
QPglczkqr3HqDPQwQ6QWbZU1IM25ZcbfvrWdoTMnYn6akD/mRKgHkQZnQVGsm11R
Gs+5iVC2aLFfBqu5HZzSa6l3nfW1iF3/hVx1RBlHUdaNmXGgO9Cl8juVeTOCSV7P
hILMaNeenH+TGBh5C27AcM9F63S1+O5tRFKKu/YfbYsd+agxl1+pn+R/QV1Nluuo
o5D3BeS1GiU8XCTZuRON2XRKVH2PAP5qB8E2HxfXl4H4uWuR8CUeGVP2AxEmn2+a
DlquhsAOHOLx4hS3cZ1Jp9cUD1XOat+EsKHcv+NbTSPuJvDcmXNPZivdlcibRguG
dhWWUstZ6rpM+ikkYwe9nnsdQ8DV+iMeYcLCew26qFYRKsPnbkIg7nHWeUISA2fQ
csLWAddbdtWekAM4/IyHwYnduJyBZOu+mjKaMSyMSF6mR7DekoG5ZH1s1K3wqUhj
ffHBtUxHBWvwd4XOWrQHSk9A05ETvbc2K4AFsn+ZeeYSiH0Op0Te0DbPZYjVPSzU
qJyM+Rn/euxnKFI0fokZ2Mj5eDhfp3xadGh1MPHz7hRpKReaB3M0NK08t6vS4mY0
6rnV6pBgI1MTBCYeUEt0dLaW2/W0ICoYrhvJ1oyC8/ocxtKbGE8PxdjrIqmAExKD
XWydgSRHjEb9hSxG2FW4s5EH9wwmUbcX0SVb1U/Sr3hYs8bMXKVcHaTYVxocqGqy
7FKUdMeyFa+qB3k1Hk5GrfrBw4sUUdTK4GCXTtTMra0ONl2ILSGb+l2ssIm3XZGQ
AgFIgAiQT78OwZL2qVMEZpzSIVNU9l+0gyzH5q2sqvm7+tfnRiNcUQBS73HKMqTt
6PevvaKi4pbruRZk9sXGVjqdKbmDsCPlKOctIwiDOZ4QtmmcZUS4qSUCooXmjvzU
pbPSVCFgK1i+HfJM2+y28mCt4A1D1w53GGPdDDaOwEmbYjtbDR70HRU0KRU1JOhb
+V4uX5XScfrMxYBvatQG5TggVZwEy5fzO2+IJnpvTmM0CMU8LxPWaXtoMlimTycH
9w5noGmmLiAQwZ0GX9zb8BtYtp6IvZKcgkSroYdcHtoVpVLwsZo/rhi+TdjvwwSa
wDpnk6bPRfe10oLex68zU360Xv1yp6sU0UiUjaa4UXcOzuu4wtRdmGFn6mZSM6kg
tzEqXRW4gN1w6nbZIff0tbbN4behJnFBwMvSYZbMTsnBWPS78Kq/S0B/hNcKbsKu
IPIcH34Tw5fly12BwCHJ9sx2vGvAPFLXBYQc+dc6VKRYYwFkm1HhadZc+g5ajs5B
psbR6tJSPBjKjeY6W75nrdJy5M4/dERpDOH5dV5hgjpKKuP48pP81TQZ0n4333kz
fBHkyBrrueyg7XBpCmN2h0tR09xEKlzRZ9dv/za2juWV50V2ccMxIEvTZMnAiiBV
IrfStJo5bzcy82kIU3Zrmr8tkkpQ1XTwq3DvzRG/GMUyUS0bgEl4R1ZIo3OxpTmr
GVJUAOUHSAN+TvR3tXDZnJQc+NSj/21DlXULZhWkHzW2WVb1klkh4V7PNLHyRief
6Dcn+xyK2EwvZTtCQMAY/cIC6Mrgp4zuhI7lSDndP4aZD5RwWM1hrQGOm33bWjwo
FyGMhmqAn9i/VPKu8niFc6rkELfEdWXF1AhN+vSjdgL08FsaxfjXYsFoBLnZ37vR
uTF/jW/rJY/NXedX8vGOdCE2FPMGqs9E/+gdUw9cf/0vI07L9rKdb4CdGiaGf2Ds
oBUUJMtp4EYo5CpIKGExRyJUQzxrIWBI2qYgyOC/JBmWTtrG0sbnNjio7ur2RHSi
ODp5Y72/yv4fcUBZ4DwYbj1+ZKWueFOafTHCFHHYsDVgIqY1X42sgH/Ptjnz2l5P
yFvy8Y1wvVQBjmotSX3H1xwUYNIlQPzChUIRV9DaFWg6jiEcluZMy4GZa2ZS071r
L8rKdo8GrLSYpGMbDkPRJpHiKtJtKB8CoDYQMbei/QuTPdpFbdm29Kslxfp7C9A3
fPJ/IhGZsUIdXewYd3ZWyem0M495fRCWr7JESUA5w0NW2RcyhDqxKpHoUPN/JHCu
QBG8RbrBq/he3xacstC80QoFdlV9IigyIJxC/0XnWd1Vy7xA8Oeipih1EiVFJKGM
iXHkmhtqbWyk4myOcW1tUqmH/Iw1/osIA32GhSGFA8rbGbiGi7/X8syMaH3R43Aj
B9RoVdh1cqNRNqcoaKfSRSoG7LueTfSBCkAyW80WZHyLtGrTmsW+BQg4N4y6qzdH
+EyEITd8pqeFV6l2V7jLSxBbyEWKCoJdiOjcCzI3SbbeDcShqs0brKCPDwvQR29+
L9neh4sRZxer+VzR3CDIptRmhsOsit7sX6CLVkoFrjYN7TuyFTImqMnaxOzYN7C1
0xZrhX1ydS2vY9RWflQWh5ebQD+eojvv9AdnpjPR7UHlXKPA6oSf5C8yzboLT/KH
3EH+QUa/bRdeoFYICd61d4pGUMf5uAjTpSSBjQmS+0IuB4vlZtATPCQJKPsz2bfy
ybsJOMgWaQlod1ohWBkjxkmnxBFQERS3ySvQKfd29fsefaqnvNUI3KE+YYmBQcWb
RIv2/WrGFdC1ca5Ny9hM8Rd9jo9OHGyh1VuIT6mfDlEuAnybomwDztzbVm1NRQYV
xpNFzRiCJUl9uphVpOJsP6e7C6bxCHoi+DLxJlnF5qRYHaadNDqLP4pkScVlzBOR
2BU6u+dTc8pcC+gzKuRFz3rzgKFJaBncTpoDCGLVPURAC5BCKDmYTG7VE+yS8lc+
kvwiOo/P1BzScv3JyO9iflmacBPG6su/do4H3Vuao3omFc2C6bWi4DZQqXXGRcnt
RgARdE65k9ffNT7dW7RutlMIWdWCqubN7YZFkmScPlOLykBE8UsD2dhoo/ws+P4Z
jcZxynEv6AGV2NaK5blaB3Pgvx8m1ks+dqkk4E30eMAmy2Xg+P+LAZx1G52aK0U2
982taGx4Gw7paZQUkGd1G+tcVAav4tkua7Jl4J7ZnoQVW228/KOPFt+yi5GtwLRp
SQUc8vzZFzL8RkNZEQirPsdjjE/I67Bxfif0BpBQ2UACpkA6gZ1VPWHmFvo7f0X2
mDtPVXu635FRh/85jn4DCIhsCn2eVCyZOt1fBOWKO9+EQv3AO7tmlEKVMZPRf6RK
vFqtYoYTY3y8Kkx9pz1cUuEm3947K6cutaTNgHdmAe0U+AYF3trBxh+rqQO3Wr+h
NpKprxtQiBreGH/0Jw6u9YY404ZPjwDINsDskcxpAG0nnoSIx5tIryf02nirJ9Pq
s6KzVBVwWkq/+95GQVb49EKYqi2zsBqJurp40ghCyogwE2lEcnsnG1qc/B0GcrIF
CpDilFqVMSBfZroAvC2exPw6cdydziq+hWAUV9pBWOejfplVkDKkXXi0z9ClKF+u
rh+Hs33Ok57j5QvVufphVt6XrVGZtsX+q3CKFbiYRhxW04lVhW4JqUSTlgNcnK80
fCr1OtEU+02u0+xnGQ79aKBPNfLIDptAHy+20fQj1Nz8bMcSBeX/NdPLiUX7PQQ+
nHbhltBH+BFvweGXRNMO+8gCuBZBRuPZfDAoOaslRA9vP3v1UFSyOECdDGCx9U9L
Qzaw8lLFEa0vGjDN1FnP8KPy1+CtfsmXbmNYxJ5RWPuUAfPyVdycpH/a1xtdslSY
gpvN8Hcx9T2rqxBCqQ/faTVbrgmo3zteQbqpUxiktyX+2EJgrCcoLyH/my+DDJ7G
5tP/kaADdZOQmZcbTW0cJynv3sXrkGBCb03268lGuSookGce0IFQCoqAh6AsRSzS
trznNnAkxC+fg7jnSEUAtXCdj7Qdofc9DzvVepTdPI2D20qOLUuH5SaFr6pEkNzM
BUqCmYe4Q1Afhckpmz9y5gkp9Ca4Nn8s6vw62EX7Qpnz3TrD19/lrEB3PksqBBF8
8OeGhpEFysdoZZEPy+ZOK6ridm4y3lhoUlNtug9IgxSKpx8QJ18nWwWJlb7YwTfP
8l1bAjLOM7KBW/ZO0Ysncr5YcacAxB9jPX2l6voDcBT1WGqXIl3YsNiYVcQgo1+7
W+RDBS1r3Q72QyF12tftDtMfCwBWTTwW31ikSLXBsTF01dIuW3O0ehZ9DrdSuVAT
BNxSCQ1LVSUfUtGjpCO7N3BShxm4RFrEXpWHxzv/qZ+ohx8CYDMWWCyj3VvwZ1R1
N0wZWeRSIlEgx2Gmu6tXlKenKPSRfSLJuPAv5ESzc5PQ34Vjg+ToQgE5zcLJw6gK
7pU29gVlMC/10m1SiywU1kFClQpMmZQ451UGOLrTmcmgKdpaShV+4A7uixcsfn7J
PybvTA05bByyI74Qb8Om2qj81wQeJKtRVsgmrkUb+BQB/MLx7m6/MNphJCTE2pbW
y4016bsRd/5BHLDihyHPyhAsPItqh28miNUYfZDjlXrKef8grgdsoSnpVnq0qlOg
bko2LCyLk+x4T4EOP0nXAJ3zUANGKCoJSeO0jyj+FA0UlwdXixELF4W07UvMojx+
0tgnAU52h1aO2jyP2qzUnvkFrq6zBXf5FjzAZg4peyUvGt1FTHGk45xCKP6yETbO
0P0hglRQ2o+v352uXLvoR371bxfHfyaGQYUQPC9qmg6kftdthBM1ctuWJ/6QD80O
V9bKldggnHpqbrRVODnpF3RkxsC2ELMcBI37Jd0BgPnhaV0CFBHhdrpSvpB9fQcW
A1jA3hM2XF4Uk+ffdmqox7xf1MTxwdbkTPABxzOhUH54rHgOS6wtU4QhC6i0UBUy
YqfQ284drSnnQgAQwhnz+o/HKnKUiL6WGtigCus1d9W2hG/YPmMz7O/1/1ABPuw1
xFfAshdMyJ2nuldzXbE1W+MzGsEMpv0VTangjAo7bqICN3sHEJlb3Uwh/PDbWfG1
VLw+s8SVsfonCNKk+GlNHZbc0E/ySHKpZYE9cfSfhXvrfdHrDjHz9l3w4lH9Xkz+
0kOVmt7QVFTrQb7111KSI8TDp0kfeejXEd/iwkYWnjL5mvI+7JFXKpE7HPQbTJAZ
kVxXfomr7zV7oDEoQIB+Pb34rWWje6FMKg+KWS0LYd/H8n2I5T7g9/wDCbQTaiN2
/5GJyqPb1WY3rzqrygfS+90dsUFIcxQkDG1uaq6KoREEbuFGWNbylGETTuM8HC3E
xhGyrvYehagxLztyPtjbtepK88DZ0KzyDUCl3rvoqRXPnN0f4g3mipa9EYvIZeh7
5go8RFpOGwyj4NGV3Yfh/qeGOJcxjCokm+j8bowVOIfrIv2Cq22r8dCDQJcPD82e
K7spg6ICIX7AZuZrM1LP9Fr17if4XymWVpuDuxP6dppa5+063Lus6uOIq+te+hSc
YvxXmpBET2Yp3azuutEjOREtm5DvXl4OPnKdRu74iZsaPyOqENBz+IHS7ON9YsMt
977e0wpdT5PfqqNUITNFRkpMMxntj2nUXVbXtiHeAPB94KvkOU4X+I/klNFWLxuS
bC8JYe9YXJQkqc4HGItiQGJoIUlPw7ZrbTB3M2YaiwAnnb7h0Yvq36yLhiIu3bct
fatKhvBK3rOnW1akIt04h5ylCYhN1m/EWdfJAkN01hRFc4hq6GtR/X5YAzByQkQz
e0vvo+PKVZWKS9AgNkmyQge51Y5QEUZ256gtLuWpXjSVbiYqSxXImZE+brncZBcS
qwujaKfJhABGDpOZYGSCNsoE/irZ3JnimFNq40S0gQCvbOFADNEd/45iccl6+KRb
g8d48mDN8f1uUE16z6vPw2atl2vbSTnOv3lUAYPKpfjr0QVXvH7SGC4ApEqbXxPW
uJEZduQJJyIXYgNPeWfBLgCDiikNULNMuUGmeGkFztFNlTli6VJYr7HpPUPMlwij
MD9gV9JQzg9gFff1QtKsZ6b7rUHzwCT89DkywU2NMiCh7memmYzw5lBXSq5NXrUv
15lplpumKSAzKaF3FE4sMtVrY0gZGfVbwkJaCcbA78PKQf9iHhCjxNdL9hFHSgCJ
xrpi45+t42+S97T3gkJXZ/h1GcJhQnuvkP4jl9KO3Hj4bwaaxsStck6Qf8FMVioG
893NLkastBTe3TXdeUTXv9Eo/brU0onoUsMEEe6k0spkD14Fnua7z7ODzQLCtTB1
ijecoMpGXY9+qfYerUNzvY7VDqqhzkaxvoqvgwt/q5ptyh2wgmAdzCAh6VdflsCM
VGMM0kCIk9hoz2XBMOSoL784EOUyLZJ4eKAUOf5Z1n1PbKamROdWDWJAqECFCC/F
0aXOYMf8IB3SjgM2Wdm14LKDE/SBD2jlanCVOtdlT5FUiKwO4A5veS5tL5BWRBdW
0ei1GdmMSu2FhEHgNyO6EJx2rnBQMZTSxMoDIVGu3aEf2zrOAX635zAPw2BLgTAS
oFe313IU/vJ6EWoo4uZrpvL7Ul+F5CCyeLHe9m3cgnC0bO/0+vcoHD1nLSSTq5It
MXFidffxMS1OOJHBvIosTm3KoL11YavXGH/u73TraVm7FLvV+AFImrKwOp1qtJqt
VYS/mrMjUtlcmsfjfOehPtReodUrElmUWXqBMJgFWnEYn/hsntIKEHYvFjsSB9xa
RJQIWfm1jVrwJKqUHyfHq562lJY0rSfoAA1S95EuaC9hYB1Z4J//Rr/WBumDAi7h
EWBVzRLtnXB3jNQi4Ld0a4ERyVE+7pSlyD6gFW9510f2EizYm4I7CC+g9asYqxP5
smYEhoyyYCzzhj9AGEJD/aW3mgcoWeYUCDBRYhfMM+V5/08YG0Mx7LIb+LCQsxHx
9TSH9OFLqQzlTyvvOK9KDWVVviLTaIjUHo4jN5edctw14CAPDk2js2PCj4dJiozp
dFvkd+X9XJWU7dvik7E+VauEvabfSut/3cYJfkV8jxY8q6+WMlYzMWz6BpQNB5kK
6OFPJV4dEMdVG4oGL5CC7X3x+a+hVI6YdBs0rIVrFbKLiMJr/NL/ZojmcPSSwGn3
ldDrqSJ9FCq1hNufuasvEHBAyBYoSp0Dh0uQkLxcbVnZ++I8GKX7WCFgsqYYPSvV
rWxWnvvp+VtGJjar+KZSHOMPbnW0+NnwLfUmHPx4t4Y4QT68Bh1MFRVvvisafspf
Axl99oXDg0ys4VoAXchT4ZFmpKJvLrd9/U83aTRdK64q9aUgh9NbheyBF7/2WvD2
9RzBSLIQlac80rrsBRIitppdQ/MQx/2xSa7FeVRTPPZgJ0tB5z+8/I6P74tEnvNP
e/iNqoDe1pPANhb3q+UcT7AabV5ODzoJSjBJTZaP5dWn64CYwxihdpIkyNXUxzFa
xAN1YOjCE9QK4v0eaPbfVvm4vbvkGgc2u6lovx3MMHyy+spcZXWPY5JbHWEUlmyt
nHZRn0lzFbYjbANo2R+pcshpKoIxfGSjJHpu9lsJjlaT76tqS1kQ/F3Fd1dLYZCb
IDQkJgE/pAfgX3goMlFbQrgcxKWXp3id81KymHtbYPGQC3bAZ7tGqHHN2HiuVj41
IfZeVM679msjXMe6GhTa1lWZx6jjHQaSsTpxkprhxkD/punEf5zeUagfXeXUZaAl
Ca7T03AsiYAziQZsIJrZeYC0ck0qGabCycVX38/YQgmAN3OpkPIW7GEK/pTf/iGx
aOnqZoeZgKYxXXzvKcnV7lnePkUxuZYJqB+94xhNGPb6tlwQa5L2DG+jFc9PSArG
IoH7fQShNqm92fG6Xqv4p16XHqU7+AZ6Qo3GkedCiB+0dNC5awuCod5TMk78eoPF
1cDkBuZ4n/85fSfrRnxIBDqonlg2lcwaJr7xqDtHJBuaYykI/Lwsjn1zVTD7Owcs
PHkWBKcmjkSQeD1iSPYf4RmAxfe5YKm3Lcam1Jp5uuE/QAN8tDelxpw5Nw5ZMY7q
NlLRhytMHe9zzuFsDHWR5d7CXirtDKd3IM+pd7sDdmNHamsPaVhxmwk7SbBj4Yy5
E9UmNYNpgsyLQgejtFXcZj8XYqBtA2OnwTKvptWlCCXgOBo5UgiSa07PXDW6TlF+
ZjMmuPgxyQql0zc2FRdtDg0JqtZM9WQNayXorw+KoMzDMHDKnksIeaTYuRnPITAl
EuvSDBSx19MlbeCa1GiBw8+16m+qHIDeqaFpIQZQchY=
`protect end_protected