`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 22784 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/59UwEX+aE7FohaWu0/8IpTj7mav863zUNIsgIH2BWb
Abd9opeuBjbGF/waQMI2vMJTwD1ie1YueHc3nSNpEh4OXp8P5ybZFY89uyGz3ztU
W1EsuUnchJoQgbHZ/sLbgtGRgsrAFn+ZoIeGN1d6RAF2wAESJmYP8zw+p00RvjZ5
heIpmLmrzD5nzvK4jElYdA2BimEnJ6fKwcpNmqwbTz/c0FkRk2RYQRtVPZ9HoAWh
8a75plMlb+PZn8rN2Q+uoNzOr5ooGoBMo4uBfChHo1bfIGMZkGa5NNZfN2H8FVTt
EKPVjCq/2tNQAvn74KfGwBQH8DyaCzl6X/HBE+tdMiYda0nDuxNCutlVjW2ssgpV
XzxxxcqWKFwlAcZD6isruejm7q+ppRE2XBdHYctPIW4m8i/6vLWW+qk4BX+47NUU
NxzmBG3nO+CEVAkMQbngwOCK8w9sU3CJ+QVAZURT5LdiT8rHuc7IoCDRBW2K1I8M
KMzfOPIjF7tWXDh5Lzaoj4MyGM5wxVVvJYjkbyUKIk2affLb+2OEQS7ouEZWgDjm
TJwCiltsyIdNy8RUL8T77G25eAY48+UDD4N4knFPJoOhhkXoYpT2Ebylg3WMw/VA
yC36aSgfI6UaTi75XvQLzQoqaZh+KLXLHd434T7aXx08DaPG1afagTruzqBEmun7
DR+K8t1oGVhcy3YLZRzp+swSdoqMIUxFAGinMIaCVJ6Jdvu29XH5FHh/wscwd9oc
E+I5SwABZxp54gYEi0+1eFynfuZAODvxb+eZwvJrha4XfmAS1Q9WguJ2ATXrst1Y
Y68PjZ2p3E49MqavR0y1mEZ72Emn3nJksRS6dhPhb3Wg/oTBccKhnVwRupq9Mdoc
5PhgAm3wfVtU3RIK35DFidgd5Lf0TO+Zs4zPlJmxKaIgrb3pc8d1UU1ufE1YdfEJ
QYcxdTQWKs/qvjJOJ8Gr2GQuVQxEsZ0GhAQp9vmiVbanNL6zE4YK4J1yW860E3l/
/oh0UcLIej9CMmMf3dlVhO9Xqq0M8F7EH6Ws4eXVfspP/t6pvW7pznBfT0N4CgP3
EiMG4motgM8+ewxFaFznzEpGLCJHmd+emXXzvzuWVwOCtHYhOidI7Gn7VLQG4IR+
1k6AbAWDPrkUXzIA0P+pU2CEMVdGtUBRO8piyToZe8H2O81BeDhxc+7HTYCw0uYj
k4u8gsFfy5yI46/o76/ljrqYG5yhkQFPcdpWN7aNnLh3IwvcS2LiHr2l0s3lGuIT
U69zz9+ehfg4lFHGD5MVFGIWo117G3P4p7KKF/FzVoOd92bRdx5U03gNLVtPLkMI
nZpb2yBpIbB2NJ9B+8saZGdpIJCypusd+2/WdfvSAyCKsPjziXV3udZSRoC1B6M8
DIhprgKBi07B1QT4QNjZprqwu9k4XUh4uVuo2QKWIWlaqzWRkEmJoTc0AQD+4MYw
fqq7KlZh2saoMpSewovF7cOJymrhC25x1t4XgVpyHhigxJt2ynsdQxZPNjtfsiW4
KRSp8nhP384ugK5SsJZNQoSypY0TDV+V4eE3cbSLf565ABeDqu34unkKJNecgRai
ahYnzhbMRSXLIN96vzn2WtrKEVd8ZkhnFd6+bUez7u+VMhbJWbuezNdEf+nOb5zl
IGk0W6dTT59wjOc47lOfdpit5MkNdZ8tVPVesMDvDKkuuExoj2ujypTZCgJQK2Xo
nsu3sjWlBBXvGrDu5dPl84zcZ0fUW0NU7EGKCzhbKXlNW1ojfKbzwUHYz+zT5b1C
KZPzD6SZqvjmuPvnZLMg1s4keFIG5AejsRZ7uoEQ8UdO2HnvZAIzAu71mrpcVkpk
8PlhEFOriZwtaEiCwpXbVeNFcEWb7AJDxUmDkZbgNFk9Kz3g0Go3+wlc9cD6N51Q
JfUag1GdVf4kkl7DYGIfvEKUQWfzCwDvNOSAl6FznrJTVwfkF+3bcR0DLp2/fr5z
O+zMGWx+Cor5CChwMK2YUfSukt48cI7NWcDFRVshgQyF4MpK/an0SklMF5cH9IqO
WI1SJ8yQQqsHmSwxdP/urQuxlXg5PnDSPxFGeNV+wr9BUJUuyT1DJrSqW3TFjgrW
zJaNefmynHhPpUuEhrXwkAww/NQ8C9s15BlO19yYCya0TaJ+RF44T+LlrNc1KL1c
upTn4bv2ptwLr+8WN6OCpQ2fzswWs7tPDmj+FiwBULHL1f0P6gd1q2Yzzbphai0A
90Aay6hjgWzJ6GDf+G+PZ48asqYm4lf7UKnLOKc/GJEBnh64upvY7zFXSkPQA7w+
1jEj+4gNIFeEY2Z0EpFZoHt6lADyHWRvHa5GtLlQT6WBK109XlHEe81lgbJoiUZ9
M9cGqLomyfsaH2oUxgxSoJBlW5OGXxNWEXEzD3EvA1QRimqekfbYuDXPrcnIxXhK
AHPxcS8FQjhhM6fxuY+6exLB3abymc1qC1L893Mm/532A3Rp3QHy4NitBGdHhKNR
sM1HZbPigu9JjaSmSfDM5l8gdIEPgQtC/FRKdZn1sN5xLY9e4F859a6oFtgXqyTe
VYccTrOtRS8EtOZBnAprhOUFMM8NtLNZc51K+hBIZtQIUigYE5ZFx9yqxfz7aYSa
pij93JAdvGrnLMhg5Wi0jpikoNl9bDSLvb2lV6VWpkrZrSl+SBdcb6OLSiUQVFYj
6wbPXfssmRYlZ7u+CL8FUrT91n/uJFJK6nMQ1fGu0JASY9TCHH5TeJ8+VnV7q9X1
Q3Z01E8hEeCIZO67W3J+iQiruPXxyAEBrgUQqYmb6ii0TlSjJaT6vYpSy8kboFJY
hhi/uB0D+Fw/XDf4elLz67hQPdmGi0nGpovobmhPPP48enPppwCe3sBfoCHKXPhb
gCJQa7qaSH4plclj2o8/wrAZylM6hx+8FQZmQmrjEMk9Z/jC7U/CZFLNs+VbOHJH
o+gmC1aw0jqqxMhwiuSHaNE21t7dBokLCTNV6UQkZ8zPmrllBnrQKiFjXbPl10PT
lyHN2Y26Yzu8qxfgcaLscV6HWGGd13lSe9BsgcBBHlICSTeOWo4Wd6EabjXY6aRN
8rvMtFdLkcc6xTdp0Xn4dF8I/Uzh+73NyWNca4Z/vnyFAepQByDeyxXO9f0UlYaS
5vlHpzcL6WNYie/FLUQX0F3GJ4yYwyzHh/4hVOZI9yVsVVSPjnp2qcseYwR9VAmI
2C5mbz3fh7sn18HY/ro9tzdIjqaLoQ9Sfeq8NBajMphnmi9gZ+WedNUleQXgvuvK
lwETaR54Xa804dCCuyg1cFgRbBqIzwCOXI8fOSdrsDs2O5SJ5kMsVlsDEPnvQutv
XmIMUi+FgH6t04fLWzww2lQdB6gaNtsyf6+Ym+DbjMm+KRxN6wRKR9qUlcRMeNik
7q8iQjj01VoimHSpIDNKcTqSWk7vAr7JK/NZ3D+RRYxVQKHHBU2mGOtHVGRNon+r
MPE+XbCSSzCHVKkEt4u+fzxyNQyQQo6CW7kt5Klk0fGHSmATMgVXeuaSS05OWZ6Q
uHahihV8d8Zb2XTgb1718FlAy+26cW5br+mP4Dw7sArrIYkUJGSRiYQ5urfCRhUS
N73zpVYzlXhQErR9khKNFu4v15n3e447vwAW5Cr9xepgVEYPWB2fn9wDSm5AvSws
D0LLseR/CXD6sAeVSb7fxtZd5W+t9jwtVXAAJOlrG9YZrW0BtJ7jPQGLnLtjl8vF
jvjm688RiKgThqcGI0+rqXN4feEJAQgXJZ89aiI7b0bzZJyyNTVMWo4ju+WPAv3F
78UXoeKTbpMac2bWJL/wtNKH8MpmB2+wghgp7/mQnFVqjkWyL5uS9UMF0Et2/4iu
w2XhX4RzXZtKs/PbpcrIgXbsJdkA/zjBZz7Wp2vNkw/V6VuwEuYEQka3STvRbR0S
edE0YOq3RmfHrsqb6aSQ4nvrbz0QIXfJ26sdGZFq2G7gPol+XeIay8gHeDz9m+4N
jCPXq9Ac2doKucnADz+Rvgy2DtsjGlxhrGZqOJZ2nf/oc332FSDeBvgUlONJcdDI
tncMIUxhXXxJvUiMEQ5GvYFaiZ5kqzf8RxPPcrdo/lFWRDPqO1Uett/RwBe+hesZ
kfRR6NlGkTeWk0rUpCG5dOh3xyzfpavmGSVwcZ7qDOokOnU4xRoRnBWKgXO9YQeb
iPjc2X00lWWg80aRgCPIHT15fRd4cIAwKiaW7SHJTKMUk7NQehiAw4uXkW4pWrQk
gyLjb1ZbtdC3RnzNwoqtZieD/Paru/EmgEYbjAWTRvI1VGzAGtiq9gX7rEC89olu
ou6IuS53pr0PRM32lriBN8wcpkHeb2U2yYODn8AXkrK1Yc1WZtTN/yE3EclXWkyC
oIB14a0rQqFMRu9mPvC1iq+rnA7qo6pGNnSnJErFpsVl84Qcj3t/OZUfeL0wU/vA
1ze1AQra/0JusCUxdAXbjqFh2HECT8lsKWLAxDOLrkjOXkHvX6t3IhselE/G6gRp
1YIcRTv0o1dlCKngmifod1ekwzsUoVbmFqfVLFcUnRFunRzzXsqyRTV2puXzXGEY
/x3fZgcU2ltNWVDxwvBavrIzbvN06z7QtiopMhOqDTkFaIZ+YEm2djy2Igbze9qv
AXQsP21h+UaQ21H1b1v4M4WS3MmJ4CqkyD0i1HaQm21ZtvkDoA/2y9RZx+4pTTVG
1X0+sxpNSeBQ0txp58vvkJrZd86TLKYpl/BnxWNjEsay0sZcmBbDgqBBT2h02sXR
qaW5WiWmI96G9924tpGGRLXYETSMmOsjiv7PJHkVAWnKCRhbAkJB6nple5VBl2RE
NLWRystKgb3qmDwngNG1YnF0ukCAQ9XiIYOmKmFdg1dkjiDbVw8x9fDfsgEbPSSj
RGMwRHu1AbZvwfMJtK+Xitn9YljtYEreEr2Ho3Q1cZXLsou2n0D9BbcNeX/fp0FN
yG/RK/KtwBqSuz9wTd8PijsbBk4ATJ6gDcu4Oy2RBqec30iWdWut8eGsI0+kOQO3
hUienGSiJUUb2XujjYb5suOtaoYSsqVw/ecHkIxIqEiosUn3qL2lO1vvyRmT1oKm
DW6xQNbH248C2jN/JdwafKyCooCpO3T+u2iiqfPzm58YMSzHF5lYpaKRafVEfFTk
C/kyoXYuJzc9miSlcQyC94skjWvxH5d6psn/Qaw//zQdTsxUScXBWLtYUcMu2zTv
r0ZD2tR1KpRmjnJpughSXUcDfZXKp3PBkBUTEGvUeWyDxT/XZU21YkPI8EteiwC3
KvufYqOh5LS7bldSswYf7+8uWJNp4Yf1wWG+DVWweOix14ltxJzOYRE+893CcI96
DLScorOJGCQ0ZA5z4roftQFoz5EojAXTZ5yx3rn97M6ho7IdufsNukjYymDDVifG
T39Kv4HOwXyyCLP9vLshr++dev75hhel+1cWUxg7dY8ycVnqLo4/eTYOmPlNHXBY
C7VnWdHpslFFpFcVMJlaIBFqrbmHnHql2x+y1HCGkVWtMBM9eyQguTiLKDHxbsUg
4iIWrp8BD6uwCWfM/7w5IUcibvuwa9aoeibmts3vygTSLR8RIZwnaW3tvMTkdjW0
ac1kvEDj9KUgWJ2V9SC5oPj469Ah2/HIKjMaoDDA42CevhaeaJDJw9QG/1y2l2SV
NWkZv1s0ydG85Ws6Y0/B3kyAL5VSEWrQmX5hXnytE0/4KMLvLO2pUCDY8v48k1+g
UBrBMb0OO9rpjE18hNv9ww4JO8HSWF0PLyCNKVKPOD0ZSRLuHIBnIoKpuCyeGG8A
Gffh0l2inb6aWlnIrUtZKVfn2y8SRcwoc2QCkC0kw7IQIQ0aN3ut8SVFUIxsJXWh
SYDaVmEh/fDr+qXclFHPuYbynSqOp8/N/x02nO0EWWMSvqEZmdy3kkjxw6/DXy/n
jF8Xg7Zb8T+dFnOCob6mOC2PaJZsXZg2jxtiiEPP/pwL7iKIViNvwAJAKt+5a6Z5
URNEso5FtW8HeO6dSLQVdFEq8jp3IuQA9Bhrim9mzNJ24zIm2l2DU70Pj88VNL6Z
5jQIgfGYkrSB52KJC1dKaurzHAQwklc4tmSfruoxeYDBoBp9p3D+WChrKRkSZ55t
GnsIdYL0KldTXrW1AF0jJ/g/71o50oxIxZeRfkyWfyKBLPbRuR+RTTlAiDp5jmsr
6uE3yadiDa+uBAT28m1PlVE58HMasAvC/pbrR7E9bsArrZbldmVa60IpoWIgs0qh
uOp/e8pZgery4Wz5pWRSJVDrSVlgPPm9fRsR0SAj5lIoSGIN8vWr4sKBzntGBG+j
jYjBU1VchhYGcgp4yipp9SikwNoHLuAwYbspguJ2YH5HkJBA9fubCR9OnBu5SzXg
8grYKGS6iRxzHWX7hgDWjfb2vbHe9gh8p85V0XZjNEQ+9mqqFuzTc0uW7tyGVVwu
a3VfK1ytrqpiVD4coMIneepXQ5WSjaMn7zvvUboq/k/5LJTSwmcwVq90nllgk40V
ipLLW55KyLczZOQ1NaBNDetgu/wbX6I2wA38hPJzxE7OEeOs26paxtvia1LvkEP8
cn1RhyNjxBYOfdBlodPzfcbVDcseFYG0AjsezThOxh8GUG3EApU+Lkj7MCCMfJ5e
Dei98mgSVT/lOumdQiBmdKU8E3K/o3wK0YhyYRt/dYN52jAPeArxtZqX9+l8t0yj
Z/op6deVcfZ3wuT6oAjGBaZG7FblQeQ8C5cLyYe9KEHSyr1tTGoMt9bVXFJdaro1
XKrI8GqxObVuN1+wvl8eko2JCZFxjVS++yJ8MRzDLq376VBC2yCIUd2vRFPnv8j7
T4X5vXH/h62GdTdxMskwtmtYm4/lUad2oD6tgbrL8rc1yxH2fzon+8PTf1ilmZTX
nl+Q0YPTHNEqmMNnrUEyeY4rk4ekANnJyJaIqUbtG3ol8q2/Fv3MLwkAzYkCxzlb
sQ5I38xa1+4TaqBI3mZKIVE5d6as9A7OoqlZx0sDSuKhG2tvaWbO1HURGV53MP+K
XDy12JxJmAvQ9Q7jz7bRI7RtTAXRqIYMpMXal754D6n42b1fGl6kN5E+mOp1MZ7s
tmfeUQdhJk0kLFaTOZKLdcLXzToHlZMhUVQaA4wfj05lzBLiwgS9PY3YsqpSb3ST
yYCQ6ZIgXypUO07WdmZTIN5eMkria8LvKywUW4Nqvt6/umv8DwkSKuKc4R2zW1U0
uFYzWkHLTZchmRgzdj1ymaWH2JZQxCr6UyXK/TyCbjdLD0h2AEaoaOh/b98a5RE7
DZpyMHAFLiRcHFBssYd9JtkXn96QCOP+Kxp1z1ilaOBoR+POoUhphdCoux0BwnOc
zhaCZGBUKPbhhWZVZ7iu1Gnipf1GPWjzCVSr0Bu6jSLHO/mIxOcYPcYOlkv/nMNq
MBbXuoK0UOqwlnd6IAUmNMd2F8NbjtAtJTEL9+zwRbIYZLgQtDHfoC8bW3p/AtIN
r6xkx5XaGeEYFAIgP0iuvvs3vYQAGmFYHlD3gXH98WT74Yg2B3Zv/3FZ9W1I+X5f
KOSQ+dmYaTSQTJ1zOdKVyNmLP3wMJvrlZGssoxq7VRJ8wvy3j15VOaWrJ4szfpPF
038qkbiYSeTIjoA2pLAO08SPAQrAfMmkOay9eVHEL23S+qDzy5HESMhTnhqhfttb
J0remRs56N7NHhUQWG6jwWXSDbyJJdh5CpRIaZCZ1OKVKVEKM+RcNvjC1MY8rj+e
Akm2bjgNzCTiUshcpJuMTUAThkkciwlmrol+ybEOh6m3MFh7e9TIOn+agvMgO3U8
KjWnXwmZZbrkD3Sp9sKR+FJI6YqXV9WItGBd4aJTaXI1zrwd7aKAa1Lp6xpHAsSG
fHKCDF8Y1OrZEHdizkLC8abeGqFaRVL0SQM6oXoWpmy2TGY0FQjgwj9t72CuPB8O
I+vbqcM5QdFptudEz0Pk7KC7mHlWxTNpaA6tGEVVwvPwZFXP4wF29F0bkfLETDeL
BO258si9VqeQWcoF0SM9QE9V9lRWCni/pFf0TIGx6LQ/Y7f6pLsu0cNfME2oOkjs
tUmcISBuAzkF1niosEZEnT8gIwMsxIGavXnNqdR97snM3kiYKOSl86n4wRDyfmNV
tA1CfTJLgJ3EyaCgrGVbSY6/f48m4H2NGgwFbQ3eQbMoaN6Jttt6Ozte+lAa5/x9
7IXboU64MTBZr3eqA8iBu6erUBm7iUeIpldN6gN7bR2jo1dYFlxSC/YNClZ/HEuP
2w9nz7sMmVZrR4qY7/PZbFM9puXrXPeyxl/0flrGR6b3c5uW1lGfpqKGdq972pbH
tnOTAkYLDdZ238gsK5qtVyks/2UyuEgExNccXIbbPAKupgpUDU3V/ToChTn3fbwb
DNCnYKxoxDfjBpzIBZBDBIME7uGWoAgVgnx+XLo+HY8BTIMuGaDky75iwu1VbYYA
DSboWnx+IOgoETpQ64I8cjQicYK/Pzn4aIyDHQLbt36fnMjVBmr0eDAXHLwRhJVi
a5OscypNg4fticHWLMvFT4pWVRrJnrFrL0iZHzJ88I4nWul9g31fU/Vk+ZIRQxNk
0IUN4UDWrSKg8hLzEURWNgYDXZuJWdiI5d2ehIfvQru/JIn6KJAVCfqRHm56LgIW
xOaabnTOlh4ptlT8CqrAFf54W5l6aVyhX6gV4E5U5pYaNfTOogj9NkphivqR+E9k
TT0BbHMsC366HCOS7Bh+gzdIddUZecb7KwC0O8iBlJHR8aEM/7eZhurZOrzSPVkw
HqxQWadzl5ZDHsWTMYCs/mahl5erqy/76QFVphHFtCKznnXzOVb5WeJaimW5gYNw
o+Hm1aomn9rJE3MTWYxFKGC0Oqjx2huJ2b14C1FMd8fuwReZreVVzqiIjVv02Z31
/Y9PvWONSuZbxrWa/iSWXLRCuyZSWf/lfkFc58dUwAxOwF3ohSbnTm3nzDW2Mb1Y
rWZ/18SEIMG7/6LYnrc7KhYtUYymIMrMorBv5gmM+M0s3BgbFC+q5mbj6T0qSerG
QqZzz95+pMavSoVqkEhfLnSYswCtCwPHpdb5SKln4F2cKNIWM4Wu0eGBT01faj7R
9/u/WOj+UxVc+5zIC6Xi0Z4lvA76FqqdYkR4Tty+AitOyqe4A6ZJmrWf9O18iZ/m
YlGiOxaZblLmIV1d9zPEFqhH5UW4QMKcY5bN4zbMb/JNxLP2kfaXHrHAjIvOn6oj
wZiljVfPGo02kKGmmLofCD0wJcC4g4lRY6mRvNXFS34I4gLkTucNImu/DPBoQJkk
/FRKfj6G2aQtoqmKQlFdyRxK/fJhocASE1Wi79n9kc7zc8i9NUGBiN3PE5eSUTSh
MY8qDnRCOI56Qp8A+PSoH/qJ9GizlrJe4y4NPeSGR/g4kbTHF6fmk3MgD5seBuxz
IsOQuOCOknjxvXfrbaAzXuxc/tLSkpUrYkor9XU6f2AIZKO//DdIAQ4xGt5G0uOS
+53zofvxjphcnaAis+FJFA1nCxWodYma9OQQAb3OA3+c47qaXe4m0P3v33DwAnsB
tDfhetYXhuWkJAFn4qNOXiXkuzqUxskAVdUvdUudSOEUp8RBi6ry2iVGr6XaVCgq
ygwOsw5eZY6tBwh/9NEqd/fWZLx/dRr1AlcbsDWOkCf3obsazyx7ANp942XOdEGW
zudh8Q5B+j46m1X1hRXQICh74I7/RzaCiTc+fKJyuMhMPu0Q/3Pg+RFB6WvmMF8k
ZP+WacUIAiHlt/1H2C5REYPlmoBGz7SVXvk2msfW9DjjARzPLvDIiwcqBrFKj4ht
7IZFrkCowY7m8ldDklxn8a1eFD7A4R9/GzlSWH52rWcyjW+a/FdrAGrpVHniEoXB
qO8T+PusF1nP921KvvDzzSMDPxg3bBzmlklN39QkCOjd/n5pUnz+iUmZlcMb4zYY
iP48eGtUbkTGnoczNkLPfRCzdvMAHSYX3YFPhrWObceO7pKWCs3fDMtilpsbd3WI
rE3YNHR4wdCK6Ig4ijFgr0VdzIeOFUV4Q2eCo+vDQNzK5T3uO3zEhfCU3uhrdG1C
i2VeXaNZT+JAAPyotcabD4sxaL/f6V2oiPbWfjICtEph6M3Fg1gsmYX6ljx1ZnuI
t2azlCU6ObCkrKJyzJsNYFu+UXMOryCSPU4LWCHo2ytnulVDdCmxOW2vcv9M0n00
1HM7J7veKdelP5LIKOThIOfKw8pYgNsb6fy6ZegcQ6vlONNkgjfVOXfV8RBzxsx4
vtvZbiWV9AgHTamKHmFPRCsTx2j1xwLdxEzOyZGIsxnD9SNzjC9FhUhjNUpXHgYq
93284gNf+65tBGfa4ejmU7+zKlaEIHTn3Td2+0DC07KKET1nHOi24CyP8uoT0G/l
AJy/Pou5AebWNh77iCkNQ1Gym8Nz5ivFWdmRZEs7noKl6V+DuGCvsDcDIQdFS+49
Lr/WnzhrUv8Rj3V7KOD6n6sh8iFfYHjg3lxj5JQ2qnopDqNu9+gX9+P5kMrOYRhY
gp3TnpSBu4uGKeNcpPOpLgcPEgQcrL/D+mr5tkdFYuurjwVvjRaw3DInCFTXMBTp
7rTAIIJvQGS+7SmElNBdNwCb3hNwnyGixO4gKcGomlkXAIHH1k/rsdP4lQO3xDZm
7c+lQm3lfhevwQdj/P6YXK7peuNr4zGK/jazqbGg7WTPhHXIhil9Z7P3/VtsTV8z
PEzgwl8Gt4tzPkqReVSiqYgRYKQxmTLeLmXNJIvjZibhOBVF0Mn/a3HrZVXDrz7o
n08sl/gb3aIw6iGWHyNBIUhN/sWDGkYITBc+cG6VAOKr0BkFpmG/xkrcsj3R4qVQ
x+b7KN3Z1lhDFvq8QaJno/9lLRc8ZjkBg4SbJ4FVCWj44DahP7N1O3oybBKrtHFk
FANZCxeXefe/qs/krkzLqvYFgOiOgqrN245/Z9tbhodu+6V02mqLzd/idgijnDrv
mnB3ctOh1+F0mwL5Nix0ZIhk7AeFhJgTdxpm1PQRxOJUpxXbxmBMG0yFYPgLuqPm
QLLXo0Ma0iO6sou63rZJ5H+5VcGP4ySdo3vYx+8G50UP4ulpe9WnY6vTiMBveure
etYUQg7gb1LSMMT++8XqJONG6BmhW5Uo2hAFcMK4FZDBXQkxsifLOD5d6HjVvYZk
SxcNk/ce98Tlc/0GCcaW/6nBFxc5OmUCZdRceZDj3mkcI+UpMQhxlC0kF+1dsPT0
oYy6jl0g3Jy0oHYtScdsiCxiTImNxU4ossrzI3Id3vHmr/8EkxKLaBaMuIB+EZRe
QWRx2QP9r+uIvi7keOumrQPQEyjaowMpwvzJq3dQvpMbCi+mIlEeHsA1JOBdB9QI
2EOBKWnZIM+faQA+ymojZbi/87us5aQZ5HUgMFl50DeLxQ8lcA3NIZuqFJZL4fS2
Is5a4xUC2Qqwt1pu4tnVe4Nz2WTbgQdrcOuugKG6qmAmf1UUcYstLLHpHTv0vMrK
N4OnqTyK1ZGmOVpeX+dh4YX/DEs/G300BG+TwPNSeMd0/zdp9mXWPrsQ9D0uGpHO
Yx95ai237L798EH15AmXFj2fwdZN24aeylFPb4syyg9IIt++0QCg6ljIRYw0bKMh
CsILFEf1vqg/i+VXV8aLKZjO61Ek71UbaaTRppT0jlMEFSdbK6gKrzPX3uwEny/S
ziDhGyx/jeIjdQsSKOw5GOgzrLKuuA5w0aGrg8guTEk4fPuI6FmBlvsTRHO3ONUa
NZay2POZiKgHr1KwSohtUC8vGWL8C8gHp2FJtaQGeMDO9QpxxBynz/KwghziCfUM
AzBJbdITUHVS2wcqtGKvYgBzq48VhysefmD7K44MIyShah2IN+Y8jyZbRV7aqYzM
tNmrDcqOmV4vwYL7WsyQf/yTtATmNnUNmKR6dmIoWJslvuuIiDWAV+PWZNjp6taY
34DS9jKJzvLup5QwAXrKHrpYXvr4pY7xO1e9FcnjmdbMX5p2Sw+iJ0cuae1Q360H
2y5D52oBJkrgLykS/eMlSVJjdTiXhd1BOHsb3FAj+JiHhpFOweTY0npjilAGYOzp
xWvXWHCGYNJ4YQSbIFhXhN/uMKuICjSt7/sAHA3lEMjpOwYc6or2p/cInpWdhy4l
kvK4GrLG8CYhr79iT1uxv5LQUP5bjx0IJKA9AI8k/1vcP8heJR/EzzI7ZRmpz0yS
SoTbpLUPveMyoysgFsr1/AbZXPxuo36p6TCIFi5iSOT4GD4kZMa4yQdK9/KF2lNQ
tGQh9Uwg2RgOjKfoOBy2J66ofo6uptzB+3xNGlzSaqHd0fVZ7HyNc5hpHkXuk89g
S7snd64tsc4Od0sf6ZyC6BmiCqu6EGBlHFSKhInVy3ICiZ+TUh9VCDwE4Dle2Ihw
9NgWpZ473YTn8je9OzIkZqGvrnTJoX45TKEgWJC316hcD3xiRQNId+VtfHqM3wkb
3I+f0HKL7LiBCpNV7WEgzu/8fBDReqOg/4oxB51EaoNoXi43ssAh97BHqi+F2bip
GpW1uhLO9lWlWYbvjTKllH8NHB0g9Ocm6aQGZ+U11BIDjwuXWytMp8utop2KVi4m
48OavqctlZoBUdb1240RfVPV0kcV/8/TLmy14dj2ytlrGgQWeQ9/9Mu/gvZnvKe+
lhVV6P89NRpKjJSTkq/bvrgAasL4fwycs5Rn7ckJk7hjlyICK9PP/S4N9NIn3ikz
/hmW+BzQD/GUYp5iTr5CF8UQsjaYHwIBcY+tSW3aoU+IyxHi/rIQIyMCC7Y7MZ0Q
3mmpwdg55ItP3g0d4lMv0/RpqivNH3sXGYEHtR5oTyfu9XmRGViT2+ze9V62RJe0
s5H6UNsaK9zhvirz/4Z02pJVfY45KE+r1RFh5JX+lS5DnzzCmQfT/heVUcwsVwO8
NTV2SHnkDodlUlslQW3uEGbcB/lQFZc8uwG4ewq6i1YNG4jHJrIFk83ZTPvqWDK6
I2NmPqKFqGGfSXXj1yUi2XQWm2XVUdR2wFt4YvIguLdx2VMy26o1EoxSERD/jG0r
Wj+h/pe5jLcExmI7tG0w1f39bBlNx2jU3pSXOkpwUgBtlsMDiQrEec73epUfM5K6
dyXdJT95gpZhFXB/i83apzDJHIpr/xuFo+rzpfLDW8olvcQkdHqLeu33muMYqZxH
qQsQ51vNbNfrThfvIrg217qHI8HQD5SMm4o3/XmLZ6PrRh8nCJohNfCTnCNFzBlv
id6vIB7PflL+VHz0fdGffauoHhciHCVxRCYD+izfjMXNKG4GWgvcv8X5TZkISe+O
Ek4VB2eQlxmkY8vnnj8vckk40/jUtbpPq/2o5oVAtVHce20TtBikVVtKV4O5NN2h
aLjt25AZC+Iu1NkNI2Byk0iFNfQ9pNCoKgd7RTT5SCaoEw5hvs4DBCucF7MbaRfk
NXaBzcT5WH+/Y5fR0oS3JBnkmGNxVtlz45J6SCl89wrJU02gWeFZZHN3caOb0Cl6
003bKEjyJE+SHcKTsVHcbtUIMcnPNVTyA831DYGpYvZPjTsnYg4e4Bzd3GLfNcd5
qTXuKz8Iet4UysnAcmfclyKc8ep9wsjkXfr9+6hL2wGH6q4cY5WRsMi2HROY59ai
WySNIAVMOpvZ1K8cNVq+uyq1rT0F5Phtl5MkvibClLmw7MB8cjjHl9JHb2/cJTb/
XVl7V9TIoWU7xePdZs/nu7w7ZsxQvzIuy1uGwE+lLFNofcDutNMiNrOV7zucyAOa
Y82sx139Mg1kRpAsPeSOKHLgqP79mRmGl2BsOZ0MmySzNmt4ZPybmrEo6GzGWI/K
FlPFc6DnUefEpYoWSHsZb9f5IwE0UF58ggw8VrTvArJSmsiP6FYzz1k0pXCi2/8F
2xgn0JGVDAV1rj1knWHD/dv0WqceB/IXRLntBPLIWLhzixh6QFUx1OuWZabGJXWq
l+lmcAHz0mNF2sFB1gowyaAb+h9oZuxb6/31DFbWJmWua6pHdbhTW7KGjmaZValE
qlfEd7fmdwFXON/90fnIZHDe4FSXmGS+lATgSCvhwC07d4Bn92iEo08WTjXKYk4L
47nez5rXhrm62ve7UDnnNIcwAeeh9S52dw0QBX5+Du9GXxZgXyqPADACMQ3NDwGJ
9mRlPtyFBpwy/JCU83bi2bpOuh6B+BeeIIdGba+41tYkmAYdrHnwmJuN0rm5Xh2+
5klb8G6VHjqo/clfXFDw+r67sQ3WtBFLZ9DqwTXDvB83tAMW1L6CC6NQo9QmkiVJ
/hOSq8a9G1Umx8RcE7AikfN3HTAJ/bVtzsB3Us/ZyTJJ28ZyiKFHemQZKGe/9Qv/
rPreOy/UVdjEwKlIM+c14GBjcVDfBdE3E4tVe7VP7aBkW54Ad6nzbxvhipKn9ptF
5UNOhU9j2qsMQom+errP3xexk3DwYLoIA/uunu3pE1kvgFSGTiMuWjMVb/VSTaYh
8yjpFMM0LHKn/9xMM+2n+r5xwSTCE3+fIsZVI/db+j8kx59SB3dSUfYuv8TbstuS
xf8dfIEJ5dUqB0P19cH5lBXhqDv0khIezgQD8Kaj43UWyPEeLsMpuKx74TAqwSey
oeCd55EG/IaMNkE1fwVQ9GZ2YS5gpmf3qPeLU8OheYthSulJ3PNNFqmS4InLGM2R
rl4O9JCglJCyP0jyd4gi4uj4N6YfNNeR057yTCTvXAABODIr3lwtlVyWmhiVbpyd
tlBSzifPCqa5nQ0db5vl/PuH8Gzc0wpR+ZffFhUh3fpj9hrYxkA/HHw5Dg5y0AFj
GiOmahCxsxaZcB9prsPh3cYdt4dvvPgJYjZ/jtKdPJofBdtxoGCdOcbJobPo6izg
wCCsun7psdYLcIoTzM7WyDdHPyxVFr5hzCY40KMJehOs7fxnZRcrMbEaYo5h/uic
9H6tWsn54VvzhiCf2Ilr1AuDEe/wxveyFE3mJcdiXv5C329GSxlASIsd0Wxl/M3B
GWnQ0+gxl91yMHo7xJjXrtiDQ4HX8seLpqdEhZJNujqudO9P+rS9b93v5P5Eszyn
0URRlca7nGi3VdXToo03dF1dgHv/iJaZ0IG/Wb+0hzjejrzgcG+6gC52G7CE3Or5
tUdeh57tQpY+4CcibfyTry8Sp95ayeN6cA3PfK2IZa1ks1FVtV/D5yxAXf9d7SiF
aNPV1B6MLlFmUvB75kr0gR3nw2/JBlKsdnzVB/NnM3d/gADyO+E8iN32oMigef18
6C45xJ40r9WzrNRmaznim5/MLkUuJ5B41aYQyEcHuqIW+z2rT5UnDLBSs8Mjthma
cBlU+198233egs3mtuFAJi3J/zX/rqdcisq4az5ImxC+5NYISM9DHhhkhILEakIZ
zT9YRYgQ5qilM58RDvU8r+1aw4oFHrEYrSw66vV5qVmqfYcSUVh/3yfdRJYoQZD4
PjG8Y8mJwWgUWgeSTvsRTAWdzfwiet8A+0jTHgA6TjMwCwlAW8+6QHKvb99r+xok
6W4uLUI/NY17huJv4CBqjRNGN84LuA02ELH2uVqUNAM0ptF8798jxO8xf5DXpjVT
ulrKB8W7fmamADAgmp9Ze2Lxj10RBRo4zEijgZemuYf6+vYsLVPxvemfMvW/07hw
h/d6rl+mYaI0nn605VnUQD9vqgOabqmTg0ihJgYc/fmHQFuR1zn+a/cN02y8HUHT
RDOUNkOwED79Mk+VC4F+OlzfsUmgekz3jvYVgVtNaZg9bZBWfXfRGY96aaw8g4PM
XETSXI92nbcH/Ya4+N+om6oDqxQ6gHDbypss1Qy9dWwhnsT/qVBiulScz5e15qDQ
nDzGWZEQRwP3XIYkuNVROHClXVvjKGBr3P7BG49ycjJpOMrpd5+3E4K6OMu/RL/g
UxQuNjuMSBa2j/vv2LQ7xO1jK6WtYev8SASIpNBMyD3fE+NG/uGhy79MLF7KJfbL
XZH1bzKwGu9+pWE+TMFhUFpV+Z+4/wr3Z/baEgo1cncRkmtmsjSiyd4FPbkCqgTH
2lPzpZuhPyqPomQAcG7APwXbYXmV564hEnXT2bAjQD5d+lQ9R7p5yooay5Z7qroL
k+3y/gLwoJ6uhtBPHRdDovaGNWosuhwD6EigvVFyJwBAULcakRPEFyl9oCea9+bp
LFp1pgXiFJJ5JU/V1ZP9Hf7kC6VCTCy4QCvyWI3Nm75QC3hURKkNWvk+3A9c1psz
dhDsElOdY0Nwp8wMzhyeP1GYhLqUovlH2wofR2zrZh6lpMmS2SQrPZn/4UtNpwFB
TXhYK9JS46/h25mHMhb8Y2C56/bpvwdgtyO1kB0rvRlSUGOCHbsvC4AAWNx0z/Oq
jCaC5WjYolD4BR4HawjracMO3MnF31iOvHxg/DtEFCVlVKmueXWwjhI47TF9V9Re
c2OqVtYXdmutjVsYL4+P30rImCMoRE1HeDp4LpgGSrdvZrCXFZXPlSk39IqqW1Zx
h4wLZaQhwYTqCPd76759aztpPpo3yizgcJMWRhQSlcuOA5yTG3Q4HdiNtlY429EB
fkhXs4pkXAr9wpRLw8Xs7JyXmGWIpq2PtCmG23p38KckpqJABrS14gKGXba8ILEn
Lry93n8qTbOweuagYNALGZMC0kN7+apjfz6BybHuRcGbK0Uf9OwdZaUYk2xxhlaG
oLD9EIh7dSGNtQjJC8aPoEK0SVfhCTwNcDnjCL3mxp02ou17cbizjl4KWEjQvPu+
hHG15L9tLg2dEdxRtoc6wCs8AvthGY7t2I4ih7cSfMAco8nsgKgqZTWAyCt90rm/
UaV+O7PcZnDFIJqUu3MaBA7XQQPX+6CCsztKCs1dt1OyAVx5t6VylRINVjQOxdYO
slxCkRu+R9W+93wZPMEd2kVVbmXm29K9qDcItsbNKpNAcY0u4pUWcGCqEIX4VzZV
fY7+J7E1UgVcM1ELW+edgHq41il3Tlfna8nGSzOz7qJbB9gBD5N7AF6dsjlgOvnw
yN9l9JH1lTBKqxLg1l8VHhObpcEsjwYSziiuR04lId/f/DBEFrEY/Wr9b5Cj5ID8
KA62SJQnbvwiZD/ncq9sux5F4DebaY1S2IP+YD6lcYZO+7wlf4+rF6UP9IxGUdXf
0eR9vpTslwAl8458JvTqnN84cCQNJ3/ghk4cPpoqNbN07SHd9cF0UKFNUqiBhT+K
jsowZf5BfmVR6alHxKUFmIgMb62p80Lz8F395soTaHZDxMHmyA+hgk0V+vAmKjCG
Skk9+DSkhvN0vh6r66KMyPRtw3wF9Ht0F6n8y/Ythf/5xKTjY2WLbA6egZMISsd0
Q+lWSQeU+vcAvHS52yuqyaPHJODCyBmqFKSOluZ583bwjpKljZ6vx2M3ZtHiunIL
KZdRfHDfRJZDKQ7syO0j+Gz8b69Xc5RS3V9UgP6aDLddhUuvjZ6biP91l4zO/Fwi
5Iivipev/gNu5Z+b48X6wAPnfZTfVqQBYKVhIwqsteY3AbqVTyXZqCMCNRgf/mmw
seTi2KZhjeLZlpRWIVhhLgHO4xYr2hip3HRc+zxcBD+YrrtDPRfRSPgX7KGHeGbf
H58b3tSLulCEi8NVZGsy7nE2eLKdfe64YuLS0iKBua3sOoJKvEK9Pf7IotAubOmm
hXkCoITW09dJTlaDe7xdtSwDbV4ZTGLatqmLGPjzXhpXMxqoL5OKnOZ8iUczShKO
x+EjPAJ6CfZfOSNgRfvhqBdy2f0X8Wxp7PkI0RkYflSxrLwXVCCRimOj3YgXdHvo
Lhi6slr6Mky1D2YgDYVvXFRKqok1uqxT5A8cdF698G1KzPTSVnXYv3wEEfwNWkIr
4KEaOdoE3HexxxmuZQXyyKUlJPORxu+VO18M5wbRkKy4ZnvjAvnOvSEUFsoCSI9/
bQ/SF9dMBbeoZJN0brASQd4Zw5Y4L1SzKWIauHyPfSNcZAIurCNGAv9cVOpS/yDc
h5086bR9Y0Bp8hlkuE4388Y7cQpLGYLvPnPsjS6fwXELBKnleW7vdeYYpFLOlg+S
3ThVhNwprQ8/ooJUbb23hiwlC7YUy+XJu95gf2zvmkJXvGGabqAz7fyqHRzbbK8d
sjgMvY4FwPuZuRP0gi97mOa6cdldH0muLALOUSjMp4UvLlU47DDD6e98O3wxAiqA
cwHGvf6c44YfSmGfKgWAmbQh4Frqb/uTcLZGmZ4gKtpgQesHtkxM3frAvJQiFmlo
XQDCx9nQ6Fr8kewOZO82/75utUKWw4yJNrYhOJIyns7wbKQPavuGl8IQkUYByQ46
bmdM9f0QWl8DqQ7E9HxckPULIKS2aAPxS+kQurP8Ik+/NgBP5TuNeGuSDznvgDxu
568ij2S7DUBv6B0swT7+qjmzoPltYpJt0iAOd4KtokM6uAxpO9wYTg8d8xqKkmAp
spYs5NQNu7/jdo5QGFXI+s7EYF/Q0jVaBjuOp6PaKh9+WKEW4BjkYmst6HWvtDsk
yjhosXZesGjiQj3lzJZESbScCe2DW/6vNK2rgqTAfZPDb8GDVwWNhFd3DoPy0jrA
rbSsttIQYD+3VPpi6mtP9psyntGJQiwZSLgaQAOYSredGtreYZ9n7MU0hPUrgsB0
8uzWWTqD9VMEFKboFPJDAJBjFLpcU8JmRts7UXO3Ge8ApBgmKMUFM1ViafQmxQxJ
OQzu5N3xVTjEMWa+xwicRw1/0V/SEbUk+NYt8j7/77yb1jVct4PmbMzhzPRJBtS+
jgfHnJdqRMnl2byGpLfm7UkGiyHdVcVlPcJM3eMMiBvW+FbLy8kmfSR5U1xZNqeH
TaTmn1CXM9TzbMiZuGbEJqlrkTfFq8Xb1ESv0QETWMg48gE6sRZhSdBMGzFZd04t
ktPTlCPdHnfwtc/8KmxJ6w8z6JAhSv9GWPokRpCRyioAzUOm48BtWCEfYeFTQpL8
f4gBzR7QaTeihysRnvdrIEWaazX3bN1zXx0vkjRaLmJ72ouKPIxlVaBQ/iymIw6c
dMa9WdzMMni9EKItw7lGmzoXlG6d/BIVK5KEF/Tq3Jyv1Fwegu5BUERDQhW28fcH
vOW56+7ZVnuDY7Q3W0Hy6b77djmkmGR/RiAOdQJAU0teQ/J3r9zZOh7Yw9NBimi6
7LgxlZx8E0USaforJKNBkf1s/X8BcDyAvw8wtW/kvIEDNJqSmle4Vlx+9DF3x0BW
WsONrGjpFIw0anVyytzrgcEB/Xh8uwFwTOvUqIrtShobC75Gt/EOPdwNXpFUdJ55
vsMVl0s7YsTZg+fCmkC10AzBVM9v5VZntFzaOQxjkPlT7al3ibxgDrLpmyUXpnf6
2+f6XbNHrtwuOIkcdbpwjpLikfPirnh87T8mz4pZFb6ROZi/kI3HV+aV64USiWcK
cGS+MIuH1QfVesYmtidXAQXF/9SXflB/9F7/GnwWNwOlrC0WjjK/5lTZyKWeiAu6
lKnLyLkVcdIgLl9IcTrZxrNBFH6BF5JoXgRvpfl/eJ8i8+/x6IW0Fhnw4P+RXRc9
dsZcjThWfiCzZfEnGVEVd31+WjWuS0Z5NvMwOObQS3jjVgH3XBkgjs+xlo2Aea40
OnjX+Q/kuxzaK0cyzspB263MOXdAr0fbzvCZawCRGBuQl+eyFjikvCSGgsTkDjkH
anD3R3Jf6WsNj+blMGqMtg5XEwHs54cV39y0A1BMNJ21tqg3CB9OQ16sYTo6+X04
dxQdUlxE8snr+TZ0xfCh9ntYxMYukI0XDnjruGiZ5uevV9c2HM4jktVtKPS94C1a
3EsIFC8dul14trcP44Zs9zKUhUhu44Cvjiw2FOe8pGAuCPXp+VXosLBhlX/wGRev
8uriwwZw6RFf/LXczxkeZcD+3/Sc4PKQw/55fWaKmNVYGJx6QuzxMLfvAcC5iXsN
JEuCDZEJkD+5re3Yu91HLq0ONcYCOa8G7ld2s9++qALYM+byva9jVrOn2/5TflB6
PplITIqQVKI1qKmvLdFUymJdokjqnqeHZvyGaIW58BFAb1IPSJeO91rLcJZuZnpM
izH6+GBOitHkVAuT5zTbHuH3MTQbIdh8bAFwMSsSbrbquk1r0DSZvwloE+aziHCY
B0WEIwduqPngHRxmH0oQSQfmpfp+7cyBbLZILu7XxIggrXAbSMNNFhuwJOn8O7Xv
NXLblBCrCk6Q+UkEPwu+Ufi/EXJic69n4aaXY100DAoewdzxSmPwQjg29/vpuXW7
h0JEuykDftrfcCAnNw3zn/4Yuj+E64e92TSEYP904Y/idso5S9DiBKFlEGb6Cc2g
3COyfclVhc86C5lmueUNg6MuWQE9senDdaUCE9c4ijtH/FjIRAROdZNRgh00NOQI
gIRKMjFICZxNaVk5TtDqqUuQrfmYEYb3hPMMOBpWbNdkoohmwsLt6CZ9FBZg9EOM
LaA7Fy3Z8DqeAmwuOLi3C+v4PKq2kttpe5quCL9nYudFrOs+XOl7RCjU3am120y6
RG8vxeVKDR+EkKRg9FU8sUFEE0PDhX6BPbgt1bpWHMIvmv8wnmcquIBRB+heVIIV
MGPOS0QzaaMeucWThRXIe1a64sWr02ohWSbwN0RabPNBSarLuHruIdh4Ms/7bE0v
HIDPrZkx1w6FGgA2pxwxfjrPAnnhT+u1l0t4OlguoGwTlNC7tCXpcU3lf/DM3vAr
oLDaTYawzt1i/BOixu+p0fZBKPXERP+EqSvRcDFRG9Kld1JXc6oBqw2XJ8grwRVV
6soNoJcy34Zpv3f5Di77NQCrRiKHZ0bYvoaXcLS098KqfKAzX+5GwYw+YbziJ14S
3byGM/pOs9EqNpGqgVGQGoNlcf5AxUrKFB/TFjwhydSTJL+Sjc8IP/53DzN8Lz7u
ERJ+AnnyEWQC9OpRtNInUuLbRAAz6DlrGBcp8pcXOR7oF7EpqV9GIeCewmKTl7Ea
3aWwdEJjCsWscogallng3joKqmNkNa/qQEEbsBGzcSfIxWAnTzuskYeBZvPukUxk
MXYsd4Gc2n/PM315/NAHSRvFCh2Hlz9kNJ5AwCh3VQty1kSeJ53AbEGLfANMslnG
SgOuhmbJkKzn97Ws3JZjo4tDORePWzc6RI4lGA3+vaGmoIPIKhr6Q/t+ER5b8E7x
RB+LfK1AmuuqcG36ocU9xOeW0/hRLDvfSU3Ly6SgBeEdS4uP1LbhJLEUAo7oJp+j
FTrD6QQIpgVk7oINFcwzXQQjUCAZsqSmLXToHO7oSJu1q+W4RNe66W7wmdZcdNcY
19beRd1KnNLxmd8urdcWwd3vPAklmlLQm4OhLFrthZZr5u3Ql93YHXOusCalLNWP
L/UouBvFXtDL3nZrE1d26BJsagZ2Xp9yPVWL2Z5+rmB7dRB1lVjSxrtfUvUgu6gQ
5MM7mtdniqbS7N8ou2J2mO5VF9fyznVx3mdF2Yvy4pMCmM66+XAF9paZACgkBeBU
10hGE3QUMeeICDxPTE/Sef8Zlqupt/2PEbrMWL8F75aZywwat+VGrcb92/gUqger
iL4mqaqGA3Q64AHEXdDi2XUirGB6f3V9a8vRNhsY8Q9egP/VBUC5tMbsAVW8wfmr
U47rUIHz6n19gL7ysDk1RkxnKn/sWioZNavFId0T9Hg0Z1e2514ZP2Vk18B3DfFE
J8ZBMrGJzYN2UlPHMYjKs6eJmonxqEOL6433S8Zobo0O0ARYjvT0Kqn6pnv3W1+2
Gb6dDs9fSVhx+2wEymuGgGdJAd0Vtlc7MZmTKdYyfg1Xv45kN5ydXxJywjEA8KXU
YpneunxsZz9+1x+EUxbkScirJwwFejQyEs3Rskiky5t4+Tq5T1PUMeI+wj4iGjoo
DmURqlFx4iTPtnHvg4JGKj35628DfRb4PbSg+lqF4F4PUsVSUbRadpu0hVAQNEOD
JR7xBaaWYbh03u/xPrabnV90i5IQXTqqCvPsRqTaEYOGpi2wmyi9Fs8I9Ke95WWD
x5lWudz0cVkent9ksqQLP9qFW/mlCD8nDUScVpdM3aStVWMs4xJXrtNyKxjCbLxf
eJE+t9+5F20WBYjwdakKsy6cx1vuF6HTag0661V85O1epE5qyFwP7S4wipc3yYVo
v+klETxG+awfuEuIJKybe8J+dHdpPwVkDDefglBHwB5dIAcsV9M7g4+1soCZcviA
mkaKufZFJc7MJSvc7d8BE8WksQUmD0c6c82r+GxF9sNpxlVOyePUd1UtTtd7ylMG
mGkM8BKpJHrU6NPWXTgo1uMfugNmsjGW4n24nEhmBnGT9dq6Vva0lqXvv1MxYXkq
9EZ4lBludaKTFn8GGJv8pDJDKMfghMaAUpyN1YSyXmbJHPoVRSxoEtvbJJLkAGe2
gCOhtNGYYWaJKwvCFkX4qRXi2WuLjhsK0WVPjTg1QR3THWGKbBA5XoxNYAkhktyR
UX5yfR2yGi1oq6LUSD1tWT+PqZ1BChUc7g2UHYWnTiWPnDMnea7umEDUTirywE6J
6xnsCXlao8iXL4sOs+88qQnQVLo1ggtnFRvaHsaCgFOQ1/vUNMwSjzo0NTqU+8RO
YC65WxGXs5fOOOmCG2hWQLlqIL3vfU0CMVWIVbl+DzWOJ0smSoB23KhxiR7vxCO5
PwkHAduIb0D2YqVoRjZsM9846eYjmQh8KON1sxO9HAZwroCCrzGWmLEnwRXURmjS
EqOhxB1q41ZbdZCe3EFwwmnfSjaWiqjGjdarW89uarOijnlW3kYUMWzALcmVfgGY
kd2FdRKxfmxISVkig5XjtxxE1hpYK8kfzS+Vz88/4KG/EzvqrSwjcFKr4CrwVdKR
3XOfKw3RdRu2w32OuJ/7QuiEvIUygVINoReFZIIbeD9FPNpRxdPrYRsm9MEwAMO9
snP9RtcpGNhkgoUOV5hNKxaduT2tXjtjIJ6TRBdJgU0b+hPLlQWxQ7T7QE3Ks9uR
pK8X/geoXfPRkWtqIMibGAQr7McC65tnjA7ZWiHMN/xK4Wi8oqJbeG230z/DSXI6
dxN6FCF4ygBryG8SngbxN8AkdZH0IJSTXcNWScZA3fSPCrwXZ2uJNjSJgPPbni1b
4jG6PapCulNyqwGBJ9LgimA64iA8nmBH9HjcNy9EkKsyr2aKiXyLRqrYgDRgkG1Q
VUUHbqrGLRaI/Al8v9LgAzqAZ9lttz5/sK0dKBfrmPvmJyw2G6Ephonwtwo4vKnE
CS75a5I6WXQh4fYrjKonmVZwYwzkkdKonoB1mb8EeIwUouCxQ+BIXFkX13+uJbJb
uclI4pqUtIrXn22AIihnf9CPNORvJRBWHJmq9gKsX+2s9jAfbmXENfgS26RZ/dRO
t1zeizWVS7r8rd2Hot9cCvgWpMZ84zgK7L0XptOL6wM+zDCUdC8alYdJiFufp5OW
ZdXZeyduXHrDmjD6WCuF3ce29WJuqcCs94/tHuDyYkm8DPUYQn5yCPe39Eh2hgrs
sJE84K/w4PyzxBmjIWtmL6xWVVF4RnB4mrJMhxgIlE2AG/KkJP1DhGRK1C21u6r7
HqgfJaR3zITufxVNYWZLsCgzvS0Q8D2XeImbdByQYAZCmdKQsSo4s+hai0//ikyr
JI+dfNuqzVKTuCC5Pb4uRIWzLYTtyTlwD7M72a81S0esAbfEP9xrr+96+GsYF6jR
i8epXAgsaFvf1BiYQJy5DAeTrYl8jIEjQD8HwkeiwFPyTFBJSaBswaB/nOPSu3Qr
tqjbrQZENCiqU4rVwvVqvS9liSaU1LyYSgSc5aQOLAEmUqNC6uV7DHDJHId/AGMi
yUoQbt4zKFRe+bH2EgV/6E6JPdMfFc9dOu3ZdTcXuhjvOnmKBEUaUBdXNnS9jsnT
5kErTElQulO7ZgQ82vFda7+VOHmGoIGwhZergH4te6t10knC22snLqv/9epwzcLP
Lwh2BF0qyYCb5U8nQG0aroeIUl3aBp7MBVn0OKltJq0/T648/fGjd2f2HL0L0mNb
l7znb4dVhm1u+xGg36o7rcjxPieY9M0Ms7lbMKwM9v7pMX/jCWxbhedFENNtJk6p
w4hhYBbTPNCZs9CFwpt9SjH36s8LzWfBRHmq0P1OarPdkDdP3EuSXrK+laTEnrzD
YZDLQtrRSQceGwoDEKTvybvw1rBMh0JSXpn6HZmRcN8DlMyjtwj9zYLXNZImvs3P
hT56q3ySOC/PFAtOo/NVPVvkmOry/PDQlj7y/NMnSW773ZyHyK0skDojznMm81pV
6H+m3YdqEJBk3UOogZF9HJLX/TRbco8B3HpXwhX9wGrkPOigdL2FX6gkzH0Euhuj
2qQ5swK7gVqchsruvsJMaq1QmhH1xJIomM9AKrUMSI4Y+gXWUbszHHz9zI3et1C3
9FhvXU0T1fj64ln+Z8vsdhUhHriPULELgt+uRHHwfQSk89rmm9l0i0YKwlOtxdkr
EhgQGthlkF7oNJeDlJPN+NthAiqNfT2m2vp5x0L8AuLBdECKQhdw0yX3wcoOo71w
k5bQyoQU/G8gLd/dDhu8/zvuAzfPG7Ep69D01koc54WtYfIZSe9Td1zqzUtrRlez
vQyE5IgE5AxoeALru0WoP9S8M9Ib9PuuvNhOZOj85/lBIS7E0uvjMGPJhMgh2hwm
CrhtG+S5bF8HTMxzpG4MJLPeEcEzegPkEp6bSayNwsEXyBHNGB0vvHNmsUgOS4zf
uFZlg5UOMEo5eJ11CcRZg8u6fMb0kEaBAtNCZA9Cibv20eM6WaESTa+qTbsToWlx
z/ohT9KiZ3Q8z/HON745nhjZYTJLJmVSMq46ISvpvmi+EM6ztqUnsuaA5OfZPgkV
L2NH9vzoJlNWFu1Hy+zcq67j08N8mbZzcYky95wd1JKMmTvtMJWn8FueHWoSO0w/
SiJMSiEVw5NOC81Qur4p1gTLK/knui6DUswohkPGa2eaDYiymxjDO+hAfnINMbe3
bOG1kfoae4QXA5wqe4kAEqr0gDuPd/aycGX2YLTNdIlKhTjnBr6J+2Tnjtbq5c8D
01AU5HwfrcFO07M/MlRSWUiF91iPp9cs2rYdETxZsjMArM6Ts7jtcolvV0CWeM9c
DOoFILxADoD6tvH1UI2cZ9D/md5pGn3hOUrRs+AXpysyBMmrrhtUBegIVnjs2y9o
VeZVP/MJtLD9aFu8KIEJwleEeKEy85wkZ9kHq+Lo6LUUjZAPfZ16v5Td3QBJvuOy
je2C2hXWgxt6uAkKG+lUnFjgEQenOKUMNxakXUaQ7e4Pnhn2/JEgV79KP5gLw98z
IeBRMiPriWwwlcrIVmOa3u7Bp9rvnPnJJ6AUFuturEsdJxRDS53kasfwUE7dgl/H
A3FCdB/dn/4fo1pWo8Ye57MfxA5wMaxXMf9yrhVCJ4+hTQu9Pa9ZAWb4oFRVFcjt
ISAFtDKW8layEeYkUBLSFP63kz7CpjCk6bzFngufab1Gy9infm79JUvlPqmcvLi5
WvQPYSjzcr0cmxKT9cVsWgKCTtcpTieWcyFRbA2b/5MDxvRhjQfdIu2mke9CLOCP
qNqvy7f+EMfjW1Fbgc7MNY7YYNkIPSFyU8qD96vYDziEdQIkSHk99HMtgdoWlJDF
eLGaoIIPkpt/RKncjNY8trDmUFyXPZ9fhqKklYiMKPObCmh0V2JDcCwsCiFMbMrs
OeWxAMmOn4IPUGxaVPE39WRxpAIdPn3daD4Iy5fDNvgNgTBgWBGctDS1XkZjNVCu
ah8LdGTTSG4gE9VWQAl+8j1f+Yf3tYCrhQYR3yMfOPMT7pp4sCIHZUugWwGKh0HF
HvtumGb8j7X4kPbTNf9gIcAy8xLBvFrpqts2WlvyplS5EMpBH10gvU64sFgIiTJ+
ckRZBCHMnZjAtimBHwNnMATUFFUZ57xevzPby1fsXA47X5tqPSFOf5uDLvUQNwgG
MDsxdunnKGcKDGMpb9eNfWNeRYix+C3YzrrDuDNxaMu8hdQtDoOyhk1gJu5dLQWR
0ZANndPYsb95lt8dVm1LLQWESRzSPmXJEFWc5WuXOeTWzkrVrQQ7x5S3KRLpLsP2
JqrwQ3aoAvFsY2mlposlB97zUxgsfKyDeLya5XnK7WANTct4XSGwMEM0qq5VMcR6
t81F0rgzZGTMXizLk9//5htHNUm5CR+UVn9ZSxFbNzgY56HefDjsghCiQbycDCl4
7yElAaiB/vIXrkrGlGpBzQR/xrRYbzbcZg/lwbS+18iS9TTQJkB3RTG7voDRhRyS
1TlkuhSpAZzIcFeAbZWYO72miMiPd+L6SwPQYE4cWS2qMpkvVDw2KeZTG6LBbrjO
9jPjRRHHB6PBqFU/2mSavPc1/4SFuTKTNbA+Tj1ZaUC7L8VP7DRhmMxqZ+XwnXXz
WXp4QWaKNOBXT2IkFdkDGD0doIms7xM0pcAOV/yAad/VajmYknp2Tw+AySnj55KY
d7762DhA6xSBcLW+VEr5sVv8cSQWENIOIZT4YQJgBDmZFFmIO+kTK8pAirT4X4sH
M7d5Z0dbAQlDOz/gjjEFjV84lHE18m9B0/mlJnAhfCfhAhgsFd0FVu+rTTOvigAC
xAp8jC4nBubXnO3aT60UDX9nrTNxkZxu/0jaEJP/CCsYayopvpMVRfEawNF9ZFKv
wjr3hKZv4bSMglIjB9FpxTCexwDq5T8XjU6A8baAY3rbuLtgKopz6nqXhHj0OAnB
FvKefzEUFQJjrlncHkbiqrU5dJ1fjlbWd5Uz2MeboOjjACsSRd5gVeGzDexttwUp
rA+K/JrrSCzc+T070EgGg35jv76d8opVnqvShTzZJaXlRPqCZryUMSz3eCJS5iBa
7PHvTESiNkgAHMVPPLdxHpwQx1+magUPHgNp/c28x6nLwS8C82JF6jg31qt/ttZ9
Y+CTdQi7IbbeeekxTAfPX7v4e+SS5Nrw5kC1x4S7vTNMWm5errtMCUkUqnZ1GhSw
UthDYMym9/0uIXAoE78nqH7MLRviKPp9GGJkPSB+oUjKVlDSB7OpjXARQlb6hKrX
5nIswZNQG5yy0NGmT07rX3uRn+hWG/aFM85GI/d+oo0rO0LJRJKJ93tT/11BHwJg
WFs1CZcbK8hZ+Q7uzlLChK5+VmuXw5iXNnh8ksJczEjceuOJLR4Rj1vX0a7+Hl1W
R8IqhwPU+s/b7FVOjMCMlYoHamJH1msqBuLLhMJfaAxzGjCkM4E5nOIaMwznQ5RI
kEQVFmxv87+n459mOqKyBWGYbqN+fCu3Gm86ajGTE5uPYZG53sT6aDceCJBSDPFY
Kdz2KSaiNg12R7Q+mVnptia+YdRtcJdtwstM1/ULOvC38ZB+nEGSbtjrmlW2YZni
68EoULOCIGGbKUF+MOdjnVI9vRulFOOjr5tySOKEtF4YpyMkdx2fxixvBR4CGYm3
VUtdYrPb3qFrEHToCuzi6lJ5HCtm/4HUYiX6Jv+PvSMpVgZ8VSxd+zGm/8aF3c3e
cE2d0GafYUBCkhSuiFprbZuBL+GMICfIpuFb1EL9vcW/7BQUBIpSp8GpFVtqRRtv
o8VXrbVjj6EJOEzjg0XyGTbcwoXAQDOAXMiMnAE6W3tS/XsXpgP0smZ8ml/+Nnj4
5Nhs+uhIbe6usRmhUNfPCDCnoDVutjzLY7Y3uehBTr+MjQYmKMGLh0Bo1BWP/PEs
7Lmyw/3DslouqI0WppFpcJND42gpz07wH7495j/5+Lqmm3hsfgMJS1SMEaZVaXOK
W55IkzIxZpWMjRV+SO2mD4cviNgaXINyUmN01gHcL9ewB39oulW5/QDX5NTLMRJv
DksNS0r4UHJ4mWjQLmvfeykjrFDeNZJsseXHB6tiQyX0E6OzhIkLI9rQsX7LfWF7
WWnmyDwUhfaq3OIc9dvsadXIBBXKpfb6rU3gP/QR1UOPYm2xRRVmiUEVudZ0ilIu
2V3rnV7g1g0ZSYeCbxSySNvDobuztF/VI70G3jzWWwIk+Yemd7XvURjMAlu32C2o
py83Z3tFTDN7ChNijFLUwAk0/QRdLar5+UHp2JAYb7haJQTmK0rCegDeDVkHR7DU
Lp/dvxXgh0zTMGmva1ikqAfPb/Q4poM3l9g+16tVSm+eMyhM2SDLxp71FGWZH+9b
tKOMsbRZ+wYygK4qIyTcrVRimkgsFbONORTEusRlakXt+cZE9AEpN+sWWvK9aw+K
J+gDtxUcUoXg9JLhCcJB5v03q1oUMcoIAhl5MK3sePVy/3Y4BKyZkX4+gCXcq2Yw
DWABWs/mHKNqOEjQ9J4TfZPknERbNAocuALZwB9WMUXOYQjzz2P3qYOuzW+60+0I
h94xtYNC/7ryeuXN7mVLC6KOSIrui1iJFTLKg7ZFzBN0cUiGzxixSxy76ehvwEt+
EGzZL8DsYjBafzihnp4apQY/W0evpHEU6QQYUFXWw7KZXxJCoVp+mPReHTo+rpqf
XFCDUU3L1rl7Tu/hfuM7s4wZ69OPpTU9TnsqSXg9LYuhOf21wo51a8gDx9f7xNGo
lb8lbNZDGUcHU224IfERqwuFWv3CAy0uw+9aBXRqK6/bhFEsX/L9iwju5u4D4raa
IiHGtAwhxv+OrLRLmMmyrCf8yF6yioRKDIFj4+1gSSdzakQWhU84qTJVgrx1NNou
tmde0dOxAa+nTnYzzudYqlnwAvtovUBfRtjJc/YDtzK9fUIc6MsRq8Zl7+Jf6Hfd
bOd6vHfpCI+LZak1BOXp6nRLl3ay05chP1yYeJKEi/gGH76ww9pDQP7BE7ULZq5q
uxdpCkQYeU2+jQ91IKsLTt+ZiWU3HmtePT2fSEJpjxXgHL3d24WcRqWfHoIn8WiK
7ZtrQbR4Bzz8HsKP3R+8ocQ3kU8rygoKn3f4Nwk8Qx8rVGlu0iJ876vp1b3DKkCs
WQBcFhzfW0qmSJz3i/PuXrV9cNHh7RdFIAjuPnbj/jdL8EMpWRcD3XzhbLtTr0uS
t/2+zcuY+ngGkTg8undC00MsS1ZM6ll1kofawBiEFyz2hp/TgRuhN0FlDahjLiNb
csAupjLKPKfcPc7uz/+lzQ8eDzdn/yuIFstZykdmssJsT5Q6nsp8DcJDgpakYVPE
mJfvu/cibK6qFuWzfaxY/xieiRd+mKP4fRZ4O0IeCb7gR//392QD1tI+A/j2tEgM
xljd1NI4O8v9Go7VsZkHb9eMniaTFHThupCCILPVwVjKJzaZuevPJT9fsufgCL+o
JjJzDvrIio7ARtmOJmpVA1C9pkQJJ6z0c/bm3U7rI5Kq4ZvD4WfSeytVGnydZQq8
Ct+le3Qm7Dt9ytc8uBl7wpBDD4BqUbS6OlBbaYb6weS2hYXS84sjxpGRbE3E2oJx
dkZ7cBTCLwdA7CRDuQ1gEnADdgjpEshGO5S8oMXFu90aEyrRusVhPVNaK/CgjyhL
S/+Q5FJZAwq5pnZ5+MPQUHW42Hhn2fqI86/Cn4Qv5Dq1RuOYSARu3O03XIkvP7lX
q1BukgpTylRcp/q9xRZwqxS+6a2qdyuf46Hl2sspwKq9/SvBbfoNp1+pA59K9Z58
D9uI5ba78iH2K+dfdkIGZtmjWw4U1rJ2egpDzLuAthqFekpKMfwbSUTiW8z3/KaD
b7dLBMThezr4SLivtB7SkwjHI680ip2RYBuKutt/sZIhC7aEQZix96d1W1lS16Ak
fEFC6MI222uwrCvFoNr8Mnu6OMsDAskfmiaM+Z124RNWQfudqGYQHnYLD7V/+uv/
UBmrvNBH4vwXYnWzatfp6vZ/c0IQe61HR0GW8hlqC8AM8qN7dKAwOBhsAg6dlgZV
d9XeVdU968f0eiQEQPjuis9x2v0aOTJInE2aB1p5U6d2kumkyElBRmowK8lbtk9p
6vZAT/Mm7sqqhu4Z3yZz5i/NST5iR5rsMylj9IZ++gMo9Z1Qkx6vhv5Iqhs4F57g
7YJhleuz6PWJ0857dYaTSC8Yj10tR099ubvQfmrx8Af82Fp5e7lliL1v9s9M48eb
IAJWJV9vWRzziXxfC6e/k+pwc/UO601Sx3NawBprdEzwQ+AE/TgDSG4pjlgP2VZ3
ob93CLTHMfuOTosTVwmOVwPvvbb+gkLfv1oO2a/xgl2SlecHTkeHsVPBdbKdaOE5
NlIaQUHFyoJuo+2p2Nv09nPxDIy0a+IU0WC+S4ig8IFugPzGjkXt/HbOCnOEePkH
cwtYcALPP0iKym5ZflE1Qvo3pHhTsuPNDCy6bNTWbdY7+dl9vk8pXQ5ICfLtq4+/
WtjU4n2ZD6EHutYSbhcXrAdVMmANHOLEfBriwsn6uXxfxMWEY81jwVkcE1EpxhyL
Vc5N4GJbRi3vTOtcpoQJZ1yt1Tzzgb7GxEdly1wcOEnjCZ/pfsueqMHRHhx8OJUG
uy2mDMBxcoWxBRd8GlKZfu+R+2kNJUhBtRGFTD49QyQ0AmLdFWX4U1E7P3CnSPqv
MOwUPtYbig0nn3fn5TOGd6016RNe5HDcNzgtBO7duklYUWCJyoC7wdsxVdfqtQBX
V5dm+u+kfXCeA00DCgZ1jAsZ5Jy2fT70dysRivMYZLETJX08LpZSsRxf1EKT2954
vnX6lrsS1iZAcfR8I60gDyG7eyC2NBTWYo6/Llh8KeaTLc/M7p5ArCsrCge8gEF8
mDFoCCLVMhXALICYM0SV4TL6emtU2uXq48hbD/aMayk=
`protect end_protected