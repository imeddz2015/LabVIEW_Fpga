`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 1136 )
`protect data_block
XAYzcToIY1VIPqVIYOouMwaXR6+iabrWSAEf0x/eFj8GuEaEd0S1cjNRhN4pe3ey
dScutQVB7r/7WEWDYSh8KlQIia3LXI2SBE8xjX/tk5LCgNzhno9H5DapHBuHJsgO
EulfYGnLpOIT24L07xg5PyOpIldedlqGv3gPmRqNgcZIXqvqYDWgoHy2h4fE4WtN
vcvhRt1HViRaEp16/uomQT5Y4FQxLsizwLuJyAnrBoJTaH4ArETx8iojRXNIkBCQ
X/fohB7U9Jv6yAVkqJpjOl87UJnytpuEW1Q2EeGP9xvMF1EdpUAPXVQ5PakA6lGh
7686QQgf6QhbWTm0BxRspU1IZ7s+6ba2CcGRNgm9gDuTSN28sCmAr+J65asau6rL
QghCnmA4sACtNJ/wnA64yzPuhlRcYM9u3Ifx8tiD3ea8iEMU22IoJlUxQo1rfVqR
sNPWiFgt1NJ3Q0W4VWbiHpgYbYINu9TQOJ1/NKZj0pxLSE5xSDWmE8aEHaslKgm0
D77BuBgk1kLsmtsZ4HS7xuYbPnb2aT2Y2mmWA3JziKWmYlKxhw/BIPrq0U3mVWVH
abHvCRLNoCBZ5Mhtc2q1sYHrOAFtmBG67tpnlZzmxn0E+QvJLqWMucEv7Cenx6Dj
ci2Ua6KoITqNJkhPiF+c7w1cuuS+ALHtgoFRcmyQnxr4A+rExit3X2R6sOYWF7Wy
2A0BGmninVTqNrDhXsWRiSWYUD+EdoMpntGlpp7v16kTFIEEm6WvCLIIGJaAtz/6
RIt0pNlnEhRsrZjsscdtL4UFSuD/tVCnzcSAvzDuTzvpiI4Xuy0IywfEDFO2Ndeg
3IL30DJJWx1rh3xLF14PEGXTazq1fspeApJjr5QLmzDAQ6jtUVQYq7ecH7TXtnpC
0/3l0U1UstKkFGuViPDZl+e/UIOI428DP2l2a3RcJxITHVK5oP2WfvwViFTZt3sd
tlfSGQhP0d/xA18FvgiDED/361xRGrwB9YePifL8Cds6jONCNq/DzJhJNIR8KWAE
gwRGLeFQj109iAticEW/Airy8HLdRN55NCobJbAz4OAOCWb5kQ/R0N3cAb/1AZ6T
dK8akMYhY+IrJdjSSX2snM9hHJVkvL9yfYD1KD+AZkV1DzqYRtlnTtywW+CHYpqh
O1xjzggStoNFCw+zywsofvcn5F5UN72R/wHvA8y/QP9V0p4bpZBVru8aZh+rxnlM
uUOXwfCj0r7U/EF78e6InVRJQnFSMbbKcMSAMj7tKlZ4qlNCmVv6H1b9Xk/zW/gB
PXwX8xvORNoG+mRsv/ECoq/MVuc56d6cX/fxu3/JQjaERgnLzoEPYafrU2DmVB6U
50DI+inShAwvO7qN/5bEugqQTUwWRMYPwM5fJ4PxMuyShGlxqCLy28DwVh35y6vw
OqEX4A5TDtvzoExK8mM44V7NEfDDp0CnYaluSw/CbtFT8FTTd3BpZBMdA6V/AMUP
+TpaVOpD5R1DXo/r1X8NDBVb9UJLTyM8UYE4bnzahoE=
`protect end_protected