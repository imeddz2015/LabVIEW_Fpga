`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 18928 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/9huKRhRMtvnNqb3Z+UU7TahEoHV+T8U3P3ufru7l1O
3DlgtZzb9QxCbOjthp9+wDkjygH0eUfDrEl1ovhZG61SKKCLZRL4u9NFkwB7fCIP
miD1tVZOTTx0hT1mNQQiakbyGyCtakwPEY6099lnpo3IoYTH8SjXwPQc7kjkPToG
JIeq0jroGgXNK/e0gyHs62wIlgx/1rMvzd/VL20l1MbGSYMW6POdXxSgcZRiOUIh
cLjYMNdHcC0m6pLYF5N5fz8aZDdJo75LTqTVIavFmgPziS5Oh/6TxDX6wHiqm/pR
fN6r6GPZmyo86rKsiZxCtVDTD4PU7qAWi1HXmQLGWknc1M6x9m/CT64iNz7pAzWM
3QR/KorUKRqufEQWKlBqQp6dZpyh/lHwRvI+y8R7krSciWIZ1IwrQcEM1f5Q4CUm
DCcT7QUycOEaXX8a46C7UxXDTESmVewuqUDrCEITeMwfgTLdqWcvDWbUXlBVtN93
AQto9Gnbv+7AnpZuXg/AhwbA6VUloVb91cI8wTSpfEqj6jz0wc+qX0K3r8XYRQ1V
BbN6iUOT9yMxQA5X+SnpwaXL4K3ZcsCFB7bwPRnrpdP+JUApAVmxWAQBBEBO2tzM
9ESllYMPblgtzYRXWAeAYwC9smqrFRaKcxdCuuvDotskRmInxB4fGVTxJi05IvjJ
mvs+0oqP3N7OLo0lHYKqQUOkjfNKIg0ex9qfAManu7gpZPuPoefIrlEFVKXneDE+
6QruPX2JJXOUBy43h2LjvYNAwatFGzavGZItSWVBSLeGRXVfeHKlQUfKx/s1Cpzf
IGny8Jo1EVeRBZb8WY7w/5nhWKFvjxxEoCKjmZ4okM1cAramPRxC0lhiEcwZTbyV
/m4DhbDGDETKfeC24THyiVRQ602aXEzrgG1ieZFkLV11bxYUDxTFz6nfdq/jtPQI
ylR7mPokvOSZzyEbud6G3wf8qGti3Iu+R0qnIjvNWlBSjy3damY8q72NBnsysKop
8wATJLucjoL6KyccOzk1JK5Zeg6EMyKtcOT8qu7v5GfjwrYgqfg9uSKf/f+QLur8
6oATZoHn1YxZOzMqU1SfUUcbkmJtL3XfagHvPN93S2coucxxdHwStWfoC0voJnkQ
S4zWJTuuVRRQBADccTVN7FGqUgH0lKjK7O9+io1FJjjfEiYawPJAEM68gFWXwaOv
tDFHnOZb1pAkmRTKXmftReuL1Su1cpCPaifOch4YrWbrIWO+D+Jge+LImVsCJOhl
fKpH7SwAw58Vd7R1eKC3+C0bVW6f0Ez3+QOZ8SRO134DeakUL8u+HP2qRy14T0AX
e+8EEB+EFE9rGFBs/akpCXOan1oO+ckdYzo88QthfSKFQQHWx9jgJ+2tPUyX1hTA
Fnt3EMiEIff93QrVuDyIAib/IA7pgun0x7gKjUa84iVk+VF6hSzJ9lkW7BoICHKS
wGM/u5R0IsQMqhbZLgGeJqLcZAQVRqyZtv1bY0oSmuQuc6IGJXwMLnc8aBzdI5AT
AN82zB1DG68kocjQbMpHxu9gby4qmaRqW4XIgIYb947JzccjKGNBz6EH8ePCc2hd
qqrgfEcbTc8e4C4Rrv/G0TGGxJv9MMrhQjCkGUSz+po/vBoztpTkHXSDEiVwLseM
kJsW6rozQeOV3rmWmyp1s0RKENQfJAubz4oQoa+ZcX2YhkZBkSewb3xjqFbkuYdK
cqy3A+Gbx9QS5aTH700Tkxduyxx0FmsrVJ7V2IWHHcSTeTWv2O8aiJZu0JCnbNct
CsjSP2GYOy4EM8xTGJuy2SaOyixggtloA6ixcMU6NeDcEUHnenQfuauj3kWdRcoM
kL/e7iA4U8cuzoLauUDN5XSxowTmNw7p8/kFigmOpwI/fHC3pLnv6AzOfwW3SoKh
AKGGK5tJfd1ii0CLoSmhSRqRo0dF2gGiTaF9LK9FbKise8tnkvDDX51Ku7i0zOML
VDC08GHiRarq8hmD3mlAEzXxnTIeJiGzwXTWAFjHArJY2FDTKN/Y02Vhf62V0QZ9
pUzIdQkxzpub3eBOIfiXt/7XQQw1BlCzvj5SCiDui6iujgbmjROf8j1r10Rc/YJn
DcPp6pY2p5bJb1sfGTY7C9lfVpfV+REXFm+FFXTjvyfdEMf4oCqikNvZKQa0o+Tn
VyunDZZxVSMqVYp9X9gFOt8JFdCMwFvalLCk00q7yBty4X0LMLNFyHM3yhu0ftuh
hBXeEpEp0/5KfVn4PMrzo0AyfyJv8Q79ZwLR23/44hm36Ey2TscEi3yJofu2azMK
GjcNz/Lx38fTSbiEbP6jvp+T8pyeaQKSwLvmCJko50+CGT0xqGadQ8N4BhS16USm
B0vs3twc6RaC6PRIqA7bhVNmnpxS2d2Tt7apzv1EuxivOz35zTBIcRlHFLlbqSYB
RmIGPqiEIQJEQ25fJ0Wr9XUOxffAXk5/tUgkK9hkNBKSaKsLa6P3i8nIKfjDABUG
BIDTmV49tUGhnHilSkMqm3y8W+0d7tQPIP0EbOFrno6zl4tH7MAeGqsbwpyw36Bv
67z/Wto4qqCpkDY1UfxvTybbd3tz6T2ttIHRgCnEnjitcEdcTvAwspSW8dmKlnGZ
dGh6WO4uctKgsXPqQt4M+N8DATy4oIySMIH5SwLVl1DwWZIvNTlehd85fpirnCMs
GaRreE0JJ0NClFgGt8jndnWi0VgY8Lq5SAPOsBCbxZUv8WapdjGDdLjoO9svUTgw
/9kU7WB7iMWxQ9zWsREeRVfWpyd4R2u3MmVTpExW+Aq6JY0fkJ+Hk6o/Cvgo6Crp
yDybT95oGIWVsSvPJqb2V+O1/FWUXP8Vosq1JEyyg0i5PtouIjTYF4tGJUOWbOZO
mEZLLMAlYXmaO+dpjToREURlq1kbxksuFo80rSM8QUwmS220/iNQW1ezYCJEpXif
R8Ycyu4VmANfUnz1h8JAesXgg4yVqtCmOkch8CDYEurOo/GnXBHPiBLgmLT7WAfM
gOi3pqjYpVcyHVSu9jC6XPZfTEIIieX3OCPFhZZusxadiYcuaWzQCV/qXqZ6Zeq0
lXmY/cbImhgZAM/c5nYVTHVCHl39u54JBla+BDydSxJo8wKrDfoOMOlZmBc2kKPL
9cQkDL9AfwTrLR2ZlW9zbtntWGRMtv0q93zWycaKzWSQbtEKGZSMMkh2BR9LNq9N
TeK1xbPyw8OiayYhUlkzUmqhpdRz7nJh7MfLfufbLb9TKrpRB2RXc1f+kBBrfidM
TN7ARe97H+hj5HU6ES6MNukv8W8MbAQJNNDUNNoJjzZ2QHP7rUl0pZvzmR0P3rM1
hfQxCxEC9Y4Myi0mF4oJawzzCIRycY4euqRT8R38OOqZGYHU4VxvcILYg6gaCsXs
w0ReNdRH/Ko5NG7dfV6Fdjyfs5X4JjBgnhyuuiffwXuPrPqSRelJ92KwhVereI5Y
EYPL02DKpFXYn9DVScxmfDeaIZIbRwTIPovaYJDEDHdMcDLWdLuYa3OAJ+WrL8j4
Vx94Gk73AjtUQACv7qNf9OWqlkXw/F0lTEc37jo54n7g1PLipikvaVN0mTWvD2GM
6qZ7MNXbSkdqryIBhQYgzuLb8nR38zk2cvPcl1HGWuh5WPjSB0gy0tIlWDoBWNOd
UHDKjzeX0rRmMxok+E2dBTsQRDcwKdNCDgrwrEDmamgU0d6JIBIaa0NZUNMI/nd4
5N04YWD2bv5Elnsz90kARMVhCZgvk8xEyJ/K1o9zCbLEMPbWZscavsmE5wVYXga3
c+f2vB5/G7GeK2phVDj9LHBAxZs7GTBLy7wP//372Q59t7ouLeQTKMrRDQ0t9Mw6
Per8jTnKaln/sxUq9GF74shxvZtDytCppya/+znS0gEdXn27TqJXMXy7ktzzr1yX
bgS6QIdEdk+VE2jPTumH7m+ns93EiX8PJQcDEFLRAPsBTqxAv4m6uCWW9MN6OXyi
Sds5bQ9j/xoLUQndr7hvZDnvi/V1QuQBVGPmQc9KfjxpgcBy0AOwkE+kcla4xRX7
fZtiTOTB8Jbo73DbY97Z7gKcwPyXVw+IjNfxsBV81OJ32Q+rSsmbqH/Bylg0vDeF
Aox4vQI9N6gU3Eb1GRVP7zVrLDyBYWHQkCIYD16bv4glDIiZirq1N6lAJ2UPtI+a
JL+jn/oE1PIzQTlGVOn8yorlTurO77cCaEBP+ivt5JnxzVSbUfUj2kwuKSmNc+O0
8Xj10LTNJQR9pN+6bnP9XBh+xQ6z8sqXw2F3JO2lnwol2DlBhd3JvdvNaDBdQTDw
kIVvUF4XbYXzfATeqwKCduavWjIdDrwC00PlbHlFxJQRja7ILkHPE47TtJTYbIbA
V0WE4qpKczd/D/JDNduME/AvifXO1iFHllqmvlJ8KmPicD+I9WawnUM9KGJpHUUl
XDlRxGnOEIujGqON9ksiD5DENm/6u+UnmO3xsQU1d3Rwh9pFrIVP8nf133veCtBT
4Ud0V9fbxonzhfFzrcMJwjdDp8Pt7cWpl395Tt9cWQy2NsaVJ8wNU2BMfx2lMYjr
vtoDE90Bl94RCZ9LHZ3YcyYo/Wh6XvBUuWdjB9QoWH+xCBfV+EccpJSuVoMpAJp5
eRfRqkFRPad6JqCGVnICv7b1/19ON6VfJYW52ddC4z2jl3EjlfRfQhbuwQ1WaXqK
tHad1D4B2GEe+jJ2m4PecGo0OUfKZSU2s5RO27JvBaVdMsQQc7NCr5QAbsvcnJJ4
FM16XFuBZPyyPTLWWQLZuuFoY2rAilW0UgbVYHMrkPMrtx3LOKQQrXjvTH+smpaL
oJaQq/I45zGkdflsGH9qtmFAbg2MVUgKH7ho5pzo7lkZi/XU7D8m0aFLiHiod01v
Ow9oSX8S1o1vgUBK7h7gSVXcE/M0lLnIFNcvwqjGSlIpgqX3cH/i70jmL/AUX+ny
TFj6SqHYlYJTJmcKb57tWKpvdCt51z+AmlaGkrrDTAZ7s9caCQdAyRGQ0msDA3e2
N7uwFDMB4C7iuZKJP21MQpZsf1Akah3eARZ04GRzBVR0nyuxNe/A51JzqNhLhIqG
EOJWDcmVsgEdfFY3WAFyblNMgJConnS0YUUGBqgUssejj6qw/YgDm0LlHhAfC/fb
M1KJKzshB7cLiE5TTyfRWnR3Wr6hbyuzZHZGWyfAVWZgD7Pi5Qu3bxeQ9wjW7TwL
HI+s1ce1pIXnGxlm/GmBpegdXqjhkq3eeQzLqmoZIbO27EZDH/lHyqDsmJzRg3Se
uAUcQ7Jj/FNOpd+E09dMWw2KFLadzrSmrf1eSGcKhUFRVX07w3hhRfDDZEk+/4j0
rIFY49Ppcrp0SHDvGBa5Zhr38nmtUaJq54nd5QAnoHy0LiAoedsVTWwyQxeih9h5
dWXmJQ48OxJNS7nvGPhHpFhGkvIHXwclyCoTpJMWiJfR6MZ973q9/npRS9ZvJd90
U/dXDOdGfYBKFIv/K+xTnkorr/2lJBetPw+315llgHrSWfDkIyCZBLKzZCP/98zF
62aBYm8RSx9Kly6n9rOfdt0o22KXj3jYJUXK1AC6mfFQwykKYSZvscQ3d2V5cqHP
C+CStt5Jh5em8KWqYkRZ772L0bLaixtjZ1sQfgmqK3GU31zpb+vSP2Lny45gF7bk
tDDY9BfAfn5nJiDGQfyY5r7Uv5tIsKnt6Sbc1GlMZhDvquT3FgUqf6vNWuiUw4mQ
gfuV0eM+WIyAYEbwl42ZlMTcVBBjCGeYsIpgcSNxlPjy+bh4QhZ2pNG6vhrXopOe
qa0G/nOgi2ljOl4jj4ApPqds0Ai0NoUL+vi3QUt094FNUbo7WxdmIsP/ozWEUE20
HFgUib9n+sUcflrBHjAE+OSsFYXdAY+d/xlwRBR4s3ZJNQu6OHUDgLCPAdRVFnGC
9Eo3BCLagjSgrA1voCKVnClggR8BpBdUym+P4J2siR+ceF3VztNIzegiOe/V1QXi
EMow39nCJKnjQitcexN9kdqNR45FJdXaui34UNZbeIeOS0Gr5utM8vJI5nutaO6s
8MfsjRjyU6M8lGLJdtvfVBm3mmdr9LhhYY892w+Te8FCV+0fN/Hj9Ea8/9/JUm7O
SpMKOva4tRL+g29h8ZmMebasAbrFzPnECmxzN1Y8GvPLTxicMxcCX7R+tL8qCf8Y
5VtBo7ZAUXSHAD/NqF2AT6VCHPW/9Bh6DSRefqbklkssrc691TG3iCUMaT0Mp1qs
EX9KYC+W8HgOZA4iHtj18KqvG1fFNDB1aYOWBSydDEGqHx9cbj5Rc+pNbK3bRBuJ
EvMF1GquUIF1VSvdsQjhUb55gjkgn4F6r69ykj4H2GDUSoqjIgED6zHPJvk1jXNH
UxqHrnGaUqS96YS2jluvVyDGcBFx4MfbotBEDuA9DWZTfyeAqyaEiULFBR119HEO
RxZxiDqD/5r9XEf4PCUhSejLoGQkSENwxvXmju+qNL47djG869bt77HlBPkhCJg2
KqTHxTD57KfIGIdF+OGCjOxhTHcVJBRFYDK7xNapRSCZmce3Z9LsP8cIS7W7DN2h
M2FdbVWCOROAqGw51CywLQ082Dk+wen88nRgyxxR/Cg/SoLdYK+X6X44AYEptvAE
iOmDtPQsQTrQcemrPryQaL3hGyBbJWM2DcJM3zU5CIN3wAQLnwmYlsbilYPc/hl+
JnNNepHtecgtkQytI+4Y7k5v7ZhheS7PR/heysWD5MjF7YiWFo4NwLorX87m2Nsk
Yd1gRQJnfCHIzwnNzgOsTmr7+mRgUe16QFjf/nsayjjjb1BZXk0o3qMJ5qpLwxPe
il/g/4F/gnSJ2ipDlotjpu87rQd19Tm/1r0E6jw8SUKH5CE6Q2I53CYVMehfvLBD
LA72ySlRcrYG+9JKUEbp4YBy6IVd2G///I98ecjQOonrlrt0/qRkh/KwBG5F/gme
6rFOqNek8t1wFOGnlt9c+8cpru0X8q0YXKccNXy+Xm2ZxuvJjoALeqe8cIFg5rt4
JvVgM7w3vlftIvkVNSKlzFEkNIr56PRhPrPTQSTdosz5SZq6HGT88AMek4uDlOpu
1NbiJoZCn2Iz8rfsl4FU93HwDy3w12xYqgVaHQk7I0XLIFYSKu8mxhB/j8Mq4bSy
NxtYRV2+mtXC6FYIqopW1fEac1V4uUxViQpXdQ/9IwrMstRcC7QBPdeY56M9BtFv
KdHZgBvVgtThcNSEU8WDXm7wrHXGEUcS9YavrhPyvS5xhKvapErJlmTXP2hpJCVg
155kaCFRcrbnqwhnTN/dNjuxu3DUY5ji1u5Min0VTHPAuCopbwl8psRmI9y96nYf
XPfiyzpG8Vc11F/RM0MeV57kEPqX/GQJYkpmEeqBAV6URKST3sCG5V8L6/es1J6L
ELYzBnr6tkqrvaFJQjdmaAKUKz36y5YZDmQPJ75SCN/O4AFvDQ5+K32uoJ1bBAej
YbYcaPNaSXnY3xdBUcJ+nnizXigz31PHwLF1BKn+G+PIYWTSQqptg1mH4O3veXCl
4noqqUcB2pAv6Y7ODJFhnc2c2XnRhpWog53IFVRQq9rkxV/FFAoVSZ7taEv2VtZx
QtBes1zkng6vuUmQk/Rb4sHm9KbdAvRRqr/wTbQbKQLRAP8Aj7CbR+yzGVB4hlpR
Dsqe5Z+aCOS5jJcaJUcobdhORXKmlynfMj7iU694T7kB6W1FS5aIIisXNsXqJCx4
7VfpMPEUh1kNXa472u/xK1o+M0RLVCHYaBWNzHfvIHfv9VEYxwZQ/v0pwWGdV18Y
xUJKDqaijXTaO7NEyLvOKjv4BIczm5Cw/S2Rt/5wyFC4RDCcR7hq0PJwMmnvv5pR
9UKg8qv0MLChrs7NT/Ll0Lcil7FYPNnmR8zfGdYuArOULvke+sFnOYKexVnwYN4r
0w7enLIhs72PbRXR2pNX891wBSBV6E3PKdLWIvZPkzNBlpeKkvutkccmozchmcXR
HVI9vZK9yJcur/OQrDVWl8dr0kgWhRul4eOeOVnRqXJi5fR1L0aEUANqpNYurK08
IimBvbqSLuMCeClxzLLwsw9fQ3JM4oCX7rp4QlfIeLCjQRXdorTGDrNggaDXTErJ
DVOrn2CDkKSWrdMiYFS5H6sTNANrLBTwhOCgjy8kWLdIkDVzDGTh3iGNsn2F45LI
qSTnnIfCUuqtdlTM4oQMVm7kUZxvsXH0qGAWkgCY062Mg+K9cY4LOpaC6DHvxIo2
d02Vihkz/8K27vhC+eCCpiBH1VbBPnI0TxP70rgJ+EmL/llgp+16O+WUfSgwQV9t
z/cqklh2qCEAS0lADdGh2Mp5CNsrhMwhomCUEbGJGX8TnoyGNui96JF1tvfnaZs7
D8fTGm99I35WgXoAIkefqPtMOIErxPRkdSC+DwRv1CAXaYOvQBkiZICTetDzShLB
kQ6NltWP/vaypWV3tRr9fnRuh80sVJ/Sexsp8dAHmsN+SSKiDIqRGCnDAYD82Cth
9J+i+Xq8RfI0/rqPojGq+E3BDFvAfxsYIvWDaKrGHoJ7g5S4zkoyTRQF3U6wxRQ/
X8yfBBLiLB6FwpSASDKcvR4pWPm+m3erXlDsiomF5dPuYbGGjblnNgmG0pqrwVc7
HgTazSD+bTImNkDdkTcNZ6jTtKpEK6hWs3StgzYVChQnuWIdhg/ukYFyPPhdGGVO
8vgn3n6jh0kUguBaxADF9uwRoxoymwAVrvp4H7z2s4N09VWNo8TjHGD/hUOVuGzm
/jM5mkSk8MS42+58oj6WmCODSI07N2eD5D18MXNXeY92/pqeWrMRzckAm1ZjIcj1
OHVmTbyBh/Fx/8amz2RD/oc5xlT1N7yLtuEBMYZI0p1dY9dzND94ycX6mfdRorat
50YehunkGsxjjSK1zivXycBS3v2J7ONGqCj5tLaUSoS8quYmwbm86UdiDiQzPgj6
4ifLLuDC8cke0rTc4SJYWFW0OKyw797qJRztkgTkPle7yjm2ONqdnOL44VHcP6fX
XmJTeyXCkECXl8cR2EpN9O+jU74CsX2uwxwmoE5v2RQRYFVMFi/cxOROEMevCuJK
bDFvnUKBMlQlKO1RbjZdT7TRYmCWamd740d/h/AB+WNUfGeK60EeTHTLzyWpWFua
coccaY5WPzZYF4YTaueWzybwuZ6Ld9HwS8Gx4ae9JLpq0qBTBvx7xyIvry/8KJM0
W4kr0FeyLnin6bWRCX5FgXCSGiwt4usgk/MxAv5ULh18/l+P08L8FHCCcIZrawJl
L0EidaVMuOULox0Mq9wc2BxPIw7wAII5aYxjCFuUfKlK5drKJ0FH19CzHt3/D4XC
QqScsi8IB2xfts88tiUJT0ARXVCZ5UeLlrnN11fVIBjvmQJNjXZ8//8ry4tPVu0o
/5rOAc3en3plpsmcisfRVFt+YG4z8eQJH+yIZ9j8fgQ5Xq0aAC7pfhKiurIP9XzO
kM6gmCLspkfz9Fpt80QhgW0j91zLbzb4pgg9UZ62vO2+Fw3iBx5nJuIXm9x7N54B
HL+z6uDwvnldMo+4jnrsX1jynVjLuh4TCIlkpCMkgqy9dOqJWrhOc5JuNxQkTqD9
Hk0bpssgoaDK4fLYVO3cQmZAqE05yH4UliTDKZBIDYGi/SGnbKaSjIkhdVxWWnYw
qTLc0xRrh8vtgdE+uQJ5OkUb1H/dm175YHkE1LyboZXytypZsstLy6uHDt9ZfOM8
oLI4ZfAhA0Ha92TsxYQWDM0udTvZOIe0sZTH08WsW7IRMhm1uulfBtBTUsUHv4pT
wBicFONI2LUN3mEJoX9Yg75pXgM6rAO64M5wrZFChHncYp/Pim8H61JbOpm0vfzD
3nAB2xaf95dombT8ZATJnox8O8TGQqha6SeHCzvlSnCHYfi9vzHcsgEFJqwZ1U17
+XSl0JtbAzqjXzxAS9JJsqW2/z8I8RoAnR+7b5yV+OJ+Dyckap4EuW1OaUJBw8Jx
+C5pPDG2h99m1VMniLuDjpS6i6n2gu1gKO7SJIBxs4btcjCLO7Q2KmVmSmfoJNNo
QHh1AGYDF9Ki+p5BGMEbO8sF4VXLjOf7w0x8pUo2fWCsk3NwL9mldTrF67MTqH/U
FstkSEeT0g3D+kM9RJG3DunGLkWc45JXk0eUSKCUYB9XKVh9PsMuNDLnHXlyNxKT
XkcNkTdKKuDG+cjKvcpadLbMBPtJJwG+n5zz55zRVyXz3m+0d9/ne/obdZIpt6i7
zCYeFWxbQmxBHnOHxfv/F6HWCedUxsChgWHcYlUde9pKCBTzG/fIAgMsBD1nCPGn
xtBckVB94nE0+6lK75bdBuwUfgBtKqVZQO4jmHfhjkC4/aQNVxiPyUSXqHxXsXQW
oWbfCu0e91Np8TXxJLJCVHev0UCe7Pdr97aSCWFfxKnHet3AhH6PyTg65Ew4FY/6
E+kXg+eD/2qR9pZIg7Kh2f2zY/UgwV5viQI7LvkPXKyT3bcYaKgIet7QhXGIxHa+
JeaX00F6A4iy/UcfxcpWPSfmvR+zdU2vFvLShBgPJsn6JEGHKtL+6+CFP5we35Cj
XVGDcHGb0CjDg1reY6lngcr6f6LVedXD27W9F0g76TpnBGWLw3D0Ovc8RsAcQQnc
DYEQNdx8SXqb+/ZMCUNRduDTQJbZ8q2swEuAfCsTQKY2wxpzr1XNa5biPojBqZEw
MzArpHjvTHgmk9guzGNZ2vi1Kp1KesNk3N+Q1C+t0JDxKAAZ79x0lbNHzn0CcXdF
wouXV2GyzGcMFfcFqr4JR0az6iWqYLw+s/8Vn7LjZc4T2afNNR6zFoWjo6luwRoq
5tVsSP5C/UnUrs+IsHNH/MyP/AiiMUl0qVxJsuXa5q4jzL/A3ptBMVLU81h87b47
Vxu73lz2fZekyFubzlCfiNIeTOlhBXU1scCzLxcxGdkcpznGq5BEYQmsRRRJZKC/
aveMiXU4HTOvWlqNnUQcI4vhZKHPY3Cf1OYrlFQLUeBmInXXcPkW9PLlqqQhj1y8
pcOqj+53mv5uNoDWurEWdO9ApSuqLq909KPGdKHXDD2WIYCTlMv5Wz+XBPNYq3bv
7SpMFJgY2Xvqd6vzLIhWMEirECdjzl5XoNC2rvCzV/Ivi+lSO1gCUgjxgmhyoztQ
qZyN/TGWSoeKs0xkMOB6xVkvZSAjql0pMvMR59NNs7pe+m9TDLX1TuL8RRn1GOZW
CGclgSGn7EtuAeseKEcQixHqFQK17d90ZO07KOoprlGnY+mYkcfB7cc0C+oF5gOr
9kL9O/Gezc0xMDoS+kfy1h42THlvg5Oz8t6FvJubK8TD4M5nAfadhdZ1zQM7F9DY
G4JCARQLv+tiaKOEM72YDpSPUY830S3QBpGEJ5MEB8txD2c43hjLpSH3xzrFJ3kQ
1hlRmXVzMiTm8DhCCzdvPXJnyoCYFTXP2r4nv79k9GjBzIDxVPKC5b4EnQmAm+eW
KssZ4u51WKfEm0qDoX1UW/g3zICAxzILNgOPYxVn0/qoTMLW8xyOCIfakdH6y8Ho
hN+4VKCvvOWMCmAr2CIZOdiO0aQAkOkz+TbqeqhY8bFcBCtzEK8MzYd2xLRrwqdh
Zegp7ASBkuoKsVDEENDdYAKYUJNXNWQr0LOyqyqrpBPXayYTrSZ6ZQ6BHmfrVa7C
PhcTigEZJfY0AwbgTeaRqCs00zKMpeUH+6ywEzLYOJpYp1+zlR+F79umQu46urW5
0vRUfZMLNQJY0Dwn3+l/Tkjtydancq4vDpZKVuyxFUMNn8MRAu2eZhrrxZBq13XI
iZsFmNp0mJPK0o+TnNoEMAkXRLKRdffQS4QqoXYwUICIUjRGdIzXp9+Oi5j8kbu7
N8LKLRW3j3hayS01nreFaBEdnvKzJgb4TQ/Yf/pDFLjI6CAjSWHCkV6kWrGtC2Jr
YtZMgNawrMaZlLbZKUbeGfzzwO/RGmaEnr2tMgujfVwq7B/6jMTto8DFdiBpzPuQ
Z2vp+8AZv5K3b1lZWxr/mJyhYLGJSbm4CAR98qUXFEJcwRzwcm1M30ygnVclheel
A79iiUyx4uW5VnAbxlLq2Cd2nCmM5yzdfebPmkYLasfPaWyIaQeDIpj31ORn9x3v
/5wNAcdr3gyRGBchuah3i/+9r80+1auIznUX/6qe8QThum+GGZGSZRlcxF5SUbeG
Aw+Kv2b25p2xBTdsaTcTg4TYd6Am2G17og/dQ6Wtomd9Xz3Bfi4ryYvm8DgwW+c9
1k60YdRSlcDU7NWV/LTKTO2Tmxb7pxsvkJ0GWv/FP0sAd/5Pqm3Wzywj/2jCeSHv
zEKUFAKATTvPPVD/H0mzTIcD112q5JhqFnY+DOOrHOXEqrNHEBdgJqDf+oBcjKiD
hC9ZeAXaP+F582f7OwfQ+EzX2BJlK7yKq0k1nfoxh4pG29knV+ow7vdwwuQzZEKS
f9mg/M0/2QEyVgeemN9fGO7+P/pBiAOnRBr+1QTq2nxSk66m0EgIKS7SO8DkNPjh
jHMRMFvIHqgmY8lfNwEqwYZScuuOkkVtvWlJX++CC1//C1Ej126A2BCj07HbpHAr
P4tBUMGn+P/8KvGklMrDg9IeSMF3BFGx10MuqM327uI7ELpwQ3pUilua7FwaxO5m
rajuYX2LBVUSxG7X6gD6k1sP+RqE3/dbgCJ+z8OZBiWIsVyn6kM5i8PnqwHiyFp2
X71mn1mu0CtKue4/972okNbhhlSDODfIHcgT3sXLVEjd4Gtf2N7MSiyQFO2Uf132
0n5zxiig9EB4JJA8DxnfJEQ94M/z3EFlLvgEnMaDFxtrDjfb7vz8FpdWKuGfDb8V
ulRYCINt8SDh75x2dai8F5LdSG4g2VZDNSrdeZyrq64GMIVycZxgiQo0Uw4Mzksc
li9qKD0FXrAxzx3oqtHu74+m2dflbha1MNaIeNqumAtMjmx+TgTWIe+IfUAhScdR
SJ8oXYfYHdBUxhT5KEEwFAxK+XQbSd+Bx4pT8CxtP+WDZYZfWqxYSR8QKQaV9/84
ev+aBouODG4sHtNT1gqyBkESYsI4LB1CxQed9jrifU98kYYD6VxTuD7Dbz2FL7ig
+cnrJ4JqWyhSbSE6rMOYvSU8IGF+wo3h3+3t5dnyA71loLCCh7zwtpIhCchjvKxt
mqxiJ8Oc9yyIPNPpehv25TZhWUEAjwof1fP6uMaWWXFzF0KJk9fIfpyc/BOjdJM2
M8MeI3V2xn+GpgrFU1d52oT67zkh1Ccq3fK5YxNRIa7KWqKUYlEGp6Jvl3kVfkZQ
0+q4SvLuzRqYk+/BarOTXUKyHdkZxvhfoVDzsBQGHY0k/fLPfYZUpw7UdYxWr2OH
eCQysDLdM7qAM2t5BNbasEoA7040ALb3Tuac+lNg4sobwe52+z/y8/8W65jJGXzv
WojlpsmKoCltPFCmY3d4/eCUoqlbsleF3KRvV3J50sj3eDWPkNFFaVJf1R6Sb8c2
w8jkODxHbJLLujPe82PNj42Y/m1Ae2DEMX8gzUaTpAJyl8uvvy/hPhalv2EgGPOV
jhx7DatWlcEI7yqDBLopveU5su8YU+VWRAeicqkB9vj1aJeFeeOgDuYjTRyMvkxg
RwzKoaJoXD0rcZ3gV/LQhGyyUI9Saa2GA0fGpI/gEIZ1g45ksTVObuDaCshjXuoL
VJr4iHvdSMLjvEmRKp4KLUVnRiIbwkb/Xto1htm6Fxp+lKt5ilYg+6O5M5yRBRa9
Iv7bfrNiEsqES3zRgEFed5DhN9Gd1sVHe/yLu6/infY838JZboRlb97cBL/SVEkt
Tixeppctr0thvMedbXaDk3gjbWgWAJWFpEk/+HKtao1fAyeDpxG4jN9WGUhC3nMP
+4x+vD2uSQDYi3DSqBaIoLANLT+bPDw9evIzirqCpko4u46Gk7QKIF8huwL8pzb/
2fKwgDnmAj3xGjIaFK/URQkWrDYnBiNeWBp8uwEhceTlHeVMX8esbPoPaY6Rp4pT
4VuACKFw/vCVFpL+ZSQ/mVC2IaRzs//uHUJIvnGAdC04ZEozydqacBnthGVQckdi
TzVj8TgtLF0dnSy4AyXhmzlaEo9qZrTwMBtXdax4xYj1yspBbwF8+1X+nUyFbjxf
Oh6vJAMlBa4c8hV9duqmWxLjDDiUXDm+S2CVF7XdG5jKXS3rYoaTo7nAnUMLPVcr
m/awYggP/8UWbdEIDN3nvu1fs2F93/SBS6YqpiB8hCFzejfO+clKZZ/0xlxdK8rQ
R1aUceVRy1c/hJjEfbsxcTtXuQjbvVSjungHDrfWPxa3uRkWKaFHmMroucob4hkL
fQ4cSEIZ9jxZABxHeTDU1pfe2z+k2o+ZfHq8LEjcVogFkR7ryOBXoh6BB6Hq5prN
q9sKidQ0fMIgU0YN55yJy/gDnmqysQUgIounDCGJqUMB5zDy93LEOMzN7amcFOi2
v94C7+5ZkxqMw+bXHa5GXSEDPcva+6Q4opoHrEEl9OWsRQ01ihCuBkhmfl4eFDjX
fH88ZIjUMxcg9hOrlNMz5cx6zj2GmjIDajtmIsU8sUUKWVCCGJZH60doVlVukZBN
snmwNbhKW0BNEFclApRbsFoXDX0aoYaqIS9ybfpmOoiNVYDm8tpKFkySsHvwXiL9
pzm6PtD3ccBNjVWOFnnA5eFvAlLE+PSTqc6+y08dQlPU3FFuxGS5JjwS4glTgOoi
WMlk5fKpdDMIOiYHo6FucHKVuZqFOjvdwXEmDbp8fEwSISSHVWUYzXg85szHFAT7
qmSn6ACy4LTNripJxxUVerUHPGDaX75XnjrGC/qdDOTE4tO7d8PJTH1GMqAHWrFS
DHVeS+aa2/z4enNjJtuwbX7xpjEYuVxdLyHDD4FGH193rC5fO0brd/vSnFlIqm8q
YyjdIRi/qw4gn1ngPZ/SrgBHylMY+DmEJfoe5kcOWlfMft+4wGYLtydyWigcUIRg
eUvP8gj5e3awmM3IMjxa9LRt+JT1goEumyjo1FQ8k9ITaRC6ecdRIBV2yWTKqAae
CF1UTm8h7d+ah3woE7ZvJFJDrsjn70HIgJo6SgMzgfwlxyhOtvFshWhFfNivEqWn
D41Ohi9KPO1yZgKIa6si4T8y0jklBG7tmO93+alzY814NsfgErU3Yl87al8oP37w
jYeBMtXxXHPEWmFztpe3MZgYvJVxTPDa+VdG9e4VzHMc54nYdx07j0oHk7Wi2BTm
uaQ21JlLCMi+Df/uyx7MFTKTU3J4Q9vIjb8dJeD2VUqEFhRRexVFGxeOL5YFtie4
H9dZcVFrShYL9yIN9AfiB5lUxCcaahp3mRAfyn6erG17cUXc7/jPp/a457w1zxbD
Wl8fOGjg/XY3hIpJHjBxEXgaxwezdwIVjZuf98bFGuzqVfCXaElWdijAAZMQOucm
ckSApApGRCog1r1mlix5dVhe8hEDdES3l7MGUCZ6vXe1a11l45MWht7Ft6MvTjEx
m83wYuYSGxuycTB6FSjkI+pCP1bj4dkVsYAnObccRJApjRO2YOUgeIl9Y3WLv3au
1AZcxmGDutCxyMV6ywMFuh9sDD7gdwGiP/t5mlj2kcwKnLD5DxNsxdRsrSPVzDlg
eLYFbtqYDW2hcuYq1rghjAUym+nxr1CKvrGvtHgZondNAQZwRb4vk/H/EAsyvtOX
B0lzkvwFrjm3k+n05N39CXCwpS8ecNA+i7QJstPg0/uLjf+nrQYO55l/gOoVAwWC
D4ltBFiXWbXk+lPWBwVF0LtXoHhIxS1qvDj2O0n8DKIS+uZtP7OlbFd7D2TQaBoI
SSKd2ip29LyvLmSK97Tx6MulvuEV12t4VBTtPq8q55F+OZ2x44FZVHLLlAMSFuV7
I+ZLU0kO1FI4ylV/XVNEf6JaJADkFvawzMtQPn7A7jIDxVSB5qZrFOYpICxAZoaD
U7TTs+6v7PiDukH/252WR9i+YuQ6ekS0vZrN2b5NydoIojkha/Gtvsz0OT4CvWNv
y+nVRJwiSXvy14tA8SBtQ76NWzjimu893+wPlyUVsxkmTBfvwCvbinGFlp6Xr5pT
VALyXJwIfn3bwSvMmvlg2Zt9lec60MkUOgP2weRGDDFQISvXweucF2gnhScQ2hhK
Q0wJ/OBQAKjOOx8HwR1N7himUk3V1ha7RwOFxNzkN/C6sH7EzeHOi21KqcjmAi4H
JrdiEdmsBJUHCeJYYAugD0hmOn32EpKub4jEcR6wB75iKFfSC8CQEDE14f4NKkxe
bcQHsae0Eh4hIy19aLntKwmd16zU3CfxrSGa4DldPdyyLuTJqBxBVqzf5VCLbmB/
+hktzF0W8FyaCSF0R/Ckhqahb+mO7GU+zMfsuwpI8+4SUIpf75eN2aQiM4xgFbN1
uUebDTsFM73o/RTiW94pZiqeq3uSpDoUHTuE4r2AlCKNhghYzImo4b33Eu3jmIqR
7mS4rL36intrjNclHZ5TgqnQi7MUJ989nWU+o3f66NKIy2nKCv4HOLlGvADGpB2c
3jSYxsQPXbhweWPxFOO30LOU2emlo1+/isVy1RSDR1c7vX0Xlucdpi3sE1tSCh/p
L2YMoOwV5mIDkY6r8QOSc9CeS2JGI42AEedSuTxsX5Py1CAdtulV14Mg6eaoHA/H
nAbWAxXuQ0n1wBu43xzomtHzO5Cv4aEKdqz2bDBf5r49oQ+VThX8vuRs2jA/hvvM
OKYLMc8xAR2PI/nzDy+ehbSR5xRUSMyG4cupZ6XtuBsY/iYRvttiPlR2r92JTpNj
t2xMZZh0hBFp6aMjA5NVEX93LlmRREYyniXYEJESws7oHZFAm+mRVGbLqbcLtpZL
qnQQjNvJVKhX7BXf7JVu9go9HEOOo76GR26Xa6uuEDoeOijYgO81S23/wvrpaJsu
RCWlzjxwIQMve27O44hpqen3jjKzc1ejtARP2igOM5cW/c1YEaV7Y5MYsqjSCUKi
mnT3vII8D38/SqF0bsohWp2fI59rGvMCD9//+NzzFAdBHI8dccOgYP7T7GcfkDuv
jz+z4PxjgyzFBgn58WGtk4P9NKCXiU+23th7bu+S+cuVnJMnDo0LyOUU3Wl/FTXx
ZP7HShDM7I/cg4aY9KAsfMdUNmDaO9m5eQJ0TuCdGjHI9QyHGAvI6u2liLyhpEpP
Y6FKXtgHQYLbfobK/xGeFpE0acrdOpDEfDYNI3s9dP6u2BvWG8E1eYi0l0YW7znJ
RoEBGoit0LxCSuLgNvm/kU9UZXV5e+waOGqwQt7mXPjT6zWitbD4VI58XPgdRVhq
dTMc4CHKm4PL1ccMKEy+FYEhIzNObYr5oQ5a2v9np6TTGDhJuE++WuNhXaNn2TYF
Qiy480zWkVrzHKRn6lafatH5vuUOFyqsQDymqGZ0KN2g0lzm7/0hHSsfrUEepYF+
68vCjibsfSzEGFlazcYdEl+lBAhJTS+K4LzKMoHXGofMf2RkSC74FQMUv4hLU3iQ
WWOY73F/FBiVy4GWZFkVmX9Wx/G0i0OTnc0i24XDXmAz8tXBv2vwDTb3urlKvp/H
dsFOI0/O60Wm6e1NxVOzlKHBIL6y+v4UGv8YAIoWAJxUQrmY15hOBE0QeLlWJ5fK
QrarzDFcb9Ih2G+Bmp/0NSrkUd5jFcWnFOHrICF1kFdbyF4buN37Nd6doGih/PAA
CoHLy5PlKuzJBeapZlajNfrcEfVkGAnbzas+Xgb6pdKjVn85jySLBV8V6XLogDLm
iew5MvTOLIzgZoHBY4NGLdoYWM4D1H/wiI4BSvgoxENN6bA/RPL0wOwDbzYakk3n
amVjdb2vqUkASMgA5mYhLlKcaYs9QGlVcAPDFefd9OSIs7R8yVyrDXoscHfLzc0O
kou2CuaqXpLCSQGW4sNpPwm1Ii118atRTt4qBmZtjeoKly/CauEqbVxSkwpau17F
5AAwkcB56Ew5NPi57XjxPTFaQDvk6BwKOIhtS92aBCXW+StvHEzF5fPgu70PP878
vjs/1HHmK4bqbjE3zZkRpopUDVddXvqCzga2DutEpjY1MNVIKBrSsK+xucooRRB9
sjC86qrRxo7qowQHbV+oJaJocXWaIGOiFfLfcMISQcLd0Y22vW5Da/JcXVWIumRK
0JWo/bSFUIqlcOOFSG7ME6rs+Xly9BaXrYagSRHm+OVEsG5p6+1m5Fq/AFb2mjgy
1QKXax9jta7pUxTAuR4Yi7Ixn/1X7+8Sy5uTUSWMzacJXz+CKC4L6q/KvapVrUi6
kq7vdRUxfKV/VOoiIWXUXKGY6uEEUX5LXhS14DsJLInf8sAdSK0wai9iH7ON3XIP
ew2BSeQr6cUvWDlg4EZmRo8hGaHRM2YzhOk9Ve8BSlLlQL0rHJsoUD/noZkPWry4
ijMn3SXZ+F3/NIKDnxNhxIQUmFk0faJGkx9IlaW9BpIpLuYCVNK0sALJftdi8pW/
pzN0XcLVqJBdbYW6DnlBYhG0JeImI8DCzwR7HhUGafWRaaaQwxwp3dHrHbqj6Baw
vOda01o3qyRJFv2o9baKC8aF/RcJXcGz8xjzmmN95adUlgJoo7moJCCRLCc9VpsR
Dp8oDg57ZRsoBJ/ENWHfzft2sFDwMevIqUqqDlE5+U6ikO5/+B2Ip8UqdZg25chc
N4m8z5/vK9itjo5yzTkPRD6wwEWrAWrWYRZGeBgbug/aP3IxEL8Ma4pkPspOYqmC
SSVc3av/I5cVtxZZW+a4l4bA5Zmju/niwKDk/2px45ra42GYrMwzppPfpuYGAKBZ
IG3WrNFDLgYSkpiNyk0nxF/Oj+9AVTTPXKJLViqg/zJ2eZ0x1/P84gr6pZPeE37A
DdejGowuyDqmnVDOWvcq/1ISqT3cRpvMzbOzdj0mNU4Se0h8cuuhAvgSegP6+H+R
CNDo9jBYYExc5QhuanB9UcQ8dj0EGZzg4yM8uwUcdMfNGG52kXi1F8CVSlvmBCYc
Yn0YYUcG3kKjvmG005+SNUXv2d9fYyjDoZw+YyIoSJT7kuH+U34rETsTln2mPwNc
oO7Uj7rGkeEEQgHOeyG6PlJQ7f/44z+or/KVL0IR1fOOS7I4zlH90LQOT9Art9Od
632xfot0nd5KHVN3jw5lkt6SxfS2BrPh9HU3EszpWyY2pMcnwT86WeWB9bSC+wky
UuOWIA7mO7n6BLqwp5zrgUNovcyzOAy2VG5Ma7runLv9ymeqB6pk0FlWXk9oIE71
O2jDbsfzEEszpA4O7Ah3eqCV+8TeWLiOb+JjZnONpdKsaEi8JjsmqB0n6vLZ1gKH
BcRp00pvsBK4J/1RFizATC+aS00YkZnqRJsHhHPzbd5jZk4bmmW72nUSsoDYiigP
67CaxZpu94irXZ8MLuZCYBbtG00ortX74r774m4y+rY1Hf8T79NXICjNMAOXYONN
0EoVOh4MhayZnEkjzuro+xnaGx6Usr5CqJo+SmDuKwZA9J5eVzy+b7NNlsPZwg7p
DRzvA52JASl702ApVu5fKchfoR0dqIOd6N8XMuV4VWpJEoSoIk/qdt73Zz4msgpB
5mxC0cHKoRwXZmRJCO2+AOcG8XJiazLfdY1VG8+00028jumO3MRB8wdoVbMhBxr8
z2ktR/tUDRLLkR3GuQG9G2VaXspaKM8RwJNT+Jibe/UH/xRbFl9Jn4qgfl6z5yKu
4XyTG/SChx+n4wjTv5Cu+JRBtls0aA/FhKGofVz9TtnCvDLIqv5xmG+5F1xAR5xT
9m1Vry3kkDTRu5xtZJ6PEix0q43xgxPozpNC/OfIk7QhaW23VASX7c83LcvYqtXa
Vm+Q9l9Pgjk44n+27vCWY1/lAEnnvAklT9yHNB+b6HH3Bbc1opzjkWHgoBkYO+lm
IrVZcj+GZgUfAJ+E+SksUiMe9Z5VI73EJjaV8QdUKXDVYvdFh0Ts1VoA+Vr9c5u/
ZTF/GU1Ghero3oVDuJUSeYbTC+QBICbo6vX5V0hp1iPHFBfhGoR1W2U68uWBb+TS
vikO5lbVo7O71kdKaY7kK8O8c4LuRJ5/MVeGYhzFzfkRZhoELqMlMp3WLn9HKbPI
BX/13/k9F2O/YMHkqtxiwITfiMb5MQLkCiDZHjbcOzKNaKo5SRg4it/59BVXxhtD
BYx+PsxA+1tmib2bCidK5smtQoGi6YWC9SBi/MlFZ2tCKzjDRIW4G21M5bWPc6y5
2NXk4qsiJO/aWUww8cogiwfaworpLT5A3vCk05O8wj18CkfrjxAYhOrdP4tVZTJg
AuzXQ40dz3yPnZP+GU6L9BYL/HL0dyZbIhmo+YLkfsR0zj7fE0RL/aiNncj6BvV0
V1pYELkr3HAoT6hrd3o2EllyUwQtRofvGWpOuS0rAVqkWXTkWxPOzEf/bA/8/Kjs
vJ9YApw9FhV5MeBrvJIbE29/VEmag9V+pqmtXzhuLzehG/7EP7UNeAVPwrfYYsTA
1e4emezWN2kK6u2Wh4zJ0tP6b2gbdVsI+oUIjT7JrVF7DMC/r6jgxrEXPe+0nmXw
ggAtv86WUauFihwbWGXPoGXRXzjk7RRZlM8k15iTBQ4W2DoWXnZFmz9C9Lm1W7TR
w4UJYOPV9taYFrl4PAXu21ZXaraUfY4YgMyopn/M+UlpZiOVJSxlx0+xfs5UGmou
D3GR8kLL5thPW1lBHwQbPHgFrW0G/Iz3YwK1Lgjs/9V9sxmUx8+XsqaRvLJVk7Ku
DH74QbQtUwNFf0sIs0u7o8zZf8TbF/sZz6i5+HSPV5SSp0LuJS3gfdRwVEPQZFFl
FTxEO6ovewgaOVfMGMLL7xzRmhisRmG/sV97ulyZRWlCnjVuWvEfAp9SYC/4QiPp
NX0j/DExsHypqcZjBY0A/GcIfttrwbwy0Moo252Wq+WjbaocVBflVruUOnTKHfxm
3EhVfG65X8nEr1FO8uKLTbAWCrrUlMo6TbbaQkeO++kXrr9xWbSKpOadO84bWgb7
QPeRj3j/FISEy9V6Eai305aoEUmymLNhVd6tXoH/vCVQcm+VkcI5taV1x5i49nWj
IAAhxJQ4RfHBHrLG/3XXrc1M3YA8KADbJbbFOE+qOpPXqc5sVd2L4q/H/NuTODom
6+e+8eeKnONxnI9xQIUO74Gb+pYWgBGL3i9WAH+Pe8UXfIavnUImEhR6shk8LfkK
WkUTnsq/89lAbnfNRZbnS0LypbhK3Xi5LQkC4wcrqdIa5gNtCXLM/jwJm01wTsAU
UzfGJM6Tu4lvxtE5Xkyt7ahzAf+jPtWWljdAoUfAYelc2ycCMiE8mhzx/ZqzZW2X
0OYTsQeYtksebuEMN9hEhgv4oy+PGT7BT71jyC0HVewLZFrqpoVrf84X5YFx3zlM
2YESr3o1Cl6c5PbHlJGIgQOzc3lJ9Z/1H/Jdd/ELQ9yqQiDHDb0GkxPjYzswwCbh
wQl4j8Xywb6c2ND84iP8b94wiIV4zP9p4K+Z+qiA3eXhZ+sR6+YJo4ON9rtg+mLI
/hMHlZaXmf5EJ1vOxEM2Z4rDU1Z7I5nK1BBzxenEiBYeh6Syjws6Aa3ktDhtIwwP
bJcH8/mDZ7PG8JnVLUwPOfNXuql4hkgtisekbba7QjCIFo4r/+gOf2zyoz7e3l0S
sPe+3O+w/GvgZ7tPQMPNqjBgicQoy78N+i1t+7+Ain/F1SM4HPDgNfMIrMcBdeOG
XqaUDSZPApGaSoJNnW14H25FMDFuQz7m+eQ8VeuAtq2GcGG5Mo6mIIlprceSniNT
XAV94d/PyV6ztoYQyMawruA0nLxju5c6X9/c4HB8TLljM7TdmkDnyTQZx7W3G8vB
k7zpX19EeQQIRoaePOih0p1geSu2gLtGjchimAZrvYq0DVFi9nLfv6XLd6ovNS2v
HpzOOiInfzgSDvQeM/wLn5sHMn7eGYNe0Zd/cyJg4gerIIWA4Cunf9yq9CbUdlv+
lsNJ/68jKnGebX5AZjjEOM8Lfz+vqzWECZF0PTZF7DtCAKIAW0wWENoPQO2tpJIe
DdMMGA1NyJACj6GR3UaGpiZCxWwDnWtpeuPsoMIfUbtiDo/HHVUexpV3981aWHJG
VFLjiKKTHkV0Aj7nlhDrj7mj/7zWx79kFiVK+Ow8TDrhq7ZczRIDDpWzkBabLzt9
v3UHSwTOi15qNkoy7xTnrU27DBKcn/60ranluAeeW+IBvzSwpXbenVwF3chZeDBY
jqAaye7fyJhheJtQspGWGcSyp4i4zKnhJY5LHaS0bSWxOVDSDlOqr8nfOxyzbGeG
KE19ItyCB7y1wqaAeITaX1XQsqnrAxfC0etmvaFGXKF4qJaWCQQ+46PxKiGq3f6L
u9Hn+s7VFrj1/C4Tjr/+WG0XsEZz3qNs01NnIoZdohDkEfRM+daQ+qxybrMXBb8+
ePLcMyP6g/tAv41fnWYHL2OcomrUGXcRC018C9Tzz9pZ0PFfGrDVVSaW4lHA1Mh4
69Z87DwKEsmoeUJMl4RUYtzNxLs2idv8sp2OwN3TskFx1kMK6CMk9ZAtw0bN6r5X
5pAVtF9s1k0ViMJo00SPREMMnGc5rdpmK92rBHbU7qr2xqQIFOsmZsEtc+NJ8glC
7/y++qKI2oja8Fkux9g+/FOuwoJmJ9ETWIP98dL2ClTsGAx0+kUKevErr+l+68/f
jRa4bP2h/4QBXmDH/deQyU9caJYOtSxvK5cmKRLq/eh6EyC4+WF6J6lipuFJwaSN
+oWBgkwxK1nQJ+k2s/tEreQowDUTR2+s9kdWFFsfulXgl5pIGzOxi2lwSlLwQE2a
thD+ZJ22NcdLSVJoIiuyDslZL19KFJJIQWJtcTjVyrgunKb3XvPxNS8HczzPNN3z
XQj5wAz/ddNZMU1h3Sr09oPGcpVxWbIk/ryHGmIHuW+XFQnlzt1vXEZkoQ2wgsJD
S/ArxM/dAGHMqHqcar0gzuNckp3r+hziUYf2vfXuBLcnBGTrxLzTxoCzifkkrgZB
S6MvBW45659vNs2Hmv0iHgQs7fYHa9ax64uGdJLlcq9xx+3abW8+aPi55cT5338b
wrvuTjyh9jeXfSHy6zPYjQCrQyLPB4RlxsgAKZ0h+OS4Qd4uHbrgIHqtbYHP0oBt
WHJLIi2Lc9HQp9Xd/VFiSe1kAoBhOQ5sHVi4349N3PWItq/2z98dWvjzLEJn4O5m
iSFys1I20hKRhbmB5dVGzqVuN6Jl3xA9lWBUtAHN17C+L4/FyqaYtXMHAc1Mm92y
5VreO4Hi49bojgn2xpWTNrYHI85vBYpK46QfDfADOYV1+moLOpT9zEUD//0pB1bg
qXPlFdYYXm29qe1jf+K/4bPf0Xzg+F7qOg9yD/UGoflSf3OvvxtFaQPpBWlD2HNs
PiADcnkvXRlAWpSbJz4aE1RziiGdzcCbQWFXw0aL7g9Y0vMZ0fImNXx22XS1Ex2x
Q3C9ujqK6x4KOgnbBIKjEILDBbNqIUGgjH9MJsDhIWjJa3aaTBQR5QaljgNOiaTb
XFSOSAhgNigxFXxUCfgVC1AesL3CbuU/ILftO33oHySIY1ftoXWjjzCAV8z/o+5U
mHeygg3mrCCagsQXO4wKJTJDTYAvKFuBDkZ4872iSJWuqOIAu0zAvHoSQ+9M1Ow8
xubnKlpd3b8dd+V/c83q6NaiKSMXuhWmX0RqMFKXloj2YlnXPysoxgO6S5jHQLLa
+KjqsCxmdS92qiCmfZ3GLppPfaet5GYM7kRIK96lSb68T0uWdAJGUSc4r2Tt9EDr
JYYnesbh1ckOVJ5KadOQdJn+BN1ZZUe3buPdlJaCgAOgdsAHoEoz0q1JTT4+tHkU
9zqzBzHtA0Zrj3rC/+dU2cvGOmKyvUlgQrvf2cZaOchN4yuJj9cLBvgtYxx2LxQO
U4mh/bPVYpkbdwhomKMMy1QqO5YwidD/KQgLfrjT0CITXCfNiaVmUsG3p5Q0JzOw
fr2GY1Amh57l7cbuC2Y2AYmwaKFZ2yizoZTVtMNI57cxVeOGGd76pWgPGFuOv8HJ
LLTHIsPzw89Vu7HoZotL7gmnwUhV8HpvF63NsBPvZFwSawLnvWa/3aa+jRM4pov9
6tpP4R+uIrikIMXF3jd8lEOiD/RDy2ZFVcsq1g7KSfmKPP0VyvqJGd/2RgyYggXy
Up/Y/K3XRxaxtDab+vm3tBwrCefSaADUWrdKNIQjEBqe7juGd4fN41RDIwy1hx9d
J7xFDd5kA+76E4YGEGRSWq3jfTCIyNorvz2pW2fG3N41jnoI/SubzXTERg2u10pO
3RHLvXR2FXvx17MhndVDt7ycBcNEtlaYrRRoaIHtTsMamBwtjLPvvX3uDMP1nsRT
nI19iXclvTOMa/cm0V21/52oeqD3z+JZhjfi3JbIAxGnD0Uc9/OMyhWbAMwb+6H2
fZ6MtVUEvwZYs4dWLRRo34nZTCHZipbHyRq9BA9Y4saavf+HvhBHe4yJ3yb6tRW/
BHHNt8z1bfjz3bjo1LBR0yCRB0TLKpbzWU3mPpgwsTYOx+8fDoP00oaUbKzhifMq
sZGGIPpmnduWLVcoJ4MdhEeZ7cmv5PjM7WZ2wMhrsANzumX5baQcDbdJEgQHw22E
4pkeuTgpaXn+KtB/mR0mQIqH8mKwdRMyzhNOLGkB6J3Na/4w24gCsncK3elTx8sZ
sQdqvu8jRFraGFxJ7meT2i7Qgp0nE7KgSktxrFM0biaizdsEtfB/Fkpjnoz8T6J4
Ek2x7XiRucm+CjUS1JtCynHQeSYrgxRh1p0BJE50Alv5RWjvvvuiGQEuuE7Yuu1a
Xv3eWmTDPgwxv5llAPgjNQGfArnNiSw+qccmlICpRNttP4G73q4Khs3hPHCH2Erv
XqzCYtl4MzcW7N3J4eiO1HqfZpzglpkU3/7n6oqxOSy75q9zaCp6OFaPby/a+KMW
dVkIFfy8KSHadQsEXYAnVNEIX8TmCIA0pCAsbCPYw3a+koj0URaccU+GR+OsJ5AM
T6dkahIehotX4BahcxCVGpswgPjG96RymhluoqS+khvMdMo6g0380MaLaEuiUIo1
eYaZ5BeOd5zaajOxBDirABR3lYtZxP2ZHSCTxPyGpXfnuDAKAGiPTAXdCF3IH57A
mw8nvd0Hivny383OrmWJHXUSbSAa0+Ckgoj9VcAXYcjmeqSJ0BgaZyoFm6gdLu3E
Eob86+kAkgsCdJIs8turRu9DBhVnkV/aKAg8GaDxjQNm4Cf5Rh42MmAGrFJf4CD/
YDm/g2N0RbXD0OXMVk57FmaOS5IXLF3UjteEXBS6mmqprXZpZ/kZMnjDhMkjUYo+
wKdQlRwvVwwQll4UNlc/T0Um372Gr3dC5UROD+5cX6vUnZ2OEOZx9Hjil6nw+l2F
HsNMkqMFXBT9b+DQHR4XFHIiwEQg+VcgLwR/FPU8l8pYTUtcCVJh+VQdM92BvVy0
8XA7H03onqTkjXg5/g0+gA==
`protect end_protected