`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 11776 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/9huKRhRMtvnNqb3Z+UU7TahEoHV+T8U3P3ufru7l1O
3DlgtZzb9QxCbOjthp9+wDkjygH0eUfDrEl1ovhZG639kMeIEY06ujE6KZGFJxsF
MMPUP6DCb+Oue9kPpaU+Xy9sA+2JdNHnLPOwnCTBa0kUfoqlkphn57kirctNt2i5
bHx5S2nt+fV1gK2il8jAzAZVINmNJDPe4GhnIY+CVFA+EVy3n3wMBzWi7QwXlXQN
J9ZJCU4U/hQIvf6AlS1OtX6eiKEo55y3kqbFOo0XjmUFZF5JcRsFppnvMv2Ja/BZ
CAgtUTZvmh53je0HWkuR12RBlgCP2NwqLohyWFCRZo9qyO2J0r3d9SzTqZ0GT863
sM1O1eisMH5MnAiuazJRfZMIEfV+cSmCN7qEmbx6FYxoYNM976Jke6YX4Xf4PB0v
vFzX4jHpGi1Pi4g+NsQ/VY7XUlKRjaMBU3H02vP0q08rdGkial/snhaSzzXi6FyI
Wv9ZNwrObWatmfIQF0SRu4iz0txoDBrsLCyXPwl6irTiO411CpQKghI3b/fy5bmV
9ApuaohQsQw00ruqlPy9dLCny+TpSgc+AH72OMClsontNx+2+xLQ/i1LpmnKz8JB
UDuAD2Ztf08fKWUr6SctMPKWNNmOf4FEcdsrmnOrmDqwifdDWdbR/M1er7zszuL2
wuXYT5AZ4u6+NoNQK/ehfvWcX7I/jG3b8sIdDeI1gSWrcSlMPEXQHFiE9/XGf2Tv
Pw55eEVPqZb+C4pzgIBR23esTUKe+nrxB/WrCSHgv05T67VvBCaZDQpB6rz+Ktd/
3WdUh0EjEhcoF0rhkE0Dsnm1woXMkUTJNTRE7utMEgslcoPyWlk7uPx3sbloxsrs
500AsBlNPrMh/0WPasCAwPaGwAVbCgEDYQq1bvghJ653wtH1jrs2dBBYFROrsub7
1uWapBrUhHW+KcbYZBKmFnoOdjyzSer8aFWu57Ja+/i/3tJ7eyy2nvk3VHOuE+PW
K5ZgLcf1nEq28dup6YsJCFJp1rFqr7jDDjaWWdvG3Uiy1sbsBbbiJ8WnE1xvBAMX
HgPa4sdZ57SaYYHDIFL0rfzf/DeM18mcWCeERhjTGWddAWgaMuIMJQtaE7Nmbu95
/D8yUXdm+/TqE8Mh0Hj2ibw0lwhMUiz9Rz/5xOVTBdng8FufOR9qc6qHg50ROkqr
fzsTjAF7H9tyHmArvUi2+ED/nbOHNVv2/wTWpgtbdKyF6qKMsSnH5XMzXFF3EC8Y
Vn9quQ4zXWaDbor9thS80oUMguY6iuoMcWyC5osVijG5oH3BIkJeBa8UfYccTiT5
QQfoBB5GYVAG81XdpFSEltY4rbcYi2N5Ni6AjIC07Mbh+vhAKpsd29bUHjaY04I+
/BHg3mp35v/5s1jWuiYj2eKWd2TXO6YbJS5GhakHSUV13WZCKD2HAnSeCvSITM3Q
lw3cUimKTopK+T1b/gnQt8XrfB5FQ4D6YPDfLS8vAyAOQq+pXaK3ZjPzsr42D9Xk
o42HBrzpaNwqgSkZxIUW7TN7XLyv3hbnh43sX7bLliwhuis3o8X8TJqF3vtrEmMK
OkSOZ2QnFgQ25FrChJLs46pEszKDLC0kiTcZZlgjOI5BkchnFxV1obzhuNfLVFt9
HuRzPDjrtGByYVtnITYJ3ql7+rJ9vIPcWetoMK64BVQ7GmqR8zbC9wFt7TsbrXqx
SI9ODI+szAZw9sYPQ9A8/muG0oWBCF1MpFIVbPj0z4+NjMiGmpMXo//CfKJuCyy8
s/+Pfdm5H0HAqyZAyMS4Nyw6OG8fbrSaEPdaVMeGviS9BkxP2fNKxl2G2c5LL1KV
rLehuYGx3/yhdb0NghMbGq8a/VSDJYoUy7UGaWoUYDMNFdytFHsz1KV2OPieE91t
n37H6R9v9yigh3/B1GyriK/qqNgyGTYxjbyYrjbBLTigHruwL+BKuIGwMC43wxt4
lkwoXWMLiV2ofNwsTqPmtJ9TK/xZWk9ESFKFb/fVS1MgyT8jNtmJjDl5lq5BHwe7
w5TWjWvuz7aIhi736dZijZtfJ8BVc2Aa+4TQCrDqSIk/I2JeVWY3dWXeI0iYPAh1
seYFbGScx/Y1FE1JSO66LHYt7GnTs2ZCfCHjd7R4yv6tsKqCT8ocM2pLps9KMk6R
SE+WJu7Q7d+vWOnnII2MzqGYSIassVkrDhWJ9HGXLq/4TOGuTW2zoWirIslRh+to
887nPK37rX48gQPCFsOxARNthSKZUBJPcrC5JpFwSgfUnZ5XyS2tEcCduugatneR
KJUUypF1oAFqd51sHckLgrgvZVAy5g2P4L/N0F+DSO95NYpbPsT0r+Y7PtYPDrQu
8IVSTDrEVEJFkDqVpk8ec4eqspW3mOXXXQ5P6zpCbqWrjTuyvUs0z7QnWdsrxGbK
OZCDGDadvmVCx9twjXmG7x3PxrjaYzYjnICdbEfCd7pbz40G6vZflUO/4Je1sXu1
WIxcH79rV2doNjRBTYsfchL1AwhuRM248gFFgS2fZaRc6Ift/O5qlAAvHnXPmOOV
CGKxyhw+1KoWcGqH0y8E/seeWBR1/R2wscpIHZOxzEmM1nPWo8h/vjZuwyt02xkR
1d7uZRLFNV0Lb/8KbdOBiqhMOfyXiP1GwB9Fv3QXoLLH+PA6EElz7Ih3uWlFTR0S
HkLehcm2zea9ja4wSVdu7tAAFQ7EmzUSI7Yq9dJwJ8oKixiXAzHjnFgyj8u2BjQq
Lv8y36V1EU84/WHDzB9AzNqjCHGQjwJ3+EurJ3GbCeLX+dqJIEnSa6JDC6uqlw9p
XGyw39LDNhl4qnbP4af8RQWRdtLaysBZA8jjLKW015h3Q1x9aKztufwpV+KlfiKQ
SyKjezJnxf9l8AX3/+/cF/POlHvUaiJa5/2aaNowQiU0ynl+lqeLWsAOcFrbnn2N
UxhBXYSNrkvGldiu2SQvwPFrqY8DKZrEREBc8LokXew56b4hpL0JxjWJGMZvc9/G
RtHbKUq0OfrA3200/JyWqzzFN/dKyOc1y/+11x8n3f9uKvtqKsvdsxVDy/5nFoDq
KQBzk2pt+fCA9Xd8zdJSY9WT2jbDlR5qwIHjrUdAvcCE6apBicQTxkM7NwRucMJc
/GlVSz4RXzCl82lIsc5EQLbLi/Hv7Nh+9QxKaceJ+sT8RR48V+Ge3hL2WHI12R0I
CNOY9upLezIOzQKgY4Jk66IIn5MxcEUKdjLOMZ80lVxzj6WRKL9LDot5FRBDHZLc
w5KoCpPvD4tEVmmvUw43q019vyXeeSeQKTYDKfd+tt+sb3M7DocQgfpxR4QJ/Nwz
701Dj6drJtz+g4BrtTsbJSeCVrFx+uVQ5868A5mIkcKuiQS8xUycutzMJ67CqOKg
nDmjQODSMW4TpJ0QFUTclGvn+DVPIToHAvi1Te3uVvoCHTIjmY5e2qIJi+Ya0sl2
TaGpNVfO4/HyxmOTRTDbjf7wtcq3gDQkYRt1TzRiZ7AFzKsd8zV3mnFvnAET2JN5
NDNSAHi0zl6mg8T2jNyvyxQy9/EVHFGHUzg4rWJbV58C4/SW6Sw0UgwhfcmosVSE
Cm8RM/c9XPL8Mb7wcVWjjaxsJfbuetO49+gcvJv5GEry9Ls4kBVr1Qx1koCPn6uV
SEsIsAapjgJrfijV/bXYM1WRI7Ep5mctocp55+0tZf5W1foWKy45dl6dQFsL/1QV
S7SJ+RtZSTO/mQgICe2IFYLd7LdJIgilnH5P0UFNGklj/w+EwicU3NJU+cfOWQo/
miXef+FvS/9aUPVwesQkGpWzqtDO4KrE4U4VWIbTxGSbHiXIbFdy5DEfT7NpTHMZ
HksAjyYe4rqH+7eFohNFMellxwIEX6k3SGEB0r74rXUEdcPgE8jK82smJEDOzVh+
ajiWO98fVE9WPtNQJOeKkrMEULIOUeu0QFhVqfOVowdWBymgj/Lr+Cj3tXvrwnUW
dglnjMDIpFOERpMpZ4/w81wzXmWza1+DQ7V8gOCpngLRMQPYFfkRVtu7bg81/lvG
WV1rRr5wsq4u6SwmmXwNhIJf4AQwvZqyRAsA1MpwWBQyUZbedmEHKA9ngK6vfgXX
EjJWMvUqCx2WpW9Ff1ZgNEJ6xt1KBfKjygyjqtTD8OYkdd8lIv4fhoY9andMMdY+
vfAIn2ywD1+nPQWWAi/vkY8RAVQ44M13uSv+pGRRGRT3sqOiVVI3yxJa6H2JBH7p
r/b5OHfUrwEmf8x6cfR0e91el4kahscncxeyxz5LEQjdwvPyhYI6vF2ipBHCbEyy
kvASzSkDifu7SDeH9LhH39gx3beoTrtjVI1CA26rCE/Ac7+NnMHeNKEQ3lNN1vL3
dxl359/9fqxPRrp7hlLpBx4OWEK/WTvJbpcjYwmlaFRXye+2eEwBaYBchQxdXagg
IW0fLD70qsJwlPo64c9E8uxQlh5WPuAtjAXf+wLSHL2aDU32w1BA9div3t/5Jwr6
LurpKiYfKo5MtsjnN0b3VEr/VDwVd2jsdo+g7JL4IKAV1m2VJ0GvuOKbG0QwBTkG
6fo0Iy5TWp2EyX1ZXLo869Pvkk61C+2+IXodh6/x3d/9mKl3WvksbAcG+lenmNWP
Xy9Q0iLcN7CATmW7PoHQZGW/GLFqYO1YZax3XkdAkyBXs48w04aPklJaQl+VFPV8
aeU8q1+KkbvQ24cuxuv7SmGr8pF8Tt9dOnsMBfvkmwEjXW2GnULx/v1vSTOZkOWn
OVJ7Qh18Csnh4xj+XAM8/DdAhP09Meq1wcRNhP8j0MRuWXuF833fYv3lhAhd1kzB
nGWCqGkCMr47P0GAeN9wUeePsc8JwJaOUwfpm2LBAYXwA00NXZo8+XjtFMP5w1d/
DtvnBd+YGIqoxethDfASdOgnD6j+r2QAkNfamjMmdDXiG5zZpWnYFqT/nHYr6m5P
ves92PYgMTVv/YN4h8g0MFGYxb+sWC+1PhECxCXUgN2Fiwqrf/BwbDOf+Qp32UgB
t8S1L3WCG5zKeM6QFDyRZZ1BKMlmvewNfzNivwIxtAj4FdR9mDldLE8RZvC6z+c0
+KIF274tMB/SI5dFW2B7fKaf3Xk4t9CxsrDh6FY95MoZ/TpfEg9oChZVDGGiaWRN
VJLI5XyQEbeuGudZtScte1catc69wmasBZvgfnSVSzN+8PS0UZYzZuaGnSDdyPLJ
xCmLv+DIA3SN+GA/qrs+kmhvVvHeSnMctka5LnoOPmebCBxu4uCqvbZKt7J8jdLX
83OAvdM296iELsCz1mNQkFRkDuixpzANMuf9DFHI5owGP/MJ6IPy9KptG71npiHp
fy9RrKcEh215tqW0a1J5S9Tt41eCSqOR6FVWwhLX0dkwvvGrJss/+mTjI5aeWUM/
7vde9h9eK+QpOrK03OQkRaDJc1AuapujGKSG7Tz9lcd6PtBx2Snt2xRsNE01m6oR
tz/kgsv/cCFaD807fQFyAnxo2jQ3aU6hhZbD+VFe0N184tIfxGHvtt8sgzg9j2j7
enoRFe8D61BeuSlIVmwmm7E+EzAqO9g7Je+ykcYiSROtzqYAjFd3o/IH6IL+9b7B
CQqrv7g8vMKyz0+BpFfxv5y07OCOidNThxaQXBdr4+CPQ8HUCzTjG4fcQ9FpmThB
s3FPT6gQTwc6v3SG3unB5KLcarr64b7LiMvW5eppdEEGmLI/R9b1GSRUHJ3fsJss
BWArKqY09emzI6YRs/26y3O6OQX73Vj0PCO/g6p7zmk2ecH9URNSQILBpertA74v
HJypL8rr8xq5fuc0q4jGVFq2cFNKGCRqt4bffwRFovDTudN3Dv1WTuVNTkBZcbu3
xFycVYTCsBc75UvOIVgRSPS4ru07HAiU7R0K7yNkCfEROcRfoFF3aBOYTaGuD6VO
xwKMdp81JS3N+rbxhoCaTkus3umeTfcy0Y5gXma6lp9b9M8k2TumClQWZWQe4wBE
fubPdSVcG6yIJ8njNZKN/JiUrnONo5WP14TJozXRpF+9/uj9/qslbvGzZwjfN3Hy
6Bg/VXHAnsdAz8r9zFp+cTr+lDsPEEma/OyNq1Y+ToNu4aEE9uN/+PmU5QoA/k4K
czIItETD31vRJEskek+tNv80cov2h5vOqSNFINum/3RT5tLItdh8xzp7bdc9yotO
r7Dr48R16zlcc4WP9USa2ACH4dBiBFSB1AuGYTFYE1oQky+3yx1CQrRMaG9XC966
ISu7gSB3NnYEegGl2xHkgv0rGIG69Cwr/3g91Oq4KJQfNGUtj8UJEDFLGioTdFJe
u1rniNRzUJm7zPZdV2ig1BqK9pFuyyUnffsl8Zzz/CTg6plrH/LBz4MWBe0UtbUR
2/PAPhbqNwJ3gGaoMptawPpMjqqFoBUESZ/UPpjFIN3O9rXoqlhKX3u4IFxSDxES
RsuHV08tALsXTvRou05Cib2GwjiJco/L2MmI557OcH9uv7pVOzQ9ikKY+Zions59
cJEme5U0U/I+u8hyZU572NzYSLefQ8oGZfg0GWDm3LSSpcVfvCOpcn6/8SrM+if3
njwVHxsYnF75hjr3vjhU3E1j6C/YZ5pDiSHZo+vgrajG2Rxyl+MoXgo1Xsddsvir
ttMouu6S0qRpL5LugroYyDZ/hea+2utzCj6xEHonlsLu5Dux+23PTn/Ikc3yIAKH
+SuTd8h+0NTkUyhmY+jIiPSlXTK1cfphWrIj5fKHROeN/fQF0qb3PXOUZCpUVHjY
rfyQGXpAQ+Y3m5oweseWNojYG2m/siKMLFxc2k4rYa22EArBU72aKf0SBwbraont
BJuv8UsCbHLLnG8PQ8CDXgpOZ5KNFWeap9g+4iPJs/Zl9pBCLYQzaY80toxQdl0n
2HyvobX9WnWbum31ecSEHRwkygEpTAd0529oSjIyTHkd88/dz3J5T+oXVkrk+lJw
vnsR6y49Sl5qgLuP5J5h7QuAnmPl8I57T6Hdo6EFG1lU5vBGPCaFU1GbZd1NTHVF
nb9ukqKF3on7xyqWlKuDzNVTtHU1LZt2CduNXZ7CWERvHUZKE/i41XmdW4ZcDwoW
UxIdrrk+QK1PF3Ze5tFP06PWt4SHHfbt+lfi86GEcJimBLwwt8bwUOJ9Ca5mX4Ef
zhA8L5vjJMIzDpla2tTow2q42p7km7I3UEVb1V7vYymMmwmepbt/xZo+K7TV1eTT
B0DBA+oMvwP5gIqCSCCwiwfJr9OLL2pEIyuz6BWR+mUqqEsUD87WjMfObVcYjJ3j
4K3XtD9PhDFYJ3Mc1L2XBVzBjiXAuLHcedlW+Mu2dyYUDabafI9iv/vgb+028vtl
RMTJnNnU/e0DpyNYJOC410NIJeqCtEtJtm1oTMz/J7m5sBpsIZvMj3IgOL7uKsWQ
Wstt8smqfDgzMuXEFNbT0vRAmcVSg3QiYEngXPmbfEFmUBYorhUIHEDmoe2IlWeQ
9eB4Kz+9SEOeIaj7LScScZ0h+x8UKvH2D/obr8U0HRwIEYRHw+iaxCIQXTD3sONE
YOlz8g+pswqBbJPor8ZbaJffp4U1jc5OR9GbETwesM9zEbaE5h+QrU1zqEXU+0xu
NdCQT5cupmvnurlZKLNg8+2xK/1NIUE3oL6P08hn+o6NnpQkTAWpgXUzUzV2QcxO
dYQmE4OznH7SfULbg6iSD1HCoWIyFjppzNuIlDE3Hx1O3kAKJh6OY+1xRsxW5tM0
INvlV2K8vK70c7SRwvhAWx5BQc7JYkC/IMIu5UyOsMarzri/qGsginvVjSEeZYiB
orgZ0ZXqAkZ6RlNN1gMfz3poxtUmH2quj+a8H69B2dX0Pxb4VQOstfIEIUpjMvof
XwoX/0SFlNkCTQ4gr2lFiLvTwrY2LH2j5+DQQouf2bKXxuYawtQGY4QSnDc47Zic
mmGp6c4fMo+sUwD96oloPVPzqaErjGt/CjcFHg0xBgImDNP8ywFMjogaamcxDerR
Poe7W/O8TCd6h9QwbmfWC//ECsUcrpgN6AFioKWtgK7pYiiubTSX3KK0qETaUFpT
wNH25WTk0O02+M9aMBMywqPRrvMFd3lvUHhaqnZbfuka2ZpTodUKBeJ5L/B16NDu
9BheGIkL6MSwZ48wXTN1IT1fh3ltyCjRbGX7L2fL88UELuMsXRqp6Ini5t9jfH1g
+CVEPaGGOn6uBCNHJtKLwcqs0HYEXgNx3GTG/GkHAmD9VUCkdPiCUxPSRZA1AIsX
5mKza+2MUEOPcVjwl7J8wrfmfE177X+3vzhfb6jAqJ28zBobJuce5Mz7fhwpQWWd
EJvC0HXPeWC7GsogfzwqYQ5vFzsNYp/qjusvsDVowWs3UTH2/iHl0If1yA0pCu2B
KMrtN0u9za30ydck3wlC2ysxgdXCL4pTu82WPTDyM8Ww6gOvDuZCvz5xQvnw6sX8
DTgfKxRpHRXhhSL/O0PgV73/pXU0+JTqMawpGFUNYpDW5KxC2RYz1OHAItkQ1r+4
HckLPmA1vtRuEs8vHfNTO4T5ekbPkJaLv32oA/22371qj9kyR9cPy9a//r9kvTfY
8jgOKaNbP1Ivxb4Ry1qvruKs22pLV6Fj3NK+1V7M4EykbeDQrZinsVFL+AZI3UQS
A+thJEAd5XzLn09ii9+udDIpzxrIGmYrii5XcXk3PMZ3Ky72UQl+cZZk1ihtuq03
BPiNIXsdIsnRfO7BiTfLyPhIYiEReqRBJ9mraprFard0PyJhG2n9+7Xq0dFFtUeH
Hk4C1pAgz6liuFdbN6vFBatDHiF0X3l1pXriYp9Bee5LI0NGUmF9kWJ5Ev6n89Bp
cIKivLA1ZoDINY6lkxwyz2QzVjVfSKAmNEiXRx4ZCLU27Q3oIQFoG7YqlWE7W9AR
vDWV/HKCFD36qhFE50kN9SU86Z7LQiW2S2EziLrShVDOBtLaMgUwHTdlhtC2SgSx
RXQeRxM0Na2nb9MeDQ951Juzxcv1ZFuNbxWfM+QMuESUM61rVvozQ+3+JMOKQI2J
1hlppZo7dfdQnyM9agMLcCFHww5R0fCaw+e5Hh7mdIzmBmPx66uGgl1u5u1wcDBO
koo5zuPANBB4SKBa/WmSNBEB+ecCcF7+Xm/h1OOrGtQ8hKFTVc5hI1AlobKRZKDH
A++ogPmm8C/7ZGyZS0c9h3W1HRrMZ2fQcl4i1tGR6cKM8bJyPm5h1noOvaG4SnSq
Pq7iSwU4ey+w0f3nHJKYVk/ROuQiWgboeyyMbA42UkHIhiGls7tBSigCOIe11Odo
Fhi8Ctn0PlSYsfTq8fwQy1G7/SFMuccJZ/go2xkKvJkMyfLOavbtC3n/Ijh4E00C
Fl5UfXAlSACakHFfZLdANwtD3Wpzl1Td9959FbL406g13RTed28/mnGp4kMtBn6o
a45fmG0oT74huyGfRfHWlNPGU8mVIdfxgQGk3fVZ2o+t3A00U9/fhUQy8xqc0pYm
IbMxHYJ87LAg7OC1UE3L3eQxFKfkmbdUvNlTDaHm95uYBVnYX2EF/T5iG8j61CIj
9uhzHS1VisqzlyIZlIezLEBJKyT4P5yVS/hib0I8gZq/aH02GBW07EhUDGFIGlyU
uWG7pYOSxJKOrxASwj4qPI60Ccn4rnyCY5GPajDvRBH4HJ4nYI4Rw1HdoM58nklI
Oqi+gYdJS5B2CTG6H08TgdbM1TxuJhj4IY2IAPrZ/zLODZrTg7VxgZadaq83Rj93
ZE3vTk7wqI1mj2KZ7cyF6pcSXTDroNnkjduOiWIm8mTILstozXbjeNwIo3154/nZ
tOafQ6LKnGvPkVHkrgcP6fzW0O3CTHGyEZlXLykmuiIepI3JQxd7/nn/HdkFWPyj
x/vjbf0zvRx4l3CMR6JCAufrpnoKd5f3NFJSfUbZpMhKCPmZDmNIlqoXf1YF7HVI
K3D2o5IkTNjab8l5I6z/fxaCWTClmSLNO/Vzf6eXfNDS0eJyrFBS3qw4DSBjLCBg
sEuFo2zMZYhiCQKNz3Q0pADW0i5ox9+hav8FYAV5N/SSzWegqoBmFmj/ChDPKa/d
hqU646lI8FfpR5jnjICMoSQLMmaqMp4wiScOJj9EOf0r4QmQ56nDsGi2b1BsDEM+
KMxXDND1JmK4tfbV9NBvfmf9FkdSIddPhN8O3KK3rX4ddkjWtuqyTljSgj44oewR
qIurwx7IXJ54EX9UN6Cb9R2FqHovZaL0zCBMQLce8adwcO32SaijaPzrIHYDFHga
KIvZEHyg6aQe3sv2Kt2MceD2qiss94vF8DaZQFhWGNliivWW9WkFPoiziqxNUj4P
IwHLL/no3MhqWAPYMhSJHZWfqg+8r/elwpTCROtOPmx0Vp/uB8/6/yXBuOOfneot
/JhfSmGpJ6d7NYnoHA/6l0x2OeObIJymfhNdBYFzmdpACm95QaBop5UTbKmDuhi9
p2AmLz560M/7B6Ktd1yYyVtKxzQY8bD1p79iCgQSF4qBEmhvLl8K5kbqTwU6vELH
D5FrZv6WaYIsbSbzMqRBy5z1DVdE9U/Lr5aJrsfnoKsn1Do0dfN/XFXzmEDjTubm
pYplL9CcZ+mkWZpetLxbqgB3JhRhbmmcNGXxZjmbt0djo5E7OUsl0lOBWStld5pN
kBPDS7WstLMDmj1F0NhKwecP4h9eyJPEfykzFXnvPIyJq8V+ohuagmtWKfQQrR6v
5Mt5ytoD9tmrHZCMx5lAdoPEq4CvfvzSIwyuvVT3v9wvCeeTcx1JSHqPn95GqFuN
bXRO++rbdbxAp7phPjHTUe+kp0OKtnySPBm3dMWr3hOZj89fGg3z9U2pFrPkEepM
yf0Z0bH9Dp6vvUNapxBD+Po2W4UFAIh6sAUOyLBbmfK+VRzkYq/FoXt49VnBiz4s
B8U0UplmisSetUAFKsl/ybNvkmbS2f6GluuxhY8/SzaZKAC0mtl+ssa2bKTOBG5/
Wy9ZSs75kdcLfvtb/DgxegzFHtyKFO56YvqnpwmU9FTTgMClOHDxEW/2+sE1VoU6
w4a9d9nzL2Kbprpc36NAdbKuqFZIWOS5jQamMl01osQQeStrZLDTZrLpstxilFi0
3GcWm+0cA0/KJP20DBMlmce/UrhfM789BH0L7Db7JZBNsieKdQlcNh7aDt8vR8dO
7cTljsA3Dxpe33WFlY/cAwxXAb4+yee+1OZmtW5UxYKP1b2lMPaBMdMjJyCKW3Uc
PlioZfweznR8Xs+GN8Jc8ehZorS+uLHAPhz2Ft5rUiGHHUswNI58SpEvGlzM7LvQ
1jpjtG1R/oYYPEC09xasKSiXJIdv+iSXeiPAe7rdurMyyPjAmpXqDi/3iHjz/d10
A0OqUWhkVRKmjt+kDNbQW9o4Uemx5PKei/sNo+wLS37U0C3Q83cmg0KuyfA0VOT/
hGZCO6OGSUziBDxJDcNT0p6VuW2Fy9YQbiePPZmxB0LkBabN2gjtlctrhLmb0ckT
l44qnJSoZTp0uHv5N8QTcqM2RE44Pot6y1Ay8RO4mqsZ0AQlonbZGu9f+R9tqp8W
a7jCu/ZLS4uQLvTfWnh9VcZGxzPD1XL8M//b98IAVssNTpEKV9SLNjUFPeJvTQza
OnnDm84ksGhKbQQPZZHx8YLZqpFlmr2YP/2Vf290PShplZfp5S2IqDBWDaX+GyVQ
y+gzYcPXGDqgSP2oend1k9yzGUV+M1WKUXyCOBousqGTLzgnTpIUABqJ+Uzdlf9V
dk5HDPSdxjIIVQkMmZ/HshlCvFGuaeJugXX2xSQMZU/kjb4bMPqsCJ+LEdFQxUIP
KdyFxzT267ZJmfyZDmXP+L6lZy/Nw9UxoF/b+g9I3r8F3ab01D2e19QvVYop1Ijs
WNwCoFw1SfLHPUDahrKrFqbm1/kgEir9ABQYK3/gvD3WlHLEdpMT2st8uD89VF8W
uAwEW9JRp/Wji1fX+TaSFnJ1JE1sikQfSlnAY5rsl1WqKpUQ21hrMqEN3Tfzx31I
HoZfqe3rOD+ecpIrGtnplu179mAmxJ54dM7pmll0C29EqU5uoSkqZ7wJ5VhI6As4
1zreLcyHlS1DGhfzVEleSBCF83JUOs9f5Y/i/Y2nYTAJNy9dNtSz3FJJCQSA5oGb
RAsTRFssu3oAwq0fmLspWdmpQ+x3UzVkO11PSzYTfztpKDRXDyknEBXAn9gbq+l4
b92sUO/VIK4JKWxbp2rYNbHZIB62nWLXHAEb5uhWXpKc0qZ8zGGhQQzAZkYgaD93
Oc8VBBmkkUA5kqqr4DshEbHjL+akd0JwLGb5kPddgT1f7i2mLyN/EaOuEneDfyt8
sJyRpO0+fcDzI+C6r4jAdPuzo1jG3Ky2Gjq7x26A0OtEToUY/vd+zAl900oA7GPx
TaEY2Q6fZt7pp1KkIYF05jG5JihzNMtNZv5h/gF//Tj1tUlwD/oT6lraknMKyNJN
ko+hn4Kbkw+X1tyazJRJrAwhvvJUElwLh3CmUUw7nPHkPU3LCmPUmWRXXi3MR3CV
gzrnWaxnr2+wD0V2JGDXSuCknM8BqvSCbWa+IbdksRpz3QwKrGJTTvmw4W4stiWg
MQEuGmzX5UjMl7dUyau98T3MGyjNqYSo4rlG2+fkzdgQhFPrGPvwYIEisG4AAbSa
4VtVvBG/ugqvE9jwFbkv55eGcRU6TqouHyQSLaVdGOeq+CFoalN8wu+8nh8VrOPL
gPLifvRx6b4OWPv9Esi4x90EP7vHyBkjNUNGwvBgq3rSDnZaBFy9LV7FkAAMv7r+
DrQZQhoZut7pfqNLYJ56OUWlZhISDenojDfQTWMafTLQQwK5O3WnqvnHj3mihwos
FTaLsybec6xF6NPfFjoUKqPR2ZO0K9zJrwvZjiTlNs4Vu21SAZj8j0bhrcvqjDlH
QLLPI0CDC06at/bwnAxE0OUxIlXElJsEd4aEzYd8d3Zu1seb4KSgeaWtdfJbTIBC
LjdFP7W4enRd9RIVe+vk1pu83HlZrTpoZ4eKaCJGr3qIJxtP2hbI4v/NQkN3pIDq
g6KCnULR4EbaUPqgP6Qm2yiSL/joC34bOtakkBf3jISQ7kQmkWD/Z4jMKHreT3nN
l9Vtk5InYAvXuEgPjDJjODyg8H0AcTsN/cU3aFbz4fmgteUETGLrQyZ4G1rtUIxi
ytU+4mSHHQmw1Wcn6fuiL7cbVCOSRCMD2sK6S1nLYnpI5KB+9iNRIy/LCk+T4K8s
JhCbpOjkydjV4mci/CZc+oQ3x63m3LXoQpNfA6glIXsvBQiKaXffigo+O2MQZbH+
OVd+g4g6SRHplRIVow6VUV+6OPjlRPrRY8xbLv24FRxbu4xPNa6MPaOEbwrTF0L/
4wNZWVlBNghroOF9qrfrIgzcKrRmjReMKxFhU+Nbkg38p7xgZ9cTzI5xbBoiMj2L
mQpuUdXbjbfcLOdVPFo0JOYODZcTHTmC2uHltkTKLS2CLpX1t+2eisTLCzq8YygL
TZDBJH/Hg3ABrDUgR8vtQ6IuMOP+884qbVy3E03QsmfxN7HpxEoaFAvvumysz8rJ
7BO0nJk+Ld+hwmXQOCFPPTzwHtTsvgJ7hFtkvCBlukbfX+F/dCBxenN+EI6ONzPb
VyhqFeVgSeLDV+04oxqdEP46AwLCyKQGPc34NHU3uJJuO9ScchpOJkQq+FeGUAGn
r7qOhDOeSzNMxwkimoFsSOnQrjVqVA+fNUu3O2HVs4fi+z6igPsldQ+HT9HBwUzT
6jOIyhGMik0SrKtsn1XXVuC3AOYPdsdE0QMGW3nV0VTKjcC1OzQnKWpAZ42+Q2Bu
Vc4zf8kYfYIU/aD6sBRXsdIgQOk8/ppEy2lD2fRRPOE3nBrTy8uJFBr63oqFdkKp
qistnrJzm9a2PwYRv6Ggisk7O3b8025Eq2nWodwuzIkDDl18ruUVksjVpzv9MK34
4g8Ztci4nxtsSqP0N9eobtcE0MWicxwTpCLHja/zJL+qhRNUCKL7QTKv2/p9O6J8
5BHPltkUro8x73nlnZXHxzoZ3nNuIO92dDOxTscl0SISUBMhvb3WJFeNhH343/z+
G+Wk9AQouJ0WrUWhW9t9Pmrh2TFJfhXRVWkuSwlXUljDB2kStupdVcqm7y4BsrKP
HiRB+sLyAtQm5mLU6fqKndi3v4w4QLyYEnSXig+M2C9t71i1mD4eyxUQQV/b6JcJ
R4SHxYmjZDnQE4tpPQQKFDsE2izvp4sCIWJKqQ7CmjMA04uoXkEHTBgeGqX4KHdp
0+hfDZB513Nd/gcnrBHPPSdIkezm5A+zV9G5eoXQbjACgJIZ6bDJ9riGWkL3inTu
+hjnY43Si9wsNehkvOYqudoH9YQOy/RI8uTGuczjIpuR6fVPj9/iQzXa97n/Scon
BX/8aXA0cT3HixYT1DEPhAFqmP0/sqXw1NFNTeCqhOEiSesLYI83IUniVcVoLZ4Y
7W/KkZzBnpRVoKnlc9ZH4H9XHEciQrhSFxp4XMa5/P4fM7uKbUnhXHTULUy1R2TX
QV1EXYVZNIfakkDQSKO6n+0+rLOaCInuPHV1gYD2mqo2ce7ImHa7lkRo2iJLN83r
2La8lqCFu58tO3iiAViMHt1TFtoWtBTg0buLJj7gcsOV+rPQGkFxPwOyS0NF6z4M
rWNqIFHT+hbTwExj6LLDx81z61w3pog61ujTbq7S/MyWD6iNl2noUTiehIlNmrSM
x2DuNHPuEh25v6dtjMTJ2qkN7W/tjdFxTX1kqfBk87x8fusWstb5Qqe8O9uGDDnQ
dA4uxrv+xzaQ1MudcD2MIJ8kwTlf9AiC7OaUUca/SJB/Qy0vlB35fXTy36VWdkn8
+HO9bKf+5b11l/KU5zYddSs6EmmFoYkB5h76+mhvIOYLH8iHH2taIg4u+lfa4C9y
JFRfi37BV2uNPKLYUXTByFQReEW0SxtjE6H78TqrRjQNkA/Cbeaz/WwAd/53uSSF
Ho+zXjntNbstpM5ZF5MzlLxIzM7UxG96XoISD6VHeYbm/d4x+1kU/B845mlQBmPJ
hI5OfkEMuwDizo0FrJ9UxgKb9vrJiFsR0G0CvpjMmUmyfE+H/te1WE9arIrJ6zbd
MYY37j8N7p/O9/cfwZ+pAXnJSYx7mAsJKsU58boFTKv6UffficzySbSaIo/N1tQk
0JSAbW3daw0HNEc/PnEm2KDquFOqxVy6WhnTlI96uFrljfdL0vqh14dVq9MiFjHe
4eqhgdDFpIDKVVhQGW/JxXbtV4vDT0uSzgwbjKuURn8rT+SuIjP8eRF06ugaBNCO
i9HsWRwHmGrBK5K5wGQBF/8kpqAGXqj+vB+YfhBjVbMusogeaqy9W6i2Q2RE7zTO
GJ3fBpjmJsHFvWlx9j2ED9MM92KOtXqzTgeMwFmbE1GcUit2CszzgT8qP1IpfDOx
u5vY8OgtXYvXE2Fj1/9AwyFQ6c/VADcfSBausbdg89eHE4R8SlWT2M/hgAdIwYBt
BB+a7tgpr7+ZYLfwwfP85+yO2sCF3ktv3FSDkSMm+T32/EM6dXdK79uEXWzLxGgq
+yjxXw79UePmpfttVl6nGAE5sN2+BuzY7oQLzrASVncA3koM5f1LRjcBGs6e//jb
MreBdf0dNH3JcrTObbfZGE07FKeT9h3oEKXT26KnXm0jWqe/HVsLkORVHYYYhSaN
oSap+r8q6rKfaicGaMeOvM0/eV/sNMAERdbn8thUmXvOAEEJMAD0HjWiGhXct1z/
tgELsnWTqDy5rCj1eNVvDXMgYUuEyWS02jecky4uUBaFSWW53VFGRmpKGC0Wsc1c
x0C6Umm2V+BPKF5HKpJ13w==
`protect end_protected