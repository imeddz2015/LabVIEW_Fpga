`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 9568 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/59UwEX+aE7FohaWu0/8IpTj7mav863zUNIsgIH2BWb
Abd9opeuBjbGF/waQMI2vMJTwD1ie1YueHc3nSNpEh4OXp8P5ybZFY89uyGz3ztU
W1EsuUnchJoQgbHZ/sLbgtGRgsrAFn+ZoIeGN1d6RAF2wAESJmYP8zw+p00RvjZ5
yD9zY/ULOZvQe9BzlxVW3jX9iLq8WXos9tOfA2C0z+Ri6oVKaDt5ZR/tX57DMPsp
+4CqSinjPQmjFsWyJdsj9u4zTAtcRtCDYkYGuc/ZgbLKJN1EQN+Mb/vB8pUZqerx
UQvaPaiKkz4enaohuKBFoZaAymqsV0I0SJSaj0gP/hb83Fji/0HKYiCfE9eX2DGN
TObi1BadDZf1TXPltnYA9xnlwT6OS1zOn8CMYowYUIXpg2tl8OMK+OwhXoEI8bL2
GDweuwN4wtmxOUlp9kuWFSipBsRnter8ws009tyoJfXDhAdPOVinx3CqTHy6gJrO
olgyS8F/fBQ4AdioKdUyCHg5dy/ssfLTJ6Xs+oREz4i3wphrd5Vas7HzMqQ7IL/v
AmyBlAinHwxAbg7y5N+nLa3rMAGjk6mT0EW/x4GhUwZ747GA5a1LdqrZad07Rjtl
4TAeqx+iv0Y3OL4/srDLLOd8eiLtr+NuvS4ZTjILIRQekxY54RjediBEO7+yb1UV
VjApvL0k0sMYse+8ievDPYHE4QWB85E/lSpyoufdC31dlM24lPiNbb1vE6Ov6/8H
k6SB1Dtwr3rvAjYhzuL7tLdqJgTjeae798P+EbIr8h1D/leo5lY4psvTGEh2ZhaL
7jqvIhQxQfMCUXKhrS57+6OhaqSvYPZf8ZTdUKrEjTyQeWSbILGXJ6nSafVZ9pQm
OfQVDYwnh4PlH0LRn2exqwdGKC/p8q/7AJEJuV98mC9yEcTEVkZGc4cFouNbbmcl
dgL6QD0p4sspjS69H2/+h/Dd4y6RLJcGu2D3R9Ye8ltPtlUy3IuIpKAaeKvHceFU
q8WxCMCXmcN3aODNp+4cKTbpu5oIM3ONJs2ptJ/EJoTAff8WmBSAOPMkxCXj4LbA
mZkTKZI09ge6TzX0veUxMT01Ikpq72H92bcpJYv/U2OSt/3PKkw02ehkWCn3UXEG
nB+cZluEX7Z7NvsbqvTHYciGCI2axBVXA1ov1+H1xuN05USUJR4LRnGLoHSzr1XV
BfKgsKly8mIB/KEA0XUPspNUhNjkFTDI6R6iyLZCrGOL6OaJ6Fb8MCZc3coyf4nZ
2InD+gjns8VdMBAHOI8gk/ezqM5WRefj7qai9M/2CXMr+Izh9B50sTNsEU7+Hbdt
6G+i5LqpjdYX1bg+kmVZS5fY8xsFPy20nk0vLw/sq8jENPDPv4FRlJqu7tXr74I5
WcWzHi1RaIS9v37wT2RpQBTkrbUFjvQhZSFRTD6D7fu6Cv+QBaqDTxWL3cOHkodl
4w/J1tFl3XUHZY/n6XLoo7+uw6rS6T12CpVrWwFStCF/Hihuc6sDpZJSQgyL+S8n
yg5YAh0bEl82TwzuFOhT1GMkhztNuomJI8s1HmVHGV/mKnftpC44Do3MOwfegzNW
e2T0NUvzvQaRkLWZsQ7PLvCYOLskt6ED8HPl5XHSy/8cNUfu+bD+zIJcAYc6Y6up
7nlduob+lLLwx2kQrVmDTroC4SnoTmeD6ed5PYU/YlPW2CvAddBTuKzQCt5sR4PP
1FUrb38oJAVYMpCCJ3c/2N31yHibASRsJ9ATXnIbwK0qNPMvlyHL57QFd+WuRYdE
y0NWe7rkQwmwlwZLeZOH2fFmCgaEu764Gt2T/UMZoYiCEp2EFYJiIx8quKH2YZpk
hivBWLTKbvLkTDdtGAV8FYyzGeoSGycW1IBX+nwTRjCQZzE7sFS8V2aA27jx1USF
3m1FQMTdN0aCcsnEDvHVNEo/sGvpCzFL0EvM/3QRJr6g7yKrT3f0gY+qdj5qL82B
ImyzDbRzuXjssix+1nq2fIouYeTRhDk9FrPHH/GLtmM8CNezpMDwGkp5LZcluWRZ
bWRLInPNeptYDp64ACMVh4QGvoLw4njlva4xPZ08hcvozLiWS92DDEsUHupz3q6F
N1NEKFkU6Y2l7YwAYxX1+Z+e+OkuVx+OAbLyBJPKXijW9O5NRuyPQNLx9/JOYMDo
5ucPSWDJjOvfXfZrT02MyxWRdboL8aGkAssJji9JC8m/bEE4UhXXk3ACIUTwuQ/A
QWQJ+jYvcRjSNL8j3/T/YQ2FgVk5zaVAdOiWLTPZIAq0vQqW8i00/+dDL14hTM7d
IkQ/azBbYJwEAwd9sQMIC6y2LtMtGqiezBP8VyzN6ymlm6woQ4qgqw1pcESzsO3P
MlQBBkgumOwYa5Cm/ZELTUiO1UAikpUZ+IRjV0qBNfD2+zZFuB0MJqe40wTY32/o
Ur6mrMKrT+wmW3zpM0KHRSVafyKjSr9zq/jzWQPvdwelM5ok+JIL5cYtKfXeh6Y+
1c/DXtb3hmD0umxliQm3evjRrQmmLQBWQUm0VTTClfVnwN3a2kz9t7Jwe1UVBuwl
AiMHq/jtXwX4T8YSzqN7DDjOj6rICzJgJ7UC1Ua+w4ROwhztC3zJL51XLcf7kami
Ipg4oRWAfHKq4fxMWTtNuM59e4gOMUadJveOMx7fZiNAz2fT+NwpOWE2bALvqmf1
EnCXBYdEcUDYqiDY6CchkKpam802j6H0X+rs8e6Nd+BgOdfFK9nYXggkSfQPvaqI
IIG3ifQzaVL6J7enJzHSYD37tB0Nw+zEum6A0p5JMVeyfBVZFprHoL/L4/DlvQG9
Y6qg7pBBxIb84E4821nNQgo//cR0DQbh4SqNZGzD0kYs4bC4fAHFU3jZGdq9ChWG
/8ReOM8o37aSY+JhlF0OlqGprKWKHCQfS9PEtxlXCnmBhvI/P5lXLzRits8+z5UR
QGag1dFoNsJ43HH/89WHr+FFlX15azDJyTWughktcORNwmEDh1vO2iMEBkfr9m0s
Mom9wGC/QMD/PiYWkcFCjHtU73rfql+/7jWJY1YdV7KNMQxwd2hSxENX7LcfmKbT
UufSvvI9jMIeh7+8jqhQF0CartbUyfucNOqEYvnmiOsNSIKuXWacOxWcHzwZR0uc
yzNhpiL+RmuQIM+RY+C5MuGZSjwJtQsWDj8icAXJtNOqDlMyReRJRtqX/PHo3hvz
gcbL2FYFt2BKHPRmuZELS6BJaUy6ledZgHx9Tluo50B3NewS8RHRF6plEmLWU1Cb
p8zkEKh7a6LyxmiA0uYSCq3BnK+RPylPy5cI6dybJxjUG9fVl+xkgzogN067N9W4
aIrLW9tPWtukOiN83MyZ5m36vlMrgLhiE5o4CW976SkrYtMURW/mHVooiNfN2fxx
Qmezh/srrf6y3DwD8C+0MVLkubO3+8DDo1HtpMy4DFRGjNECwcF7zT4tVM0uSfgR
RXmPh1rvRmlJrZ27bAe1tWKQ7AspDP013A2Yyz54bC5C+TkArkcWz7BnFg193ZWT
4VKM1n0vZmpA4YTsGyPQTBETgNgychHmO6QICz1/AkkkCYjt4o3UI/EIOwZyiMwX
csl6jiwRJovOxuNmYqNhdkd+cqI+OgUa/8gWLKw3XIiG3ceOfwyA7VfKF/cruJ74
0cyvwUM8JEW8FadMuiNrl/Zzj5TJZ72zz3WZA05LRB5gdj7FkLJ6lodvflepVg95
fU/AJQfphrhULXpKvxKJ7lDJvKv68Vv02EoZDAiZSHpHPR07dVgRvc+PL4ZqPdaF
rbTUJkgvDfMuEXNlHPw6jVSzRFgZ42LhDpc1xjJ64TlzFIN7VcgUMFqONMexUUJ8
3xVFqZso7Eme9E7N1YDKpQNLZf3qWPt7u0bDaZHFscYI/vcVH2aMXtBqUXkqzM8l
nlTJfT3XqgQtsMsrt8b41l8FajFsUotG4h7OEreJQmwVnsGZn9s8Ex0MAfb30G4D
vLEHpBuWGQXcQQYXCt5/jvnfaf/nxAMGzDzf6/slXgPDoz5q5E3VICrahusc/8CN
pCy8L0Qw/UywOIXJHTtZknZ538kH+9o3tR4+JEG0ItgV5IgABDwzVwLEuIDEGqjg
MCkQYr/3PZCieYVIMkNTa48X4cPAfRf32BSKU9TG1L34P9jvLxbLhTZL1uf47bD5
NWVRCW40pFGuvaPMlS1/HryLiOSKXtRbjx1yFW09cnFs04pWifgz5+U2MZkDXo7J
5zzWjKxZM/ksq5p5M/qoRiSHZq6ptHLJ9ZFhNrbPMWskEzj8qnWD9enJeLPyNDD+
MnIAqY5k1V49KX7N+/qLPkulHmgVPNYiYEmKh2reg7ZKBWHAl3u1mSpHKcTtHhzR
uQJcnkWr75zNy2FCfd9FxU1SplfiqzYOsbScMXpH6nk8yHWJ3T2xNjFcuICzqwlw
hhwUiy4b3BEaeBDKakXuyjLLdOP4U10fvuLTf/y4av78jM3lINWIbbPm/k3pV2PK
Bm+b9o/sa5bySlhVXlLZ7EOXUUpzy7fIzWV9vEivydsvDVPRuDeetAwkMkqrUyur
KxwRFAabDbIqD8mgEifxJ5qFYii4pO+jPnKHtsf3BkdUC8SHcgXc7lc6NkzjKmww
D9oAf3/N8OoE4DTHa2/CZXHdnpZdYtE4veSQyS19TS4WkJfGQ/vho+Yg/A5EaeML
3r3tBOuEaWOsaadyGVcdSQpGlPnI2zaxkqujcVpDw0vKA4DLb9mWzA6/CMNc54VN
8LRbgfS68VXN4+4We5+kZMclXLHGNTrXeB1PdzDWGL8knJMxIJPoR5r4zoFJzMIs
6Xn3aK+ccAt5+poFPiPT18xn4aTznIowZRFl4mQ/HECfZTxI0ZT0cV5PFx4wrAWL
XrbwNR07dBXHsvU/FJ2I6DfrRD/k1KFC/VlSbIPf1/2QDVa/o91FPpeuRECbhWAk
a9EcNAmhjilz41UyvKOdXtJNQgF34/frIj/3Zb3NNkV/AAjSHsISjwJsU1X7opAA
2yhEWRU67u01OOtQ7Sqg9cTkhibLnlFOWvgUZakp2/eB2x86mR2aDvxCK1yoevyG
cX//AIgwloF4Wki0BtXxM3jfhBaulYs0TVTb4mrqeU27uFPHGVfl6Ci+QKhMKFeh
nPd4tI/46i8KSHRzC4cODkr3c6XL2ukL9DkPqQu4XOXC/HMZnNPtH1ftrjMBjhBL
AXH3/0SMRGTDe3aX8tgDcOKMrwUBY66K+PrqYSY3Z0Wte9UJpuESypQ+hRfwjLTz
BEHuMi9QOPdkhVlrDkQE9iQV78P9BAQEJ75bV1ofwKzIDyr++5yxs6PepjGCcpTO
vJN4IMx4nKvXOK3dxvTQXfdA7MwowG0vOpEBuMu861Lh8M56znRwbkKmmT3VsEoB
8A4x9egM+s1726Qr/vyTWGGkiw66g0yechljofhb9wz8ab/C6Sv78JOBTI3S5TXr
vtTVab4zU87AP6f8QPLwReqghLExA6C4RVrR2KKLC/QnDbaoJmR9HEiPAwi2VlwH
yRUy5xWGNuoC9ovWQhaJmE/Qe4PV1wdqyEVgDwx4DoMjlI6Y1qNTfT1IElelaKoM
pDLwmgKGnK1cU9Bjd4UeR84ePFQ+9FcoOxha4HwV1OTWZRasXSQvLnO+ZiO53YB4
yhjcmQMxg4eNLdxw/u6NoFxX+fpLVzsqAaexUvNs/EQIVF3JKOXqNwvr/MTvN5Qk
D9ZEsp27nNIOdNiFTZSrbvI9V9JZkZs2xear22FsMG97yRHgVI31jdHnCDyeFqjz
9IjMgn48acLnoZ9hB/DAN6ADovFEawBC+o+//uTZK6TOQaFCjRoOQsFvPZui8R3E
T9CWY6+BFN/DSDLi7eNr+oawuIaQsumcXPmR7k+/4t4d4Hfc9VLLf7nk2pR3CUts
BDzC0kwaovD5qOvbT9z0Dt4FqQs6nFn/uecQwJKsMUcjqYPsOlSdh2fCv1v/Fb9X
hFFi/QTAIdB1mms5LqrOsvukBfNYuTix7WJleFmpxsfZD1kns6B6w04sKRMnbYdk
FoWi3Pjr4LaO6wwb0JZvD5sITo6VuogIJTxp5uC7YLyrngTpKLhP1dslSVQIBTDU
inPJB0IQI3tSWj7/9oUXhhR+aRKuQKRq5lAe/ZDDXnfKIdvamJcVUdYG1RJUrFmO
MviQySebBWdkHg2kA8UY5pvnVY3k6BVhc997exHyIyO5iCRG/3kQsO8YTkZOOJrr
iVvFUjTcrzxGfbr1md+5WCiO7tfNbTlsT25XkyH3tEuofAO7xDf1woe2NvlDUUZk
5P6mXy1ixTdXO6jZo3Q2Tvx1ykmPsSL03GwU2QniTA4cC/Go9peOYQy7PSbs1q27
G8ezkbvsqjLAApcZZL6KpFY1a6S2MXT0++FfMAtUkZsm/TkBgqKv5GWHF8LWrxhM
xWGfDeLkKY54FGu5oG42gIWQdAcTrYFa+qSjdH5OXbFvRHdFovO31A+7+dXKk+u7
61N50jbmB90r8OO43iFRNLIChWHLlB9EsFhBZPyFRfFl8P9O8llhz+8+vblr13YF
HHOhUHCzZVK3eBOlACJgfrEosJXz+EJpKc0AAfRLi7cgqlgegHER9aAml4sX6gMz
6LcI70GpxBB7MSDTX/KFMBeuEGAK3rAyrpqgJshLLmgjCd3XDqgg52EYFYllLPCC
fV23yK16udmTCSJu8u67X8bSUHH1IujyDsRcCyGm/aiS1Ey2f02kT1JM9LkiIklm
PO9C7yNqcRIJZIu2agu8enGvwigRCL6PJWfahkY0xQwBY9GvnE/A+S9Q0ZASDyim
oKToHTgJgiRBaBiP+aD21HJM7RstHLeh8+spBPNWu7VXpHJXpXWna7pCDB/aPHVp
n0CNBymEh/9WPWidCtVI2JrS/aK3fFQw28qXjdgf5zZnJMW+uISn5Oe3+JG1BEdm
G1Bvo00mPT6PsbFmmodsYgCsyv01d1D9qrS2n/axCtCUX1BJQJzYr4Dfe0lFqaGO
7jVzmHfwwtmm8XojwLYiWz6UcyOMQdJSkxVxuBobSLR25BGyN4CUSKQ/20z/W9uG
R9bZrcXP8PZr0n/gnSpYUFHch04m5C1Jot+zZ9vlXkp1dYPdktoJOQGnTm+riy0C
LV0tcUyF8zQGdqbG/coZ+QogwMLCkuM3e1xScCMejctvZ+PMkiuc06koQ+Drh6oJ
kOOApXmnBctr8CUsGplBGWf0HcLA5uU34DQ76B1ag203J+W0RW4EBAh+jiNUUK7x
J8B/94uqO1seU3unpgLvqIYQkWLMWeQfNIDjEbkDCMk5nOc+ebRtH/68EX0aozp/
67vh2SH9K6AES31LS9h61xa0lfVYrshMzN/Cp4W641rux01aoTMIFJrmRBJ77zF1
z6TdTjwh0ZXmQeTK4fMCs0V86Xva2mmLinmDg4BXLZE+dVjpLSjYfUpcfwwSfQ6D
DE4EoDdAVFh3TOXr3j4ncjIOl7m4vS0JXW1a/bZp0kHjqvoCdZS34ZkGhT13jks9
N9i0juq3k1j5u8CdSVjHi2DZrbwrPGSybt3Z1T10T5xKX32PE0tw0UpUkWvwaDyg
/H5krFxiq9Qlb10pNUXpsitE4ZwQh+Y8nsiOW4wrWrssi+Qej/eYE4UvwFzGAoWH
bkKb+Rc2ip1X7duDzXaLjb72INxPaqi8xWp0wN/wA8+6/x8Tvs8lGdt5bvL1CND1
wU1YbhO0zhRIeyGdkYBRkfduFF+s/TQ8qXZ5GSeMaDwltBzhlZWR2Tp+EHWVo+x0
69L6+h9vTPsZQbmPJb9olpADj66cStl54tf+WddX6mxRmayIPCKqmzNGpWHwy71F
9vpzfxnhwq9P7GTE4Pyi9YY3pVC0lHC4i24+qS9eYy79Ai70cITHWOSFue36fc/1
eqUtp0nYQr8X/aX+U8ztToHmGMl5pwc8VXVx2JUJuaJlIA0VLqgzPdpLWkawySlV
EryD7YzsLVtTE8ekaXCo9mSBpKZv1qB4YhRTKd9LBceFQTUzHqH2yzk58xvi8nBM
Kxi0w5eqmUfZ2sveaJqVaU8XB2z+21hz8ENpSpxgFSVqVAFeqKw3kWzz1qmoyQTr
4n+qxKhcQO0rj550ZemxaBCnF6yPsGnXd9+G3VaEUvvz+x9OhImblEXJawyjfWi4
lol3K9oX78TRnecUd76GijZD20muc8D4UVrmVjitDyTqW2UXP1EusREhMpwGVSdp
Y2I5jR73Sp4t3gMWNTK0oWf0WlUl3Eh8CONVYCThPjgYUHQQWhfd1Q0OPmMSo+sY
9orG/bf759p16TmI2LTVEpUNKmS3+C3mDAgq7f+702CLMLDnt7DU5pRAB15dpWRd
ArTw2mlklu/uzfu/YUyBumtg04ZV5IUEYl+JrSiqPBeQZoIVbqN1zhuWt2ioYms9
vgPSZaIIBfgnV9qrItmXfm4kgwjryFabIct66gYof5VfggH0mlZ7/LtyYJEuK0lb
in06hGiCEuEh3tPI+JiQKM1IVHDzeS5cMHueO/iCYWdCF1wXzyTjtKyavZoaGeGm
43Nl/5RXC3vgJGeH+0BlXwNi+1tkG07ij1x/05tc/8PhZzHRB1Q7fs+he7l3A304
/4gBDdT+zCWswHB5bOPwr2/IGQBFt/heTIsnMQ1TrSXBZeL62Qzkntu4MB447r1/
cgs2TvK524qMe1XxoFmN5OTJKeE7QVkA8jOl4mVESn5bmJDshDdqu8VBBpkLhXfp
fzcx6CTx+Ggjp5gm2el947Yli8YOys+XGm/ZvfOdVitNsxvrRuuRIHBnDn8sOpWd
og0sAmdufdpDqWEuToJlREjNw9mmke+TyoTyF8G8TYBCJnNjnZUWNIqkI5RtmEIh
nKVUmb/8jM8hzk0WF5qM2OfpoP4JpO/lqrzrDQM/A1pFtpl5umQS5Bu/tjAor+ju
YrYUnWVds6qyJ8dcYel4h8loB4yrBgJgRvRblxoGsqD15X+yirbxCAkce3xZhPou
BLu+1oaZ7x8SPjoQTf9qJdm7RWcnnHx/qF1VKGOvnL6QJgKXEXFyNgwwy2i5Dheb
qJ0cCayZRCowxtReuzdpfhDTbkC8WGLbua8yE6fCZd2MwX/Gf76Fy0TlGvcGqAkz
9zS8ZlhxyEsLZN8WxbDzIE3R1Hm+EXdmAVN8ZEssps0MhLEADyKGxARneoUofLtT
vK+GgVy7qkG45vlF6EMnp6pQiCujE5Xj3MBqdgIpjUDvi8g4MIehnvXl68FPWBGe
5rx13sOuW/6+8wyvpRNneI774ljS+vt7QbaO8xPcgmzFRpD5Ox/j8HO/4Tj04U6Q
iwP4AsR3VcC2Jp0iEJjjcZzk63J9UxMHtGYoeOQQKgjVfvsaiVOr/PonVWO27tFT
fPGqIdXG54dUYAI5qgipymJf9C8BBfMN+sdnmfrB+Izm3MEX+cisZVhpARs99zyC
J1hh+Px4t9PFAZTN9hhMzZvsux+jx6AAOwEXoTIgdelmp15eu7MXwD236jZLgPhK
q0k0PussJt7OmTxmpwpbwjD5beY5QFGHc4n/81Gx+j7IXJShk1V966z1kg/HahUy
mYiss53x+ETwOa4ZbYeAbWDjjZKwZ5jw2owEg0DL52eF5LvD0YwuWIPCRj6pvXjV
q35J49pNkipprxtkHRMiuOG8xfMdzCRBFw8P6z332X5KCPUagmzQY++w0gEyrDDr
N3gm926appSPKYUx8+/IGiyBx1nVWCINBySI2JMBuoeXTPk3Zkk8Wuxyxng9CT+T
AtXUMoy2zcjp9P03fXFQC4vO80W3HJg4guexchlY46s0O/psttGeZZIiZ/Vx6vx5
xiwXdMeKHpro70GBHuT9vOfQOnRX92QXL13uYyWIhBzKNZkX37dKrU7Vh6ADStYM
sYC6WtNEexv1wPrz8z43H/gNYCkDN13qj6cOedTJFL8K3gTJ5h1IQBb9JlQ+HfD8
3p4FcC7Qn9OCQfZFExveEMmoRwOSs7sXXFYo9vhkgNbx7auOCdHiYWBVKMtYJAu/
rXSIu+BNf4gqETMH4QmQ5xkFzzY3Bx6QJrwH7Xjo0pJtvrT1vr6UosedR+Yl++gh
kWIrQfyZtqv3kNx8CMQqS+Zy9zQY+oGY0zIH27InOXNZJpPc54JensawslQHxfkw
rXLUP9g+HAD4G3TFceW2G/Ps2ae0K3V5SEZSaDlylv0SSgqhBt7/Ek0PC/2c90AN
CD8OAO98da43YCS4HLSYxdMpI1POf1dRfF0kDC9eFpJKrKb/zE4eouQV4H55sVaq
Txyae/H2dELiZSgtjyoc2GbRsjo+PMLw0FxbtU6SRstUhMQa2Dq59UoH0LL9JKSp
NyT+u1LOtZ8UFmSgKCny59IZsQRMbrD4s9LT8JVg995093entXvWN/1EnBOHDXqS
D5CNHrW67PrbFPioH5qyX9qy1MK3wo0cIUni7yq0g0n7FuIcxrqaAgHaxeO/jQ4C
oQr60u7EeMMp9vRX8JM8uZiFfiKu54rdrIjO4hK68R4MXBH5sabiiZKoDmgMeBuE
HdcZFhkW/nGFF7xsDVmspCPGXyWutXX+I3pZeMCs4oD2KA5QGIFprK4yBBAH5Kqq
eWrPixohAy08sntn5Xgpw2tjhV/VrTklno3lT1K/99IXGhdxOFJI3AIjZdmYvsRa
h4Y2n8oWTECFZ2Q48z9omHbZnjzfRbDqimdlMR7gKVXAbjJF9LUpdhVh2qzgWp52
EPmb7WWW8dPQpUoCMT94d/Re0Qz4cS6YMkdDGZ5vneS9Y8PfLLVlDkx6OgzvYb4D
wej7nBSKhM/n6fK3lssrZLk/wneRA100iVCMq+P5nSCYg3CfFm00zAwSqBarD2EH
+o9ydLw+rvuZieILjsXGLapg/2uhhtZX/nRSYbXut7E9oWodTjqe+/fzG9nNxg/1
+4+8afvDXzxTzqqXhhvW+ZMzfWVNDdNiqsI3aIcrcs2OWA3/wBBeQvrb3XQhsOA3
w5g8ti//m6Rug1Ffc6GYexfRq0Z/RZkZx6RxMHXCcZKSDh1U20s14HLS2JG6itfB
Ts42L9FjklJ9pLO+2L7fUBlnw33Nc/h1EJkEjQOhgGp5ZZsnpCLf5bbHlFHgcDfw
a1W28nFr2rOxeHcmXrU32xhBUibor8t1nqKzg+6KikgOCYZDEKflt+v+yjivTHe9
3m41RIPVn45e2i5uvmU66HR/7B3mK+Hk1HE29qq2AA/77NzC6nyyXmfTg0sw4FOr
4JTin0F4M0jDPeRGQaBHYps5jdGRSC1/3/4NbHN9jXfVjKnm8AJwPFLfIuB1Rslg
0Em5FB/4cWb9/NlUyU7RZOrJ+JPsylvuvlvglewJYQe78M55cU3QEPpl4PYeOQJg
xiu6X2C7WjFk2hb2l0WK+xgmLQ0sBeL4w/pP+CMpyskOZUdF1OqQpysxFULPInV2
g7g8euTKnEmI36o5nHRokhBh7tfEjvniIebICvctr69mS4ajwrChi1bXOIVMTk0I
VIBob/SmVgFMcgB4P2CXnpenKsv8fyQ5kGwZUmHFhZGzbavECkSRUnPiVXWGp9qy
qFksaJr/fLo59qMKghBoygPoDCltVFV5iFeAsCxHZV2IU6sc8TLdPuOs4/euWyDz
0CZfIhQdUIyg+MtaHlWu56nWY6oZU0lbDvQ0W/o5ejxKFFrJw134IhBsW7btfTFi
eMmjWMSWIFGTSZToflUOMAVRcA7pt5uW6NfVwYhnfXVQhR4No2RJFE+u2JvQjrZ6
RNjrUIQNH5Fn7Llm66+K6DCRgvklYMedgGk2wzz5vK99vlt18Bzv23lD2mjWmU9G
lL9zUAsN2VOHS49/Pp1MyQb/KXP6kupOOWf+n/vXW+TZijJZVVOZ6Giw8RV8UtoJ
wZintHTp7Mm6vOpcvMlUx9DdvcDXyPJvl9iIUzCnQijKoTtmyt6jPFqriytJh2vZ
/3wWlFhn+WDSBzww3ywZGh7ugXzYI+mpYfMRvE7uR76r/AFUOmsE/19f/b7C8zRb
Gm7xS99VwN6ggkoq3bt89zPJmRJVAEDa04L64C0Fx/gTIXFo5G7jffXDVkLnwdG4
7l8Bqa9pP+y/0tb390uiIoQt14ieQvsiUSMDitNQjRPzg4uRN2Qqgn7tfsvEhnYe
/JyKIczfBLF+sgBFG8Crxqz13MPWwS+d8e1NPQtfQFQTjpZ195YFWKD+CT2aQbzB
JCnjP1ab9Vs76NrK5trWoP4d0npg/KWL/dTc9sRMGLBssLT9twURTcL7Hw7H6nFe
CCjh3Ab0Bp2r+SquWK/1LfgqzcC6CXnkComLwkUoCq0NuVADzuUx4vd11OmiVWNi
YCnjtSI/tF8nzrkM5I14Vq4WNtgZhm4+A3VUk4KdLrC1RKG4dBu4hbGKqM+VBlOB
fdpMHAgy2yT6Nwxu8hfBLd6bzZ2YNszwUcU6TtqZTRm9WFSjywJ2ePfbk/1Btrdo
x/znLyzD+snNKjP2wMyOmxZc7NAUGuJo6/JPd6st/UZRDJYlZhL9V4icBQGbHvhS
wGW8ckHj4QMxb1uPtyGnsmKKk9Axo/PjHne5PD7eSIMORZCvnIfvqqDSnJthWdNX
yOgGGVwpCKpF47t6rB8K7c5WFOHRGdRos2W4ikXIAG8wAaFpQOY4TstdTgiUY/i6
wXOAgw22zOrTd77Io4fPU7sKmAhcclH70L9thnsUH7d6b+ONWM/E0cxT06izk+Vd
levt7lvrphb2hOMdFGoIAezX5emer+ul1VOEY5yAknNO0CURA++m9y/s4n8vvYm9
AEjKfq88jA4cxsIKF1NhWg==
`protect end_protected