`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 12176 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/9huKRhRMtvnNqb3Z+UU7TahEoHV+T8U3P3ufru7l1O
3DlgtZzb9QxCbOjthp9+wDkjygH0eUfDrEl1ovhZG63CmpkOuGPb7mnYPAOoLRvX
2dfKOj/k9PDIv3PsMFyC6yuhuFbVl2+Tam4yZE9I17oV8c7hWE4u7+9iOkfNVcBc
6Du55LJsyaHqm3pkFbbQshH63hZUTctuUIc8pXXZOafFmWEopjz8AWW/kszi8JhJ
7EyKSH4qoBYuLKPBwDCs3YDiVNTDYsN+a+/fsaw3onB6v76df8HKA7uFHt2TJ46L
YW4wMg8fESsWUEws3287Px+IBUWB2gaIDgvw24FXlQmyR3Xio57zUeMQzkBgpcpD
1tzIq7MAeFVdYoF8+H9yt9Nzgnckbn2D7XHbJULmwsGPj+/s00GAZcV0VrOrHqLW
JQzIVdlgc54ebVUAo7TA6rCW6adIzmSIaKE5Tf9bVIBKW5cgsfLruPMlyEi8Lunx
QulkKEqyJKO5BzBHH4bGiq2f400CCJLjZyOL+iwYL2vBH22uZ4V21wTgworsiS4D
5G0X+74eaq+NwAb7GiCAZu+9L+RUZuO4O23btofVBlUAjD5QzY2gzgH9roCF2OtR
uznaBWT1ctwM4YRVp5CVdeseJO4iPm7JNcMThasr9hNFeZlNjQytWWv7fM2dI8Wj
+nOqsWUS6klywmVFJvV/wMorh/QLwcApG0m7sesXjYXKWzyLmeVRf0NcyIRikUIi
tfg7VT2UyjtR9cDbI2ySuaidkuhBCjf57LJzE1kRkkHqotMz6nEuZ5w7AqXBqL/S
5RL06sGTacdQbDQY58oX9JliqxOnf3B91Yh7n0ae+6jlBMWOGDhVWWoM2QnsL431
evrEUa4jh806/Qy028oeWiV0L0Z+HCIQ824BJ9gXWFhUzuiZ6aIgGNUCn1txgm6A
hUMkAJ9VhdrMb2mQENN+oVm6TrYv5byswqrJ6A/oUOnPvSop4QlPi/+/rGJkSzsg
QFOfzOs86saizoFiZPYvt3ostDwTgmu/iRM5V11dmq5Yns8hVqsk9/MYnA7eResp
ug3UDBOOXfDiqLkbRVWVcnG7MUQln9otZAfA36CwpEsxSMqR7sYyHAUNlgkfpy76
EzWU3assD+n9Nq7KZ7VjFsW52NM59V57gxLGr00KCUxPw6jbNwUI2jzhKYS8fXsn
TXtkGXhuvzew1XvtWVDqbj11AjlnxXGz4Bwzq7mURqHg9irBywwRCx1qvwtD0x/w
Y3tOWxnAukUeVpf/GbgDxvae5tdULssPRS3F6IbZ9EkIQSTh6gVIi3XagvtBuRvG
42RkcK97SJTRmLueacI+1HEElQ2UhxInqvYfEncAmBovYHXpmPPubyHKqiH9kxeU
NGlXrF5eXyZKJOBqpmKciRHO+KyC/j/R5O3hUNWGUtTkhzb2VpbR7XuWRC3p36uM
IH3heMGlcFLxhC0SrRTFSC2uy0rNrBF6OCflozuEHA9RXZDsuFhpTyPDm9xYas43
YMlg4WVjZjDRibkPRBghvK7ZGya+e5CWObonH4/B34+D9u5xZUi87Ou2JXMMnSgQ
28w1veIswmmqiob7wHCKO8voYyW8offtu3KKkPjEZ3XyNpoFg5FupueYbxd2vEjF
P09RErOPaDvwycWuIHbBQz1qgwbswB49Oym2H/7jWEj4KRww74tgz/3ClucJySEH
/Lnz4Wx6y39FkkomflN0H86gHrqq7DIbbHgKaphm5/BZ2k5vawZaZd+lOMl6r9p7
CUWovIb9hbL+dT0TP5RLs4mONPuBXSvPHOtxIs5yS2a9MLqx+Gm5GEftofOvqXHS
hAHa9IXUvUmoSvx/L84Pto203eoh+ZSVFrsbS3YEAVXzyN3KdBw95D3YyjDi808M
cJ8mt5Ou+wDPWDIv0eD3VsXuWNfXlEt9o6/EGBrCR/s/wa6Qx+NJLK/5RYKbwTLl
rTVWVTL+D2Brv/kcyIShrvLwK4J/xpHx7hGeaeZTXdKyXRi9gck31RU2VjYXxeO6
CC/gCgCTEx3AXeGvR8DhAWXGOUgE8410KUCtWGRJvqly3cHIbCZN3InXdu6k4LZ+
8WCbmcjgYCyW2U00yumPrgs05MPbOAkIW12ni6hgIG1klTMp9jaMmMS9G1l96wSb
M15oUPU+IMGc70lPRZDhAWXj8hg9IDvXHj2SQJjDdjBZA3zUKJ8ndWZ/6z7Hdi5r
8mPFLrJG5u0CEDigGHJQXCNXgSRpIrOiOTLL+ciQJsQsZreOF/hD8b3HqM+WhRzb
QJRxmykYPeBYmBB76xKc2xPfa1VbYpa1ON7un6ea+jlAQGUtxodtJY9Wbxb0x6+c
FXLtOixvtFIDRi0tppnMEpCdeft/jDzYVcZUgtsq+sQE14yfAuDDzX40l2pSTqZJ
dwQ1UTNMtmXNm/LLtkWZIebf3g8K+AnAaXt/I4uMHkoX2s6oxQegA/m1UWtpLSat
MMbkCnRsNE7iUCzCaDJDYW7JS5bOBQs0rBA363mexO69HpDEwEpYVRQ5N3QqPCVM
DcDDmJYvbErR2LyPJXhUST+CR1lfOUvskNqpys3k61q2a9L+6wgRaznrRqGLvFuj
XamkLvsMpQY+nLGrOyd0GKw3d86N57KcI1D52hz374RTjB4BeaW2GP2JVHDUs3pq
NndyxV3JjhhXtBJr6OVLhuEb7TXdlPXYIMt29KXPm7eUVpzky957CbGoxRU5VgnR
eACtEE0tpH8zSLvoGKtoX5oAP0wehayuSNNVOlRXDjYdDoU8QrvC7NZSfPXFwGHe
2JMbpX7i/ny6gyRmMZSUV8yTgqyHSSa2mQREVSF0JhMmIYsMWN+CK0WtsNaXH9yd
cWnakXwXUjS7LGF6l6uSVIte3+AASPRCQjFDGRjW3wwSRwZlECXFw4jHJG1VPUOj
EJrR6fA/rYntikfzbsg/ApHDJukgnFPxBmWuE3YfCrF62ikf22TfKaJNlntYOF9/
iA9BPO7CYhlZHvfMvyXLDOEF3k0EM2DVWtdBVGKEz3i6kCnv/OnoFRY6DjUO3b3L
UNZpbQihPFv46S+Sm+mHP1cMvq43++89HhXvNOoccPqqe3KppbE/nvplmtCo6KSR
FWS9Js7m2A874gCi8faE4HE1vib6PdLE+FROtta304FIXDjPfDrJfuvZlajY3OSM
kc65tBQdrU8m4r4777wYDIqo6xVN7E3/uvATodL2+xwFFLOzauSVTUOcXF6Jd3oc
4Bhh4G8nT/d3V5R9A83GHq1to3MapKANxLviBnR+3OnwPQ9Z78ONDiN3A+hiFmHL
ZT5RMuUbJXKl+tNOX2D6Qrvk03nOtoYBTHsX9I3LjwG69qoDyuWGnG6CBKg5H9v4
nv9Fg7vg/PuHNJdZGrhGAl27nGYoAkvGTpWTd9b4hIs1xAjLvqqIQ5EX1qvAfdDn
kO5waCvWCret4eKjsqE9f4+F8LiJNXrnxhZIQquw0ArhQcIrgTT8Lp+J2xQXorVV
CXVIFSBbCJOgozlwimm9/ywjpdu70Af97dIk8fnSPEfWTtqIghQU3eJyrKcbQnlO
ArX14gi9G2akcM3AuA+y/rRcYqsr6twdMZyUURJJLilMmN9IDKCOJPNAHQABXlt7
+a0kARtzCDWiv6mnUwXETIDhY4GbxJ0XA1IuqGLXV09qYxAU3AkNp9ItMAf/fNIx
HS4taOz+PCGzySSt8RsUV0K85FKCGn8sSt3vXuLKD29LpVdOnJIhFm/Fgd5uWk9m
qH3j4OcDJmr9GLNarAtdznD2/rAa5uMfOM939swzKxYTN/5Sz7gAantUCL8hgnuP
UxwlAcLYFYccPQbRa94d7ORRm2+gWpBQHJIfJhu8u0r4wKYUr9/jknWx+tEQEWw8
binNfoPvTxthksOywUsiFE5YWocAEkaIvaMAurIZiETSeDfLEA0RIuca25Q+XaH6
CyrzHzZn8MbRbkzSXHPjfoHe/Lu6iKgElO9avGJus8CCyBlvSLp/EnF/USZ+0wRQ
s19jUY0i4fHcczOpErpRn9hxGHcRTmhNhaTW3Q38uoZAAgFymTZlvrOCyqWAX63N
xokhqVa85f3AiNkyZ3wLe//j0e583M+qINVeVI/cPgB4SHlVtWyssDWVQsRwLdJK
jlo1smoQborb+fGKE33oBRY8anUlqjw/H0ni6X+wUUmEJ8DOaNsybDlNaehmP2VT
t9xtXSLafcnoxK5iQZw7Lk0bGshwtWbedtPrVFMXJStwJ9XPmRSm9UK80V1uYTM3
2YyT0zTNDMtVIzWGFF1bR7dKCMZr5jVu4PyaDbxTe3tGU54XnJuWUHBNdvnURW+D
p0TmT/8wN7TH6jTk8z05dmEaTaypb+/XX6fsNMn6rjNvNHSkOstN8QI24Cn3Lqyn
Q1gd34NtoGxIUvNyz4aQSwOTBiMcr9vRVKHinQcS6CQlVbRhsth6n+7uIC1nnbjn
YRNJizqyDwY8da5iVbCCHzJCf+SNj8VIXQ4uq6XEcztsxXaIQoTfXkX777NA+Y+M
Umtqcbx05zPSCkPihf7t6kMrWM/yj9TjXWs3erfRdlqEnnHAtJv3YK6yK8IMAGCp
d8SSckUeY8I00UJMTnsEWrfysgwwN0UTlfDq+LRuT7Z5aXxXS+42LBMRE5x8b9Gg
XryEddiA0dbfIGxxEehrEWGcRLtLMQImXIJGINZtBmj+I8aOJN2PQepnhkVXvUW5
sEOKeSWK2PWCbGMohU6qeW3dMlXgqlEuMouWazhKmawv0Z2Be0b/Bvpiffzq6z1R
xp+nMwHcr/GzEfoTG+6I2U1UEtgkuCapP5CEcQ6Kmsidyqqt1yJzJNYgYaaw1IVA
1D1HGDENSIyD3zHHeQiXSV6yT96Smz5CjjwfYxpjiRmifukD41cTflAMUhhpdOwN
n9w0eGAjbqQBSzO3NC4o68KN6dWHaGwfII9IeM8GuiDdO3N28iaMHqaQhUoyCBCU
+f9OLabL+KfEJOWT9pEXvYI+b0cXoZsF2sbQZWHJodgfwDcVTHZq+JucdhVLV5kZ
wEov0OPPH8dundpqa0qhR77sYfsnypjjdCljgoAqJ7m86heMb+cb/PNnUHZ0lLc4
z3eNdz7Cgfo0CyKO/Nja/T7srRF/nBVBt2pOFVNvDYJXmOTvprJ4PTM2b6kAa7W1
uNWtYHfrQ/divPfOqwe4aIzxNC27pOpbet8SHk3G9P7neJibv1wHw6f+oYs/dCdA
AvXScQtZH0Tbj7UTlEKf1MKuDWPCZa8UkY5O9/Bd/FID0SMFb5dyyd9RTl7KSJe8
F5g55ECX5D0CBSUu3RDIKrCQVnPgWe95jn2SFjFBtjlkbqno7CAWHUkbZZnaGBYA
pJyvUPa0IbkwRCuLUAkef0ebl4PoXQeiPL5e0wIwvLB0QFS5ztXTAKHDe4JMNl+v
Njf6f+TzR4onYr3GNVbrtDNa94eqVDAPxdo6UXgehiBwJhvcEy/z6D6Nhh+0ZBD7
VU4++vVwg43KtotRpornmNYA49QHNZw3k/Sc2g3vui16DMUE57Us3qQfRyNsngzz
lFNpLRfXm69Og6Pn9D+bmCudJf06frEgCFs+H7y3oezAc7RXu8AsVilLNDmW+Dq0
KIWHR+xjzRjwhSoXbXeJeDLAgYJZkgPlWWLycMBa3DJp56m6/mLJqjDiDPvTkL0X
dEx3mpfUt6FR0usVIFO5g7zm54Hip+aEQjh1eKldZIKXzVJy/EDkSHLFzI7ktgRi
SZ5261tLf/JRLECTlbpC30DP6HGTES4mQaVEW/g/lNn4A7t6s86LA7W2Koibha67
JIvg99HEQG6cgJuXytx1OS2K24y9/lnD/lcweKqu9Sv8khHnJNFkkIQj+l1IAVCo
iIMJHEBZ6qdWBRohorK8j28RYri9XhwF8H9mXX9l+h2B2mPHZ5A2qU3/y9mChOaV
PGn9RSkLSpokJTMtKfP1/An3QmpF3ReVDoYX36GJX3P4RMiJUqfJo2zI1cmL8evQ
5dacs5/Ip37wbRqZi6K8y9snBeM223zWWk0vqeK6vp2HqGkb69GCyd7QydqH1KVm
d8DDyMviCPESssKSzpN0hBtUgW6zaUmgVwloQwZtxqED0Q8F2z0lWokut0CmayMX
kL3uwkb5NommMvGYfej+92lSDR4sPPUYXknOAMCPUsRvO0oPGS2QS1TdWJB7gw9s
t0tdoDR8+MDVwxapdWvWJfOS0zGBJIAqTQdIGFYmvDg0TpI8NdEpFa9VP3UswcLg
UcYd8a61JABppkYImJklyOJq2XrNNPzwu8YXGFqIdhhswX2P+uXtKIkAzrJIGp1A
oS3TuODp4NWuLVUWr6fpaHrIzwjJc841nIa2VjXRBnft8uuLk2XR997GQjXF/KJO
DIkXxRqFNiwLaYlUWLurDLKUq1Y8Gw3QI6bFKT4OgN82c7dSlHSv1lL1FzC9Rgcm
MRItBzccdCNL7NB0W3WaC1eX7T/gWq0D0p4AdtrPg2So6U4aWHuqWfMSKhpo9CKR
AvLgrC7Vfu73mmtGYu+trabN3qPRrvE1jOu9BmEvuRxW1LxL10E7Xm+GqzMUTsd9
3YLgWzw1faNUhCzPpfDCaMGhtqFQVykGAyZH0Lc+scIONk1rEqqPct0XMNQInJja
Vq52Zx4Xp7Y3fn79m59VA262/v6Xx1Zw2SCvJL7qKpm92qCet9ac+FfnAnlFmsHN
WgOlhdoAaAwSgDBH9jkz6BgQza2Gkzs9NWQnMme/6B3k8I9xeJ94mbymXl0AgePu
ujnlmQvwhSiKijwBwF4+UQq6RBl8j/6Mv4xfYMLZK+0DxWiRw2dN1SBlIIE9X04p
kfX6qmvqGJI3gw5JV4ZPEDhaWmlfCLs2B9+Yzf0qwaf9Enas1DAQfnGJ9weIOVMq
eV+MtRu2io6DjYN/q3QyMAe64X2wkcPxGBKSeQ3MDbPi9PYMge48kTzO/U+YyCG0
f9rWVWJBuZ2H6U5hegh97ujS0UymRO7Ka2cpTSoI4sEtJbUfV1EY4sTyWtjTeUvd
763L6r0cFLTH3IZOg5dzftIobK9QcGYaFePfG/7X1KCS3N/IR42NXRUpEJ2EZMmh
Bn7oFAQFEHZdGPWqfHTX083WfDjhWFnmJXuir6jl7gvEMnkdqA26pF+YEGmo/PxT
lyqhFqCS9OXBUb2WByLs6Wbgjd4PzXVqX5xyFZMrButZa0fS7eywqRvjCIJiMR/g
jWMxRZZvX0aNRIBVu5+Jc7THskX5a1qslawCgfRAkcqRGufktnY/qC/ccmR+DVT1
53y0Vf7EzbAmMHV9aSJhWQMU1fbjyK3OB6m6OWlg2XjvjGSVsDKIcMm2Lx0vqbgh
BGW+0/kVjHZqS4/NY4RPxqdIgZ1h3NytAZ26Y8jG5hlRZrlKzN61p/HHi0fTiQVk
GTZ8NNMwuiqqJDw40faN3Dp3vf3Gh8+9i6cPv0/moje8uy1Fp6gWL5DACw+2Mgu9
wENKBa3kpjXc6sJ5yoJAQ5cOQBJwRWjER90CuvcBi9HoAZNRL7jftT0krnl5aAC8
akEkgahmekFhDhvZs5eRvy16odAbDKWEfuty+cnw2r6Lw08dMoTQAxt97LxmlCRw
OqRovGSCnn1W9dzTDRjPDyLgibos4nHmfAAzDxTIbTZW2MD3XzVKJSKeQWHc1wI3
j53/T859a+vQ3y3XWm835ZZtBU6hP+H829A0XrYpM5VKzcCoqyVv+VoUHAO0wIKO
K4k9UpuqapCw6D7ZiPfZRCebFaT7yf6cWHORRbEabuoPRepBwytM6x0+GHep8ciL
vSZ8O97eCHN5SRzv9KkRUI8i9iaoW9ML1ccKcMO88YOrJe3IwPafSMvjUxEjRk+Y
fIUoJFVCB0uYALemWbWGTANSiJRRAwRoAaVUlpIlaKgQzdEOWLCH2cLcpQmMru6e
z5/KfpnVAxbowY0tc5COgihvUpF8fwli8/0FFjeXV+mvm3K4OzU1k8RC29alMIRH
Etg/nSfPrk70g+ViXIfMrgUCfFvzHbTi48rKZ52ML4q3gURXO7xHj6CUdhNJHkM2
355f2tEVke/yh388VaFt1AzvIaL/CjC6QnP1l9UaL5Ksf3oYgSKt3tSeZxsBk0Y6
cJ92r1wRg8tVGFH7rtasRU/NGkm/C9ZDlgUHy3TGJzMz/Qht8b3KiuThK7nYo8ka
rJI+hsO7ZMJmB3g0hiLuUSyMHvIp5ZSX2qKlPXnKJWdA05k3SpQ5IWdBG8sRMSs8
1b5kUTGRjQn9ZuJ2IbTivd9dbIu4Cp4bjvcmhX/1EbWjPMvHHtiyqUartNNefi/n
7l1A+IPvW1LQsbCPTIhISggiW5H51vDNaXmO6R1NpUSmqdNM6U+EVCm9Zbe0zI74
pBoXVaKJKgtiLH+yFupFd5T4T1BEADzTDa98KcNP1YTjUXiathMzXtZEZivZGD+W
BbDST/ibnYAPSnamLfwGSOKHTyOCYgTD3N7A1gBDCkZqhMGv0gUkSPT6TOM/j2wy
QeGiKo26dx4Ayk2Piy30RStI+6bm8iQMfexSXGd379Fpu2RXaJrY6wXYnZl64nt8
xHCAnNBIyLRS4KT9HGd9t4o1FWVijhhphXPwlGuugfg1KSG3g3pj7nyoCCfjnVTD
rOzodgvrhvMQB7ncvS/tRJD3cXmc5ffBfpDpPWBA46cV2dKafF1PVDlVi96ZbGOG
lyZwf/hIkmfAt0SCO9on94je9lSOgac26zyXHnt341ti8JRYoHEFrBY0C+/rIHdx
c/N6lqWdo4pLi9OY+dVqz4pDjZ8I8MAoW5Nbd5GdsvgoUJZf8F9RGEi1vhvZF4q+
j9SVvnWGr1XA+xNiTYLkwrAQeo+az5gLYuD74FZB9WP8NdpbKtEC+yCN2+PfZG5r
qjRzRbfmjxLdy9zfAna+388Z2kkyZ4oarc4no0DfQD3hoUrf8uCIdnL5aqXBiQSU
EYJSj5IMKQGpui6O2kvs9NMweTBwl4VTJyniARUSGouGbD6vW/M4EhiVUA1PbMe4
eNgmUCNOaxs7UAyLkpRWTGbLdZF+UHWdcqSO6dEOgIRx+vgtDaBdHW9xYzwSRBVn
eSil7K3i3JBPvUhZKw9RB74jyR2nuMuxYupLARbSWq805HUP4kY0xvYylMIYfrv9
1OFo2vyrgEN14eL7qLJG3oYCIWcRvTkBfdn3aRMc6OwGenFkkTB7D5pqkZ5AHcmq
ORuPm1UEbWu1MMRbWvdMsjAxKtYePFuPRFhXwPmg5Vm+GSp2jrIRT5XtPA4BVJkW
Ks7EmcNP7lELeyb0vA0OGTa9Z2P9qA6weJdI8Y0wvPk7NoS/4SAlX/YYNs+0T/Za
xFr3wqApeXQeDKSvQeWdj1u+vKDdtYu+BeShSuFqgcdr00ITnAFu/wBzRBzyc/XT
8+sHLO8LPgr2V2iweRNPhdbweuPTJkw7qXoPpOPysnfuqBHMI3VQv4BgPfbTa/e6
JF8oGUrTeyP8P7ZPPiSmuw+vtMtE9uOuZp12YZ+zmSnLahl3Whk/vXrYhbvDBKVt
uc7XRaak0JzwZ4jTV1WWbhz0HeD9a1jjg7aYfzoRcp8txkSgKmdDs/ZUQc0OqyGP
Vdl8kkOS4ofKC5KaBRc50STz7iMlmD5SB4j3MJqGjz1yKeAjWTC0/3gIeX7uOOiY
UeKYUEEaCG9TJJJ5RA2CKCgTOcEwmXMaCQBZRP8EPDihiZkDciOvqwmsDeRdqMDO
bmOrEI3YvJW+dXzXCcQ5pDaiIzhi5K9BxNLdv5inq1fOOicPgv5ldTvxKz0OWGP/
a+8v822bDUu92wdoKgLgxp6Ahlmcyw37eFrZ1Il3eSDRZxxM6yj8awJ+fyawDMW8
K6PIuVaqMO5zy1DkWU/GyvTT7Ioxsc0adGhRh1NRYJr7xRZLAB/yHMHuOHeXI0Ft
hjV1jGfW7N6PIN/8sCBcHjVR3cy+6dUqDLQgrTnJibUzaig7jcOBUvjaxZgwGkqn
AV5PToamplc8ljx720v0sIa7XLCjAtyaIlqvUKTs+TG4UeWuFIrvUxC6/TcVvkIS
ArX3mgRdnpWIm/EZNN8RpduqdTeHR1onKirregBA078ahSIUiK836JZICvwtBlJX
YIf8ENS4n6Cyks4Q6T3xVVSi3nEWzslLVONc2H4OV32dBNli0DRKbJA0IzCr/Yf7
9dbPpz+4Rzm8A8mU1sNvIiz0uWJBBZhk3zXHmpCOHZ5fMFk8U1xVRfUsGiZCqEzW
10lnXc8NA48t1t75FdWepV+KacsGkHbAaovtzSA1ifanjK3P4ZGEv37GbJ9NXDbs
lEfgOF5B9ARnkQ1dz/FneVZm5hAYdajekKfuNgg/d37gGW3UelmW3H0+6myWW5hB
bTwLxKK8geWmxZara/HVj3W/BFq9AmUPSOFv0YSHcYVlFllrhKtRddhSbeEwudEf
Wz1e966HIa3mjANF21wh8rksZBMAZfDsz+mxPiJACa42IrQJt4ju3okbXcg/GhvS
uvixGJiAg8SqE5IsQdX8eLKUcw29jkAaVaFfk8HNpacecyusB/JjxG0OqCom8lb5
EV6eFoGrD6u0vLR2uZobmJ4JaO62cUJfxf+c5Qbs31BH7U8dFRxRptwYe9A2Dvp+
31A+xuIiZwUV8137tTQ4SozPcEQUiPFoac/aF9gG8B67weVDkYhLefB//pifIxAz
do6bV3DDQuJj3a4pHx3UPCTGajC6RUNGNd9LL50S/MsatAI5Fm4k7XmdVMtifHPf
Eae/BJnzwAUBWbUIWNtX8Td9HrrQJ3DsMQFB0bE/YEve6YcXAQAhITQWyHfJrjpv
Dhce9iFTDGp1DcxNPzQ4bDRus/JxWYm1eI6MlZGsQRPk1hzBycqm6Yy3ANFbFcCJ
oeW5owQoKdzLSDWKRs3xyzGtma+/dbeE+UQX/CDKryNxDcuDUCBnMsVc6aIfctsj
maV9hRVp7AODCoyL/HS8lICR4QMeqU5FVkZKHcAMXd7ltsoMbY/MJJJ0l+qNZ0Uj
qhgS8SvCTepYbhDPUTR8ZAsAFWGOEo7O/gDyjzo4HTPMBvUDSvDpTWEnlPfkilab
1oqpb+MlkXWrvZ6aLxzWkOrXFPooBwPECAMUiisXGDLAHjvgpTZvkf7BUbI8O8eE
iG+jkqu6cXPL3wsvUhwcdILcWZir7ZKNuTgW2eWeVByHDyQhwrtjlJDwtlIB2Ntr
MtCaMJ5ugRXIqIZDmgZ8yJlTGRLm1z6W9sRpWKdi9TO3LFJMJ7kd9INnoQ6KGNcN
jidQI6+08CkAnwhuu6NJIJeug1dMVGWHc3R+Ta96B8kXyPCZWLAwQLdOV3z55BXY
BXOTX/LwM2ftu+GQOzal0jgMlKjVxQxEYO0L+vFIHQjNdcJbfrBoz4fn0nDvxAA4
7M657ZUBxZEP+nWBwcVljwelYfsesjetmVCcwrNNxg0AxOwslk/jWqCywndQdnz0
wqw7ZHi4itHSmYS+ENNuWunSWjJPaxoHXZ6D0tptjRWnZ9ni7H7DCt7xt5SOz8OW
C1I/YJsqr78QQfmM6ZdiS2gQHDIL4vL4ZsdB5v7mpkGGumQmvbIkKF5hQpxySbZF
HlKKvJuAWMlOfdRFo0i1QtOmWK5dqYwSab5Qg4D25hrErukvZM4jdqm2U6GbCNlX
kyKtqIeoMiyKnS1ZZ6kvGWbebp212KDyYvuIG6pB8BOUJWrMn5/g9aqPyqP2LzcL
JryoXGEA+lVICAJW7+VyhjJI2PJbL02mnd7OmmuoQNNirpy+dVSrl3QR1Pn4Odw3
C7zhmqoh3UJGguKR75DhtnBw5qCkCbrq53yvUNLaIoqcJXgp6Q78GCDBoBtl69ca
pAqmB4cvkBAs7csQ2ZJTRWKVu0fkKFQmAyT7dZQwci0m4NJ5EJUR8xVatdvwK7yf
BsbbF1a1M7XLoZpywxyJ/D67EF7Z1q39yZCuWtI+rcQOGwBEbLfhyHiJBOOJJWub
0hAbR1k/GvrhHttvsVOFJtdU9tdxKWQxPW85U1m2VVjewjSnuxR1APL8gOGlHs3j
XYXfBT2jq0Iy3M8jeG8iKYz/5Bq6Xc0jJkxRkB3zteloQtd8jmP/8K/RKdAHpwWC
EmK6J3hj1yMs4HwKbXwpbLZOj2dyTalsyGjNanvD8nfL9ZlVgPEidNGgif7Y0Isc
nD3ayUG1pXyKvGNb5J38UDpFEa92dR8XW/gC+7pI/FkdtFu8AYS3lo/hSfBrj9Ce
yAiUSlmWppw7mcsk8SaRNt0LvCA7t/Y0RPWrRHHXr/iR4kEBSZGoioFQ5qlSe/aE
g7fadbIvaSVsSjxxKCyitkRwvsup+7F2Ui3BVMYxi5Fvz/E/E0z1GlhILP9uTjVE
wtNze/tthxN/Qx1emj7r2NrhamnA4xORmTBRW38xQZH5I5H9sVb+r2ODhEFKAtqc
tw5r7vhZpywvAT2LPtaFQ7INQY2MqqIxM0xmhdoGbutpupUBwCmn7xSM4qgci13t
EPl1KCmAw95bqs8jMfj06iToOqc3QZ33WJoBdQXc0NlfTxuCRtMPREi0B/HBhVcs
oMAyFhkuHOAFkDRuDOUDMj6xU5tkbe7SQWQ0hxPyvx3or+2ZIOShV0lBzUv5u5lU
rIzL+tPwzN+XomF2ouNNm4ECFl2Ho2q/Wwa37yUvk3nRzfdhej6AyDQrX/0HYgAN
keuFrTNSxrDY+2sFWuAkWrd2qfF32XlKHAPIrByurELyNSgD/K1MeKQk0RdUoSc5
3e6NZMdMMmN/LlYqteSXRJjFH1ZL2csyEjftwB2sfqUDaOCHQI/fvQRyLZWdPCfF
arlkj57uK0HNtQL2B+GzJUvHNFlHC5uNdgXJgNoXQT7OA2KfH7VHwlm6afCWW4gg
itZN6iixNZ1UjsxhVSHQ4uYHCERjtt4IXjGs569IypGZUG/dpMaFpPe0Mjuuxmjo
XGIuRTYeSsCQAXMcR84B/+AxESGFVVaR2P1jE0keob01qN0g7UmKFawJ7BVDlUMe
tMCiZ5T72cgouDy/rGYOlna8w4GFQoq3O2RIxIsEFMcrfQbYxW/YA6c6sELl+Al2
qZKvIwvbBj6SZfHQLz0OJ6rm3sKDzHdr25TgvZERPI4j8Am8Xv/zAYZJEIMiuv7l
1/auVLfs5j7k82BOtm+CyMLFm6PcENNMvvhapNgG3O17djTEpMtpH1h6zqAm665G
5SfkrUUckXaB5Ypm8X1gVVT+xSBccfAiMTjT0jMFv1R9Wt/404GBz43/P2BsyhRJ
eR4POOWCZDhoZohP05pNmR2J7TjnfrfFXl/0Sm7L2LISkKjSsfrMMyRpLu3q+YzQ
WsyTHsEWEYxotaxoWiNgqwq+4XR1E9zGqYG42xPrsDUVjHTKHA+qvHXaMGrGZ5Mn
rttigCxLvvRTSIBqKCh5QNHq+C4nUHrrxA0ZnBJrwZ0HsvxupDFrcJFejBMpjydA
/J5fvc7D4U/1xJ43wf12IhwIzkZwZQerEa61a8HNbKrbM4mmIKtR7ZnBkCb9aynK
8rGuZb2xRwTRnbKjLA8D2/l0vlQt2mDZOs1a45zWF6BcRs3MwHuWj3PsIfDHtmrg
uFnVDDM31nEyKEifFwDvIrONofFkSKDnOZ+wxpZcfAkHMlaty4AVPGYHFCXfShZo
GNfI6U2dOVQ0kZcmEtLqeU7X2Xy5KPWSCUy2nygrwh0wuSpJg46+TnbQlxvoOT7D
SsGoq0w847kc+k0ZZ2QYKcTLVPb7jrDUHiYGmmCKd2oAUywLca9FwvRFSWqKikBe
0SBYIxZr0ILJgv+89AizlbT3vs4gW8oIp+Gt6RLS5141FNNXXd+Jeo4uPaKwTZBN
P5wb/rkabW1LeKvQkeAXoLCUjt8HEJ0yunTtvtRZjgoEQZ1Tl1qZEJP0NzjiwPVU
+6EY5FQOHUz1aBKY3pmm5IOnoKnSfTFHvIfdJHlNciZOYp3FdZ/e18pcZZefzO5D
9yP7fWdnz2+tWZf66wYg6LoRpOTlsnr+EXOyjsAV6E20l1qPQubC48MIZHAK7ca5
ZJVWcWhixjck2ihladbqFURd4+H5lPpNjB8L3He/RgXXHmJPZrJ2DPQch4ilsjZS
2V15txdfpliC/v2k1vBu22dPX9/x9ibGM5XaTfXCNAWTMaqgyh1C5kOHMtqin1pl
GbVupR5z341MLajkTxwVv4PNyy0aaiLy0TVKJIyjAP1NKGm37MNLJUsaKReJ0jEV
9cQFB7DYr4DIDkBXn/DC7b+RG3R94g9rdT5K7ktkxc8NBUt6qnBoZuzlhHCshYrb
mmEOIbn4/C/q3xn6Desybczjee8mXo43aaZNrEjaEWF2oQ7xNex/MUJF2E7qcAGR
ic5p3/vV/uYPr0VqKbPqHZqo+3zP7rwsKZwpX/kY9BwI1a2OatLyL9m02jyideeM
eVIcsMku+wS5Juh49cZ8wpMQ2qV0pr4JVhFU9pC0JFjOR8i0T+AMh/0YtW/V33Hm
JjaHhSIsh48I8hG1HsErT2Rsh4CbayJYeXLiX9MVYpHGlzMaB7JT3ae4LXkZiNMU
WfD7aAeamDaW6ZvOJMoEhZHekMhCAM9LAyLXZbenL19RFz31ituIDk3LAmOPTIhH
bi7CLJC4X+Q6WLFYZ4AG6UACuDZRPDWHcy0vkrdOMmtox7yXpYbIedUzupMLE6It
OvJgLHie4TY8NcI65ZKhM8aIEeXOqhLmcqEgunw6xBkygwK05wD8EvPx52DMbP4o
Gzozwh1wf6vQP3yYaCtJWh4Dye4NIObxXgha+UWQkNNRcf/1E6maXB4iD/MS7QZa
jdfWY0bcBFUkwhMaLj+qVhAEp3Uw8cjFs5CkDOdSwbyQyrNJ6SN7UHwZcm1PChDS
xpvW97eNcuyhMstxfnzg5btvsu3/h4yfQc+1zRUMY7PQGRK7h1KooHEeOaXm6wc2
6z1SutMseBEvjHYGZwAhxg1Llmft5yJENwvZUVIVLlZK01tCXhgJ0Mfzpo4JWSTm
2ybT74CrEmEU951lBVhU8cAXWYyBR0sl69wAtPSpoMyLXb5LfV+kMJxgAOewhy/1
ndm/VsjdtAv2Cg31LTXDZvAlL+o9taFrAVKCBf92OFbehP/2TT7UxA9CWJo8wxU4
NrwhAU6r6Dzbcfr3ws+8NctzAgpCpSx8uCjPvgdPKQyDwrYKW8MwnNbQyyrQLugN
bCpr8eNRAWp2vfOcLcHq1q8u1XUaFtVNZ54t2t6OPeLGCzeKR0ll6oJg0Z8eAeKD
OMouZPbigoQoIL8XFJrtJTTafL+fmnHePidB4hZDDfAv5WFrhGYVsI5lnwsDD8KV
Fq7lHSmMlVIDhF+NU1FapLBP/LVRG9R6NWW/jN89sJKkFNYGzEY5j2gPJxun0rR/
jH16XVhu7KdjNI7edgT5Yl3L1L7wdFnv6tC24A6IsKUVkKPSXw+nDX7omUFnzLGN
MuWE1H6Q9HDQiFim4s6sD29qMsps52qouzDkpw5NUtpGNH05wYCmu0KEj7i3f5OD
l24s3/qHZM6tqhC5M1VZwbNWOW97DfvyhzNg7XkKL57gZcP56hdhIB9+StXjVLhe
W7pjxAB5BgMfiE2cWynUDu3rq4SXWzKEWdyBKVq3aRekNJExtMLWAbCqDxXYFNPp
qiCB6HYwNAi64uRXteXKGWedoPgRFMJzcO5Hb3EipO4zH/2Cf8gvNwYXwJv7ftPg
Dz5lmCzzX1zsRt0NJuPSJO8GSIHxjTBd69G7EK/73uQ8+yKyQpYroxMBIQ87mZIO
GNlaz1BrwvBNoSq3jXfjKAZnUGEAcew6nV5OiQf0kNHt2jOFSNdqo+7MXk+Dyw6W
7qwSmBBXCUdjYWF0sMGmY0lX363OHguvyiNPLA+HmPRIK2S708mj/zqeYdC9YPF0
6fKNgjdc83Nr0hN8/23/97PGHWhtFnY5yBrKo7cXpZC2WV++AG3o8CU3XntMDsLw
1wADvGTg8nhBo5mrxgYhiPHeghvodek39YkZO7bGXlxzKfAEDdImVWg9cxiiaZzi
Bs0MJEGpRayH/rggrNhibRoLuUZoDypZAPeWcYBaBnsQYGR6gCyqEc/m99BqlIZ3
bf9s52AKXdXFhfnw/ATwklY8YtQJ34ZG5lfOCkFGU0GZc3f4G1m8m1YQXGANVrhA
2QoISg2DGWaQyPFrdqMCscqhCCmW/fc998/YD6j0BPhLuttseLeL6Bf3FdQkQhmJ
x/kopHeO40fUrM+hdJ+dspjT9SCRfWZ3TFY12d/FKiA=
`protect end_protected