`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 4624 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/9huKRhRMtvnNqb3Z+UU7TahEoHV+T8U3P3ufru7l1O
3DlgtZzb9QxCbOjthp9+wDkjygH0eUfDrEl1ovhZG6006P0iV5mmYxfFOkqu8mfN
aHoGdj0YkUAaeQ7O4AzMRpfjdL+cjbnnFXyeTxfRs353M/Q4jSyo9/UJn0WboxBF
wt736DxKsuhoYvuj5t51JXOYy1Xrct2IueuRTrJe8wI2jTKbPBwmaY4udY9KAqK0
/5k7U74zAtw+BJeLIAzTeFzDr4vf2Faa8in/QkK/14jiMI2CjZS/jYEuaoV61owL
nd1NcNbQ4awLsKBeaTaVRPBBsVaLb0+ONieP3gKSAn4exoaFxsqc0jvAHQiN89YA
fgVPtt4XCjRf9YdkuFQ4fADj9rwanbWBpr6mFcAlvCoPYZAmAvJx9W5YpLS5kmMY
Q8zF5Ly5yLnxava35VIQoR+rkAVESLBlBSaUQ+HaXXRBxgItRlc5xGaR5u0QrSq7
dLMCwW4oDleP1sQEYYWdWoJ/NbX374Ow7xcrYNQgEEPr6mZ+nf9gWkHaW276wTRx
qOig7qMTnAqwx14pCqv9Ba9UymqHDWWhUhZmn7tBpnJwUyTUNAldjHUF1F3jCUbV
wwM0MLaPHTEL5Uzba9Go58fhC/DMrfaLLvIUeC8ZpQTAMVcp7aVsoIz0SGETpC1P
x3Pjvv0j49fP3qdN+vi1C0FiVvyWOEEEOx9yomCJ5vaWz+pUgESINxb5L7tfo6we
559LATN/i6Qch3DAufiUdpKYMZmvkGQUzFq+zFoMXxPvK6UfK3k7EXwRW4kdOmbF
7moqpLR7YZ6wvIniMEXJfhW2NQxKMXmg+sy3mUHd87Okjbovrx4R6AU9eor/CDMg
uJbKYd64c0fK0LJSobaHehoMmrNJPdooepbCNApgzg6jeywckHrocy3Tn+/Zlq8Q
UGCifKFQGVTgAL13namy4DQEup/GlI9dHjvRiLexv+tq5zWhIlu4kqTT3n9GrNdV
WCFclW9WdKqhoDoBhcQzljN8hI2UDUGhfsUyufgMZG/PjoYjaltcJrN8ZimP05Gd
mnNL2bGO5/8jyEyLuwuzGmrTgLwGy3KAWCn+nab3T9fXIsu+EaySuBcbZqnzNIrn
EOVxo1yb2TzKVQ7zM/13H1ILpd4qjxj6kuWlz7p6W34eSc0gZKsAmWwzcD1N7kLo
G0UaHEih8o+anTOCrxmM9+vbbMX4YjfjINz4IcAjVKkfPg/bsllibCagVDQ0ZDoA
LSM4Gw5xTugCnuIMvGSTbr4Y0ruj31R7hYvwMssukaF/FMpfTnye5oHpSxVHYZp1
Ttdkq0tykvs34v30gKmzgZuw0j7b0GD9yevc5DLTzf69evmOfIkFca9e0lZd69EF
ZWwScL26REG0F85GXUpuCihgiclw9u+R291juUwIOLmNxVJ6g8ip7IoBwp4V+m3K
zFYEZntM1fb+ynZJ+yi+N/nFfbiIb7/h1Y8wIynHnLe0bmbnA5stQI2dGpKMNpni
TUWv1mgHCtaBO/l3V0ldgLYC8hz1E6Ux3EuhkSq9QbGJHILXDlvBACaiLXuvF2IE
AM3gdlYuqDSYB3CXkzIagflQsmIRqjomqUvOwJkOVPjy/nS1q7MUS9ZjDid6p0hO
dR3tEZIMpdnWAP0pT3+KMT0dnTDBsaPJII2pLei/GABzikq9c21dIjks9Dbpbytt
8JPEyFMiBAxHONKQ8PEN3UtnmWMWx1FoQMoJqZOWBCvV/pcQuYhBgjerPR6lGi6J
cp/leVebo54cJLnczaJ3waNt2rmXAJFikruwd5Tb0kmpCpjHiHYFmEr0dk82k+xm
8NQTj2/RNarPvaGpzpEM2vmIv02nHT36NhIkRoaYBXzUN0/jt1d+3igkZckbo945
stZ1JQxrFaVBEybSkayK2dH15MVoGpJyko3SMCN7O7pFQtPeQJRLYeO3T5dlNWx2
HLiyHLNhtiKy4MBuL1i82KkdfZHtHak19RnioFEc1NvypDzKrDAWUb9oHcG9qU3J
37jiaP7pHDCwWi8OI85VxOcAPoBEC+ZIRqeCIbM3sVPWaMFLC1wq3OwK7CE73Qj+
55QBNOWwCltDVG3rZH0WgE8SffZUVTLhC19QqwPa65hn+TRYBZHx/BLdMNApayUN
W8S5fGOGDu39n3Owp37UWpMzdtlv4KMdXyYJuzHESPflBHfBDO5j5NqDrSo87pVw
1H2HVieotf2SH0aB6IqDk8orLdRTmuT3F6faqr9qSjSYkQQDKDQhWoW9NT+r7LCx
2ZTGamkWmyWf7Ks4O34z1kKxuaLpZfvw2GWImgAq/Q+Xx6Zk4+vSvhGggNtLIGSo
oBJ61k1Fgy8dW1hJnVpDh+aEJk56l6htUd8qTH4Sf2zbN58Yql5412aqVy/jWYYB
EpjAQ+kl5I0cqA08xLngUOgxjqm2A1q4DI2P1k1/eLcbTux2SwABkIvJInBfAUSe
MmCPXXJBNdCofIvKrYq4QQKnQyXTkK5/3JwQM7WGhjYc1Mc00JrQB0pw6mWaWhqp
mlPcLy3Vt84LQgYD+t/AeHJtE1SaAbnG6l47noXtZ6/228uNELCFFBj8F/T0cjjk
bo02q3a9xwpAUvVH7XkqWQJm7qmsgGrQNOVTWGwhkY9XHP18EV1GC455nWcGAjyv
RSoX/wY3FwJqXU6lYFQlTutn3DEGNqRKLLYlGQKUTcgSlX7Qk3D6txMbiDWGxaee
YnbTyenLeWDKwZIcR3cx2oLxEGTVEH70tk6NaUCo8Ch5W/nMVK2aqojeoH1VWc+P
QFrkZEP0NBVQS8fRZjrozC+05gIxu2NRyR0WSdK+SyWcWx01OTjlzQct/DK9dSAq
yQwW1DAT1c9uOtAfURNVdc6Fa7UhlbVTDeUzIYGCEdHzja5a1M7EVoYzNgO4S9C9
dO6WGMeJT/IXhOC35b5SjLq4KCV18jjv7M3dk+3bWPzee2n1rx6+Zf5GAq8U3JX4
CumHWoylXQBmI24zI/bplGwRGTSrK7kyJmnsr5pTmlUf5tGFNgtHDiJm+lia2hIZ
BhX9I46SRVk4D1uMK+QuolOGjnlvrM9uXovtuTSsOPYSOqor/iYPWY8wg7z2VUXK
QegSxchXRTVm5IwJfyYCRT7q3a/AxQdk9irYiL9/rVHft5fp9tiiq+2XgJvikrrF
r7yaPsqcdUGtxgnjDa1PU31ZzKDFCg1x0/5Yy/gmsY/Y8pLDx5Ch6HKYed4vFxhd
ijcWJcL2h539dhFu6rb7g9LUVUfNA43LFFLst972E1SsRlr+8fR91ZGS8Nppf1c7
Y2CVfVt27lpjkisOg4179dRfO6OQxU6/D++AotHA2Hbf0JOa+ZLoD2zRtSve5MQG
kbBnj/aXLIeLiaamO+TJzNGiqWdqaMrTYVa2CmenUFUPHT2BhJ7abwVw+mPUjCaU
xENBTegbH6vdx/hgsdxFSyA20xir9IG2JTCjEs1WC5gULfFbPl1cRpNXKn6XgUYy
+MKeXSdDq+Dr9mbZd6kirN5o6NtcNLcY5/1hEn4k3UJnLf4qgArc8xZn82Lr3szT
UoLi/2ZgGQCWjKFiIhwZVC/enw4FXNg5HReZmzFCsrvRXUxPej49dJZAXxnvp6GA
eJdKEso2SWEUY7HK82zi/a5hvzbrStPIQ0lwEE2BBVMaG+6ahvaSnJcXFYS2MrFv
UzTCJniqKsMzScETo8nLwaLuDUZgw2krStipnLB6CcWc77rgqypnf9aKub9ja3fw
dUgZJjSVjDEL0HwwikhY96K7M+UdwRyt0nbmQ0D5qlYaqVjK43qAJLjCYxIXyp+w
dyXyUef5ykqN1gMAfRpwTWo4vylrocFVGTe8yelzNALd4ctxT5Xc70j9rcG9ENkT
3ZnHFbztKGr43KesIxs0ALjQOPN1DWNNQhsyp/LItoB2RkvcvsiPrRxFXNPwnkqh
rgA6s1pQYIdG88RuxjiDxfsR/VKGvKTIZajS8EL5pAPYUiccSIXvjnpxk10UUYcL
MRnqFZP8GbkCapllA3aq+nKNiPD+PKxiCC3RDLQJbp6zjcUgw/2Su8ItHo7IYXnP
c8flLkToNXD0gkLxWOhE039BR5Suhs6BJv/KU3ESEwPvC/UqIpMn3kWQdmBxQNaD
o8yCJgZ6dC/AMSJMLR4dguiGAxPaNpqXxHHNTcbOiCx/Jui10ZTQb09votUN1N2+
o3CARhbJ+E+nnLmcfJR2ZIkfPBx7ejnyCUXTyAgVJYBZ7XrsQRI1EM/yM9oq2NU4
5JQ0zH6f7fdf86e5aCdca5mAMXY+aoTohDFkeA7U/sRXnvE4yVy3BPUoyAJDQCWW
PfKrh0yTUtn1w0gqXTp4Hn5GCUJODQ4I9ymvs9bgV+nDe+davDIbGldqYKxCPuws
TZnGCtZfI3mWPsjiemYbsw7w3SbLVZ9SzxcUbCABerkn9l3CTHw6emIM80r65uu7
sfGUTdqkOSQ5uyx4c+YNe7UGN7Ka2Zx4tAq06dBwp7M3iJv0bqf1+nGLMO3MMlj5
R1ukL6jUfO6dZShL4vsk67cre5kHXIzxFeF6gNHJXmDTHPQ5wDsWOmW5ngx/e+/y
xerSwXI/zun+ROhhSVxifLYRcCL94xxtBar7x45htD5UnsY50iVN7RiusI1laA63
XLDg+dhS2CpxB/ngBJG0FCdDH29dWc1+NL4OjLKvJxn4MW0BMAQUvM0L43xjfQHU
Ubc7oXX2DQyw6ipxCCNVBvL+dfdfa4DJM50gcgFn4HWqB+avGMHuuRQok1o/XQ6n
E0on7/Ouu1X1WMtfJxkhAvtmLnvJxUdaqdyWJ+wBQmtQW1NPESY3gJp93ezfBpSp
cVaTNKnB81x5TqC+SE3trd97CwJov9AfeOycw7brMAlHd1us6ng1GCUb0WnZtdeN
2zQCSefXLo3zkArJO30R6xz6NZ0/kJ0+7ZvJEoMZLnSG54vdsFOw7atKkpqa1RQl
pZ3BUnfaaugK+T7qYuqFmVgvN29sumXMEweXKoEMOmG4Mosm5XLSYT6FM4jNuSms
70U42YriohZ/sQZ7SGwgOWPi2KWLAZtTgvun5+EVGtevY51NOh0wGE6A4WwpdA54
5PDGCRGBhDHOYFA7KzZagKixh+6AKX36jSBMKduDmFYOdSqqhOEU5kjCwHE9vvJN
hZKW9KFM0k7tuVGBtzDXrSNcdINZ7h32UT4SvQhl5dyMA/+Z1ML70t2jndOZGdee
1pNDB132moLSjN2dwmMO3oz8dEMFUFFVkqKW6vWy4dsXHyeiGJEY8ba+Q2mcRJH8
ivfLNyacaQelwjw4bYrnw+NDHuf8lyLqwRhkJe73OVXTBmES9gfo9sv/ORi7tx2M
78XyQH63vVr15g4x7CCbMBWcG98LyfU+NcY55vuRcbN0jsBTEQHvSmkP+ikLErl2
JSW6MQQUwEJ4NXufiXiXBEBeaTDINK3qLbonrHdHkOyWUhT1CVq5/FIUA2fNJcxP
fk6VXBaWeIa9b2OwuG63gsQU5Ct+KmK3kgnHrIzN/42UYvQFlz9Et8qWNuOTuESt
rhRFgl1JSon0xM722amaXNfJ+yZ0l1Udo1vmJjGArTEAXdT1ZpfAec/h2yfemlcV
8ErZKucRI2Oy4OblHhASZsoynNrYDigAZX4qgwlacnK9fN5tBVI4V9vZ/qGSf1uR
02/CqKpJ++AyOOi3vvomq7a93IaRMj5RTMSqdGt2BJeOtG+j+8Sq3obiVgrx29Kp
eebiHWRIwNHByRiOHImE3vTtkg9w6C/pUvTw1MH5ivRoyAhEtx/9Ph0Saw4+Q0fZ
ci1vPc8ntfx7fVvnzx3qqMSyL8iDz//x52sxWIt6SzHytxD98gN7yGHLOQ4DMEH1
UKWxF+eAj37hcDmdVhiFbWj/RMXoyeTJpQr2WnUDYqTwf8qgjFSiPCm5UCu2YZMb
SRizMALYJmlKDsq+yxNF3qZ9DWGb2fJ+ldbxTE3cZWOHqgKN8g75/NkpM1+UpctO
IXlRJet14RdV4aIH0tL5rBbREYNXsc/MN+5/NDSxyXqpXYyLo4HxIPhWRN06mqgX
FLgIECt3oQXjFcZPmIMQxVhBw6BXxHd3dNkdrrmo2Ywr07N6x9oMApRfnOOlw7A6
v6DqKp7rW7W1C551YE04HA==
`protect end_protected