`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 4160 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/9huKRhRMtvnNqb3Z+UU7TahEoHV+T8U3P3ufru7l1O
3DlgtZzb9QxCbOjthp9+wDkjygH0eUfDrEl1ovhZG63owkcFKKSIxnvlMdDpHe44
QuOadcbQaGMuVBJjnCsa6eG61iVFho2rwhM6DHyDpE/Yy0TGQi29X5OZd6Biw+rG
Jadby9JblIN3GKEeUauvJ1x2Ls+KZsLJxhmvV9o6t7pqfRntsKCan2mPwsgztsh1
ZUpx5zZvvcZuaLJnMRnIZpybYx8RXEJDSK1lAqMupro+s796ueVhd6g+hra3kuGo
rXv1c+ObRJChGuj3/VKea65PTDLfSPxtcaxTCvPUvJCLmgxAI7asELE52kvHKZQ6
DmcIuk7Zf99u1zaxLM8vXjuFgL/hqqB/ZIf3Wob+27dZZ5oJESwkmiVc+Cz9+eK/
qGVNYJ35HLkV254ztbUluUlNTuOyDv/vFmOWQLVjx8b6zHq+x3siVpuWerp4kJXo
d79NHglZes7BOb3ZXG9YTw3LxQntdwcx68SjiQe5W+SatiV6xl2Vy1ZS5+gfI+lz
mXiehAuxgOhsjJhgpqN47MZxr/ccsQ37r3TcqHtcIIX8+BJN3SOjgF1geLgG3FDo
UXkWTdLVfZvO865i6kS+WA6yZK7spNw20Fkw0567P6HWwiZeiTDN/SSG2ViKnAOC
N0sO06Yf3mHEdDqCNe0oqmyVxOCZ/6pE8TF7TlJPYfpQgTgDXjz3ibpZqcFOnw2L
DsxAzYtHuNz2yunam4MFt+lNys5PIimUvA1P7mmY2z4JJ5tgyj6YPEY3VTYCzKhm
NUdIHi67QCTUpTJ9MKORKib3m88TqS/OJ+6MQEe5fpLbpIqsN25CKx2agJVrsRqu
dt+9iJPPXcRDyTXJmMVlZHvkmnk0RrTF82VX5qn8+3caQ6p22Qe9MIA4OHVWSj10
pBcf1Urn4/ebX/jBIF9c+8hEDjZbmhQLMnJs47RCfx3SdmC5t/MLHeWJ+l+Eb7xp
mABb5T4yFh3bDMRrtrWlumdFHZU4RCgdTz3Ukzyp+wxWoyklbjmprihXrC5E6wWv
/viv7YW9nZFbGTObusWGkqrWk/FSFBeHH4lHXSEBzpL6dyzXeP0BoGLZtUf50wni
oXhdwVJI2BUtrvzdUaL8mdY6VqM6E8U+VX1ej1HfxyO0FCisHf+l8CABkfxzACSA
L2j1X4SPlUDJxNyhiJmmveSnvkpOvIVxpv3iW0+z+UpebgGjYsbhc1f8cs7Tb/hS
MAwGQgeJNfggOdEUq3EPb+T3GQkMmoXPDrymSVsKJw9CeSL1l115LZyiDmTJkUUD
uS9GIo0Vk/blAibcwNOLnzc1+YmILDUA5kygEz2vEQCqK1oMSBts3edIPvB9uXGx
9cMQxlcUQ/VgkzzvrhWwdvk6vqFvc6hzx4audrpL7idII09gJC8Z2gbieGIBV4WI
HJAkShRe6m7tP+83tsr0ld97HKbv+oPSyETbs+eHZkscD3kMup28nLD4He6iJU7q
GNuxlwOnfsWXXZrOnyXI8P9NDImRFkNKWE+NouQoRBQsbvWOwzrtW83AlUxI+TCD
+Z17we6u0GVaiq3w7/V4cXG3wjqqTmk+2JOHEQClM+XkJZ0hZsR4toQZemxvht74
MwbnQT4YiZa8f54SsGePXrap5bB3/RN4sfKzZJdv/uifuBUYeL66vfkkd+XHucpW
QJTP7UpBdEqbKC5hdP7s1BnVL87OJw8SfNVyxiOl4j+lq5lsDoMZzWUPiTdIfC6I
LboV3gMX3VeR1wbWlzfdFOJTO6Acp1MHPQ4th6tclPz/1p+DFO2bOOZP+uUX36aN
JswY3FmQCOCC4pRpVNgpB0eYk6QPsBsmXOolbM3OCD50pVq/6urFELkRq8Wf2MFd
nWSgO3WvBPMUZAtCaPr9ajTe2TNIWz5y97UFBwy9D/vPndlgV3NJ39yluXFZlWcw
BDq8BxXeOCCo51sfdBr5uTjGdxPTGPtTA7yqPPF0noeVCwvWD6QHWtA29tSh/Wef
JuSJGllckkLpe5TwIxxW1A6kn7hEyD5r+bp3DaLNw2mnNe1v/meuGCMV+IbAPCbv
TQsLXAl9cxEN4APG1LkKw17GUngFYGhgVD668oPNSrsqb7qJ0IM9qZFQ4iwkuUNX
uSIArRbJgr04O7Zyw01Gj0/ahTAS9CM5u7lOYJc7R1oYlf8E/yFDHEMXm+D8dto7
9XWR+69ABewOja7jziNy21tSRFQCqBfQRttFUn7BqrRUHMWM7VjFXZdOloKW3FAy
ZGH7DRIiSLcupzHiMJGNQA134VuKpIigeeqFERddTbsF7qzXJtshSIq2S7Aj2KA2
1Bj1dSwzgaqREulvVUHkG6k9JzqDMR9Pg0BtsoyHd9EmS0NqUE5fypNzEh4TDMQz
uJfeLVCs4NQlJy8esdpetx7sE/282/GIR7fNmFOMXfeSYDb9ZJKcbVc+K8ypaJRB
3YCOLKenSE1a0BL9Rm+TcvT3enO7URh7U6YMFwHJlfu3Ga+0mu+rlRFLy3qGtu+x
NZ5J6dwUeqDJt1GRyzaSUgHvmElyHXvTRlYfB+CjbWs3Pc1DrvG0jzCceqcvePr2
80r24qeWEnKqQ7/HLJ0FPZze5IK/8dmtdqkDqbIrQaRHv2B18WAqLTN+RRP5z714
rqPwNisnd+l/qqlOn6veMuoKWCVNRGi6twp5k4sagQHWjT+YvRtW9rMsakdJPpMk
hFkGYCYLevQ0CZR2uPNp3L5CPEjubA39G9f1XLLrKQ96FPIRwWEeKvtKKAy46BsA
s/EBtF2Vzg82gC811yLs1Q5GQbZdpFXbXlwC87LngXniKnqnlUei1lmiyLRJtCE9
2PCUxDAxTRNIQom3cvMcHtZiNWLkZ6yna28FyzzUFv3rIi7PJ4wjFXNK6O7JKoqG
2SJrcBG4yaDhu9HzOL8d/bG76YPgbnKyb9K8L8FxoBmkGMF9tsDD3+xu8HozQeAf
38ONqxMvA06gNAoW0cmAjU2HowEsG/vBmY3qzVWkPfQ7KpLrWn1eIIhDZZkV8eVc
6E4lhHFn9YycOY5wK4wYTuMKagU5ttfw6XUCw71flbzC+8nx6hYFX/7dKlVs66qF
GfAYmS2cxl6R/8P76n5c3i51cZg2K+ajbZ6etK8yjy0CgnWGevD6ssuwvC6FAtdz
FO6rIjDGN6ttKc+fF/d881d5upe89471jiKBu7Phe7Kom3qql2hIeM/JLku5Rtaz
WKSHwgEEM9VzgEdwqCdejGBPsigsCJNg9e6/g9KsvU8JZxwAg29qllkh9ABg9Tmp
IRhFCCEGbPpsc0Vm3d0eXsRskw3QM4+ZPM5eadItPtzDtz+9t1FhrnXSFNBW6M+7
MJR2Gp/YVGVV2Xmz1IvEkSqh+MLWrtvkB723r4sHUKHrzODfIDFZoRKxVXdVyUcl
nk/mQRwLnMIKA3fhfuF9A6nBksjgEveb8tDzIDW47ITeqOABtGLyUDVg173vL/QT
hAEdK+LHBXkSCt1zw2BNEGbqC9P4BiyVaiqaqETmZkB99Ua8ORG6mnRFsps2TSta
9kdgVfhHLGJkyLGglDRlgwPB81Gd6kcNI3slivrlKXRxeAtb4iPYFL55o9FCVp+m
yELGHY6LYb5RaZ9F/4w3/noI4YiqqnOI/k+DA+EtqWPCheJ0u/f1qLClpS8dKdxu
B7FDSDQ+XZjHIAUk4NpDRmOWeBK7kZGaF4cuBQ3YO4vheQknkIm3GEF71tTh8BGL
HO7Wn8S0aaRrSI9OWEQNPvMV0qSPUh+E08HmCboychW6Yexw2ybEHwOE+vGhKTrA
x/xG9hcrEemTPrB9gJc8Q2ZVgkKtlwQQEcyOqk9lsxxUw+y/PSMutGg1ONgOpQlP
rO0fEyV+IY6nnlgtak9fTTuzxr20LkdyIYFj76iJUD5Rm2F8TMBdLJXqFs4/hA+l
Y1xb5wOM5VtmkLWQz56TzaVfxGSKguKj2WjBJZoDnG+lKQ5FE+cvJPGZqreqPvzx
Bok+bxq50f7rjzru89ZKTZepqBDEpRqzpV3Txf25me3jt+MAJd4S5LWAF4O0EYE8
R9AUlRF4mwpuvKf2Kcdd26HLTgiqz00iUA8axH/wiD9L+6u9u0tuIK0D11zIAAa0
Jb8V29NM2CAV1QFzcM1p9dnEb/Jb8XHkG7e03Z1LNpis9M8eIrpbRcvs5LoD5C7V
HPfKYwsaz0L30T2EhJTfX1Zl9sS0YfgK9XsHYUFdrwutg3V0GS20paNt9ygVFi3q
G8lhyXczVzhuzszqGTDfIZN8jtDNhig5vwSx7WBcOJjtXgEBzN/uJ3at9wPtxHU+
Kfg6VopbgmBb2X/SWDrGRTk9Gu0WsJLBIeql4Qweatt1ntApvohP2pvihiNPoaVU
65ywSnNSEkLeLbVDvju8JAo/ZAAEUUBCVHs9Wm7aCN85dGfV3Q64Tzd5GxC9eUk0
LNK9/H+TkSGSGIIiUbqnJ18ByIdEM/7QZUuHEn1lLGwo32HsBIKsrDapY8WOWFSh
cDdBM7jbSACjsXp7jaBuxuaPc2CtWmzvo/UYok+jRgWvzGD1MEsI/QCJZKOMZNNY
kKMetCGqVGP8VgZg+pMwXtUgnISxDcsvy1t4TAF9AXnz1WTB0Ao/SYYZBjMTYP0c
SMFsQTfWuCYbQ0X15aWY7maiP3lZj8iXZH11RcWNj34xmN0uonks4dMoo2EPgf6E
Im4xUKzCb+q5Q7E/rUwJctypRAdT1ErzsuyY8iXGobT5DpVrXLx4Fp6Enr9fncaR
L1wh1qHbIXC5BH+G2bzdn4P6+D/Hd/Phh9YmfznyGyqtKPh0eghgH1E9cKN1PSPf
yBAGMz0SZM2AWzltZB5bQt0fcNkwcZHmDi4dXoty0GyfcI50pI+1g8QJfwl9PxyA
iJIDzvrkQZkNLaWnQXzItkLfcBNPSyi9ua6bjd9XYi0MmGIAaTKJ9dVaEknoMUOg
GVNxxmItL7IK8vYhGzdq9dTaZFGS1TERivZYNMejblehaPlAj4seiSoHNNev3+aO
EAhDHZULVcBSvqmBgWwwUfcR/dycIex0BKE9gisXr7iUEg1aHdB2kjuHwPQGIYkY
vx/FMbUcw3V/nVo7TXxV/wxCKTlBcipkRGQtqx5VZainI/5pVTTf7Ie+QI5pz0+q
8Ny3b/2qVkWDg91BQtzdiiL6eA3pqvtoFCXWevwkioS96zPS5pqrakdhuX52fWOc
kH40sJabyn7HhrGK9kdsXzfe9EuavtsFjLB7VCUPgXKVF4Ww81UIe9NthiErTM0Q
fYXi/4zeUU68GsqUYlp7loeeG4Ds0IYSOmEGDV7+M1tI+BZUpW9WZg3BgnkFO8OG
9cM/J2hBM7ubF+ce1H1DeTUwOZhkt9ontfjcwRjmLinWbV9KZGckYI+47fMvKgi1
3k6jyk6RAHqpBIk7BLpGMjcqv0cbUjSEiSexfnpy72gsAYtcJfR0xdbVBxzRST0z
Tvz90dyPRqXxDnCN5YWfFzAGF4olVgfKwhK/pHiDIw4=
`protect end_protected