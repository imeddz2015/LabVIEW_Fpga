`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 4272 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/9huKRhRMtvnNqb3Z+UU7TahEoHV+T8U3P3ufru7l1O
3DlgtZzb9QxCbOjthp9+wDkjygH0eUfDrEl1ovhZG62SsWZDA8M+IK29KW82H0rI
IcCLHukLPdnk8vzIWDugz8Uf9ISCCMaeGtK6HM8zgaaocnSs3jvwhhEe+F8uhJB+
5rgnPZ/uyJDGb0TehsOsTrBWx6L3xq0PS/V9/qNJYMVg1/StCCuQPtSC+R0oEyyf
3rHxvS9YJkmDY3x3LdgYVbM4jKwQzJcWVoohefP3CUwWV2quOsHjWyLIVJCO2Fxj
Ck1wxMoJkpa20rZb5XMQPGevQVdPqGCOBwwaWYffmj7GnoBtp6NIQa5QmalDGUlh
9IwzzU3MVtWBydHAzvmOSOZlqzN6B8Nq8UXaWEKoZbC7FZmJKf4FZZLPC49kw9ai
kzH8YtWglGglKAOg43Mk8CndYv6TjbDuQQ3tRFfahFmcCreCLLeRaP7GVnjxSl4z
qI1ugMlDXmuVguznQpwVDtWQOJReazfb5I9tNz9Rq3jCLuU0+RmHwfrZn23Z4r3U
kmRQ37uZmCNj46gtpZMcMJhEeD8ueW0N0jslr1pUpQpLcV5XMw4E1oINqcfhgivD
H3g7duB8KWGZqUL/gv94k4SyGgAChtMPtKGJvrE2I5/EF38HWI86F8hX4xJK4iSE
hq3mijhoyGhJZ8dhV0qYvkz2GsltsgHcqe2kkCfUyJoQx8vJWrM2NEgGhQQa7YrW
9JEPdfh0GMC+YSytw4613AcG+mbbEp4su3UHlqPWLLzJTEj455yQpGhPgBFag0Y9
LkvOlL79rlo8jPATgqjNwDUYzMOIckWm3Ksc5GlQhDA9GRZm3UBAKaRmWZ7cujrx
e4+1TL3+4JF1PFNQ+7WDEl51EMiiOtPvf636SDKlRwBoH4+wZj+BJviriiCoRUUk
bHClJtgqERejmfEugj666FxZEMXwlOTmmP1gJbMl2hHEpS97B7f6Q9r6ZwSHdbRb
hP+iJXuJVjz5Fyk/fRIawS48O/yiadi5zp4UrXvGK6emNyK9mQwUCdljLEUUaX2x
RyGDF9+rAwnchm9AaI4ErpjmWS3I0MbC1P2IrIhwi7qq9c6SitatY1ZnDPDykqp6
DyRvS34Ihi8HYhCO4HVoRck/3uxfJ9GwOOoQ73UOKz1OMx9ov/aGAXzUugzlEerK
DItHJwnHvR1K+CIFZPwF+DqIbSM9mlRWm/Lhow7q0B6S0ynUQjZkIx7fc9urZXaK
86/5+2B1hbFcGFdSIPgxbjxzNuiMyY8+OYJdwQsXWBV0UaG2zANgDpUdUBE01lYH
iwwOrNIgHFEkuqeQ2XGdPQVoh/zeo3nrPQFyqQ9HrxGZKTcCRPoG08DUgJ1pl+Cw
tk77rPd+xU9L2HGZi/epsXLGS+a5PerppGlbW8djZkVr2MIysf63XB3ZYDHF3ty2
X8vHDs9HtrAAfVga0ioafnTZDLEournGJzKrodiP6Gp8eRs2TELDZ+yziMQJuMpG
vrd5MSFrlF0GlOoJEv71I+/980JhCE1DxS02lFlq5AgRcVqQIPnyqqjvK85a1f27
IqfaIFYBvoBLSKwJvLhg49Pqg4OroamG750AziSNk+BsBJscl7cMt9gktUT/itg5
pUyNCxSmRogD4ol48ZWzuxh5MUOGXKmtC7QVPL/FRVOMyu2qBaY5yXBNiJ4jSXuY
/778lkqofDOfsWHFHVsP6231nQ3bNVFCcONSJwqzkYezDzd6oxbzJgzZq/MEXoy+
GpO+jt8rzf5HhoKYXkRcHqUBU34/wmtj2I4sSVHtXeZZCkUAJvBRJwGIxIm/ZwN+
BPlwDf1RuA0mDlCfgiRfEcr+eNkDILiq63nzhzvcWsbu4DYHr0S679TH1uTfUxrD
l5ajk2xpm+kl1rsNyyXNI46os6pI+TWvnvkT5kazhM17wbCyHzYW7WcSD96w2uOd
usYUk3X2dM2iRMmE90F9C+7U9YH5yBz30+ABVDhCHWvb2r3FZXdubeC1lUZ7JbDH
+Pg2RDTF0snfJaIKWv4c8NarDbwc32eX/T4EvDF+qJB3iluiEe45AOkgRBSmZFZX
KwAgKO99FiHDBlKmTPOPvZ/MONZ3UawRlD38WbUsrLPH71+PmerO06P9/PjGzLdu
TkSwe3dQaFp7VwTTh0dfarpw9Y5pRk6uldNFtRs2dUDAH7JjobPI4zGZjxBmy+ZQ
EoX2aydWe52cRkMZX0At5hLY1BIih8RNq+oD5aaSl+YjrWVVrl9dm99bNPrxneRE
aVs9LWtVmweEwk6M/WhSEsil+5YQSoW0WV2L+prM9PCfLgjon9pQj1kAVvlT/PQ5
T8Z/IEiHP7l7CsMsxjPIy8H7TUE0yp9NeAzb25T/ls/9SZKUmZOa2jgNeYb93hJS
NRFNKliYQFbU2ti4MwMXJlV8oXD+uJnYAM4tw2nvndPBcwJ/YJdg/qicqjSkqCeV
E3KF0dy7rkCoFf0afpU0LbA0qlgC+U3Yeisqtz2UYVr/2gVtzsDgTHyAv7ZYpZ6h
HOGD3aWnRw5Nj95FjLa00Vscu03I0VmmK6QuwJ2yjOhFyg5Xg91PVmjIYz8pscC0
b1SIP44PLc0G3lGmnMSaSRUA+OLfpj8GG54Yowj6qM0W9OpFwS6URRlRUBdQS7nA
wXNdRTMKYbOj/ce87SMRJXaifdS7otIK2jmRFrb/z+gPXpXUmYNWhIsW1lI/FxtF
2APOyo1i1OUQSl6OwOve63VfldMQXSGJG51O8kbkCpdbkcJ7n0jGkj6YLPLPK13B
I6mrPheUBZgP2SsesLEvZ89IeAWjlOdRpprijo7BYmy8eeXPaeXvgT0S+RhVbuFJ
XzEHaGjArpD2IAezKGjkvalRKJCw0gx4p9x226FrfpAQEGopWhfbBluX3VK0mD8u
F+BUYN0b3LFyyFoZOHjn3bAXfHWjc24sQx4Lh1Vn/sSIAilXK/jb7juF20Hb5sqo
4Wg+h4pQ38v02NbDYeJ4oa80go9LhQEzN0eTrZquN40tpf3f1ek4WDuNto2GRoa1
cI5THSp8hwNHk4ejKlFvsiBxoce57Zgx360suntNSVrbJi4sh5P4dXuFIStrX/0a
R4MM3ylIZ34QGFVy9obiiBcTV3mE7fkiaag68VGf7f1SogWBP91KC2cC+zZd5m5a
NBZNhRsYoeqecgW//aerX2C+5fxkvvD6R7UTgjp3VofTFlUzyL3W+aGQXTZk+Vmn
vIsLRF9mQ63xVU1wQ2AtEQF1A2qu8MLoBxueJ8uQxcW5wo32Yf+c7jiVCqTPXVUa
0FGX5aNHjfvQNSXbTqWU+TQW7J3jxlbS2aO8sIyUnos8OKW+GVsuDBvDgudXQeDc
MM68IZi2eE8Jx0x5vRLRgrmQh6UrdUMf6FV52+b3jaCZMvIfuBQIn0ZfWM01W6Vh
c4UkrAtF2lco21WW2jfnqxpB4nX2wmbI1TxFvJ95U92g1xgWtUiSAS+wsQTiNab7
9xsCRqZ66d8tkodXeryqglY/lCJNMWo86NSW+03LsIV5wpZh0GR2jdSvm+8E19IZ
aK7zSKZGHpyeu1d/f93k8AVooh2oWCcoX0PTAjLISsKQ80dFy8iSttxwD9YYkgxX
s2BUcQesFmFnC1AjFsXI1mdWt8mV51FNJIp1cFbewUlLxEPTelejZ+MIyedWU2zo
bf8FkBBmRGv+K7qcM6hzb33Fis1gCNZ/qLHXwM9vv4t7U93fDxxgFDX/5spD9u3y
NRoEEoEx06Bw1ikPrIlxjiparCN5Y3oxXzTVsrGC18LoKoBAD1HL9/6J2RT8hCS4
ofYKD013UVERiljh8huk1bKb5tmxqPv+O7N14r5dkgMHhJEp0ndDNW1vHOQ+Ct+m
m9dnmBhOZhy9Zem1iBF14M3x2Jq8CpFOueLWE+QgJ6CC8XzI7kzegEIvETNGVKod
s+0DRtUBTwmy8elAx34bSrRVVjJx/yBOtfOYQVR6rURVfGSLQKaYFRlQHppe4PWq
cR6U9v6Go4Q4BbuCVYZBB+78ks11vQKBJhIGyEzx0Z5eaqJxSAiI9k3ipXBUbDde
qkfA+249sAwLkct8+DpyzVRTCJehB1U1JR2yyr7ABWabew9ZHC3NvLVh66TNUqQl
tCqpokLaQ0ApMKbDWfaU2Cza6qcVH6fhQytDbI6hN0r880Hiq+zU403TYe1ltP9t
e2KcbdOp7U93DX3Gkec+d86fr1imTupXj8JAkBF5l/MF0Dve74R2Oo1ILQKZzo+Q
qDkWRn/+jaG5LhR61eZkGCSXOjzIwK7DsfFjTvtsn5xtdZWndwKGjjCByxsCPRXt
WQrcjbWURmPUZ6L/hZ+TFI4BX/A46dwKQKwrzem6ghdZHWFH4jLYoLI//fyN2zhi
f0ptJTYNOJxY9jdfIKEoAAyZcSn+wCTejsmyfTHafpUFnvapJ7CZn+7eVV6jULGl
zAsYCHyorcjWitjy6JF1D81kHkEtDqyuAY7BfJRNRgXkfVGxcqGqGdzorqsMzVa1
NHQGTX3Rz8ptAouvxdfzax8Yr9lbXpzRnPdyh5CYiNWHLrTyI7vS9F3iHDcR/el1
KZ1xAfbX0LfUHRgFQ2s1OfzMyM89gQauBTOOxMLQP3d31NRCakKE2wu1CH84UkD1
mbTphkg5vMfYxHy+QJJ6w7j+6+dI7963jGJn5h8ee6cxR/jli0C8LE+/7zL9nPX7
DFHkPxhaFtQCOIblru3uY5WcHBX3r3VP0LatHccc0eo5sm+zzY7DrdouYCZjuaOF
par/M7r+kgJFD/jFmnkpMvZcwCyAxBRwFMx8lDWmJa6p04d4AAYsEAysxmSCnqdp
9nEO6lY9cJtAIe98JFUExE+rULuf8NHKiOYFLdlnvG/4E+sgjb9YLHYwO92vh4Nz
sFCfYYv1v3gVdZOuUntBxflGuhcv+/nME3W/sFWOB0iu7JpPHViMf8HSMfXE53Hh
FmoBkL/rpcjTz84pAO/JMyS+BGfkqaCc9VQGS+ehTo6flNRc/zwfAuWMyu+w5F9j
4KPDgRFdzT7bDFQJKXU0gU52IhCSGYRslh6qtO6BBbnOy4VW8dzidq181l/AA0gP
fwu+03Fhs5I0A0w2rVeyYsx5FAg1801SK7AOgoeRQqmN+jV0BnKiOYqjlK0UNJUv
X1TPzNmElWQ+uTLCI50ogMOIA7HRB/m7R0sjToMKr9+5CIwVVHVUR3rL/tMDbvzQ
DCEgyvgoIxrH8+G640Giuu0vnxFFv/nV5ivynhX1fJzlHijcKrZYjCQ5y+VGBwtc
jl2XTQZR3EO1WebKzx87QRM7RRehT6bXH8jEDlvDI5/jl1iLQJwGpXvLvF1Na+BZ
KzSuiGt+opO6fBYQRfOvnrp5DHmL+1yK7cFPJzgYMoDfQDHybgLYd/O0u5UWbA4F
pcKJOhQ3d9T9NBsusSoO7P7Iyl/kkiQt+guritcfq/1xL8dPELGk726JjlHwpmGa
DvnZrbxHTEglnum3uXc6a9CAuDv5ZaUZ+yJ5cDRIjTaMLy8yHpRve2okg6CmkTB8
ixM8HiZh+lzJoGvROYr5m5zXJ65q9wbYQvdy3Cpbcw7QonSgwS9U5edgbY+a6E0h
7WIYLmNf9HiyoSQe4hqqGpDYKIu/YD1E2DYQB8Rd3PkzWpHHP2EdUSrz9SbquIzt
`protect end_protected