`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 5168 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/9huKRhRMtvnNqb3Z+UU7TahEoHV+T8U3P3ufru7l1O
3DlgtZzb9QxCbOjthp9+wDkjygH0eUfDrEl1ovhZG619/hkYA0Kh6GbX6Zigv58I
F83K1o9tiRDBzjgxePD+9cjI2y18+fm1lHKWVW7RvDgfhQxPMMPXkp+aDVK/GebX
Ecg0O3BNCdqDHO85ztBSgpO3pKtlynOYwjoKwPrXoQjVsE3QvD+GHOQ0nANDEP52
TJ/5YSHieJcSezP9tVmcY6Gryjc4MW3Y3KwE4/ip84/1NEw+twouqShG0FxjF5Oi
3nAYy6PfAmZH0zpbj/8puLtnrp2crOvF1D0DdGmo8WA9xc7kZRF2zG4d66YFCAy4
zlw16x5vx2mwrni/yH/thHna9ihaVTnUh80uQxvkpqt5fhnQkrXzdLIRB0C1swZM
i9Jlj2bUlM9wkD4UBW+yBxYhR6GrB53vX3yEsnw9mg8T1UAEs2nqJu77X2LvY9OG
Kp0Re92Q12Mts1XTqAN3iC6FOUXULZ/0hcPmYYRbiljl3ztMwoQTO/El1muuw7dI
Nf4qUfBXRft4SIBBFJ5T2mWazsZgI9Rd4FVdMIJpKwb2/Pn32oatwmYQ28geCQ1e
AMS1tkIj/4CXgIKB/4097LcavytHJp9N9sOT5rNDtBwEoUpgoThhMpFqtjXUy5ZW
CI5Nmw8SpXEUN9TdQPT8CWSkyoLSv8sbY1gyTXkcK26/YSc9eAEBoUQ3+4a5vFmF
7fhlGuPR9/NQTEhShLvq/AZvzaJMUAGxu8domFZfTDwXopA8qld22q13JP11cG+6
xeJks+obxUJ5vj7yEKEBmOaF3YtSSpiS24cj6gF2Hp9lliI2UURyEN8YJSa1WQF8
k0eXT45RIiTWC2A1ZN9Eu3+H5ouo1Yw1uzfbVuCsITRBh+NHgEqKMPNOONjw8sZA
FVzvQDZPcSggb43LrMneeJdF3xliZYiOZJsGyD7FjcJYgW4Z5MYvmd5NuctG7qPB
mVU9CdDmAMrai7sLJHMkl6D2kd+UjYhEU12jzoQsbvlnNDEQf3aRSjkvBwArQuSH
mECz1klEaRBGBJfyBQm7P3I6MrfTRG1e+Gk1JErXWpISlvTRgGcN3Btee0cNf4EI
JzVcze4YLDcUZ7DIKxFr9p+9BCqWVQP2zVlOV3RhtkPkal9JRciwhOPeFqUekRyD
4Gca2zEp6g9G2THqRfYHFSiYsH7OlT7O2mbK5ZK4LkgpeXUR2l+n3LtmiJV7Uk8t
zFB2m6funE8QGYeHklKuKpy0TX8kFISywTwSviwqD6S54NeQ6pkjRe3ZUidmaOzH
IeAaNnsWd6s3IRX9x4oXTA6ngdj8flaAfm0mz1Fl4A8xFfMLgpfcMsWf46chs7MN
0u9LGPomRifBxwvdrmspxmyANQDgCd+pfczs7Cf3aCDMK6y48iVGIPWfZHstIVx1
msCDSCLm4dnDQYxqRts7dHVq15HXh3z/BTJOKdi63+/oZaHkTVWEGqWFgpW6XBjj
xd9+geP7GFysUSJzaxrXYqA45BLL9JNy0C0uX5p0HKJwTxntMx+yYBIpO/2BuMWx
01dwYR0Vfig37hJT6fjllTDpY8LUdW1F122P1cSu28V2RTrtSPS+ipn5pgNgtOMC
NAX016e5FKEqfSCDFfhBuMcX+mzQLeucezzS40laQB8vkA3ak5htALaEloFspUEq
igaSRHLnUNp8wsJIeGoxp277LGAtRCggSyzu8ddtrBHSTSOKvzYvsenFsEDpnmO4
z6sN9m1pnzGlflXM0eM0Llwcrr8KzELoI3CtUcrNbk2JjU4397ftDkQ4oqyxwDwL
28J37kwzLrThQkLgpUxMncZypV0co3rHzFehR91LsCfif2T3d7eMbshdk0LBo8BJ
q5ne4I9ZrvCuvl1tlWacjFEONZNJWvqZ0lt+T0Tolu2RxmAXlrjlfWH8tOJejmxH
jkwTIAgKHEqsAgUvwJSVJo0M+ZUEMxXzb4YH3HgBZ0NJUT7ecYtfuu11CW/o96bM
pyBYdHU48puHpwIofzjc96vdOL7lgoaYD77/rox/ja3IRqAw8MRhf31iaIqxL4jW
1fq7vmtlLP3Gt6suJ3bqJq945sD3OrCtglMh7/zOx+rniRXPxOv7PiS0+mRRpUhg
gzvayYo9vD4HO9eAgVcTFoULk/pScMoKCzWeU8VJHNTEIw8lzcxOHIT/+7rkwvD/
K/9yubTSxBshQXzz2o8zfJ9zG6pnTgyU2eq328JKw+dLOT1QPhGHXC4taPiJCO64
4FeXgOSX/eyA+grRNFHrPZ7Xx5/XxfQa7zclioOOmUp08caJm268onVTUUqXOAs1
N2x1a3JUEqzJZdhKu5axtosbowMLOq77Pno+/YLeeCKeTuq3U3UmUhkFSm9IgiWN
KmiuV49v7fdHk82ysHYM6w5R3u3iIncqwTvn1G+SBFv2Ud4fyV+efNR+zrkBYK+j
hGeLeQuAwNiPgDUIFQEJYA7GXW+EnHxGpp37ndQis06d1+6N7c4CgknlLbumokVy
xpbDRWg0pvN9dK/AY27ZqwesblqiVyCGs95b8DFOYXVxd/qiAybK/ZpqRfpp/Xsu
Hs4LNpSEL/TON1llqnisGJK6a/L0EIEcil2EZiydjvII9/44+qproE9EnuTSCTpz
/KIwS5dmiAFmOeAxyaz+gAwlwDKMWvMgrLXrEdeCmPW5kcPnK9Y/VxAnjn6u/j+w
yRsyZKRchq6Y0DM+cY+qRoex2HpwReLtzU0q8jrUmgUSbszF2OfT9rGtrBdv8Q8h
aoT4LCJqeExcx3NP0J7efVohe3mK9V1kvkLSTch8PAKpxtebXyan+277yP4qhYwU
tutD6GPdoPQAwLoVzbkf9slysMc1GE4GQuZYS2QWAojYli5T815xEidGh8hwGltg
QQVvl3bJHUuPZ5SmDxEfr9EKruKuYmXIkAmbcT+zKcBpTG3ecnzn5TXnT9CMmZZk
EtTpXh6Q+0no0r/p51Z9EkJ5hnGFI2SNplayTY46DRf9sZBOVgH01p9NKhKmbe0M
tJ4iboHm7U4yyxE1DLiA90bmLMuqnvmMVss9Mtrdu5G6gEztQOPHhcwhne9w7fmJ
+z/td85s2skdtUVI03hwK7WL9YLKrHnNux1wlwsyO1wpcWtENCrdO91v8QEzwnqA
yL9Js9s9WRklSOM8BPbeDr7sxiq4uKLll/MV465NkvS6nCBG/VrlumNxJiwcn/Eo
rDgU/xbXrE0NsXiaz/yyO5OpTcdXLXUVMxBVoXkMr3FumuqCJkiW96H5S7zyM8om
QowQW0YUa5ihu1uVYPTHhOU3WlGe29AMliW2FIiFwr++01GEBM97Gz5Dixx8M2bF
UDjuyZw2CcdriMJGeMoVQFhSOvEzuW6PBGDvYI/MnsASG+ooHFoVr2JWlOPnYN1I
WFy/WWldV7/KsNtiQfg9nXdsUf5QJ+eijTiSiitr+pa78FGZSQxLo5gWv2xS6Qac
/OMhdtP9zX76Eg9pq8+9OwoeZLF6VLean/wPbMvERDkL07CW9CPv1Mh7UXz+GUqm
NRte6B2k3pPFHBmFeS27g1ln2Le6qemSsNskd5zqalUUphQX2TdCZAlQYvqH8Jck
+sEx/x/SywflMOWxnmjDLh/jCFA3NLWwJTbYWHUbNELdWqUzKgi1p4Rs7A6lMBV4
bsP4Q5Ka07cJ6IB3j1cKpogrX55ZdTvYBW1yKnYzoTUPoN2Av9ingNI7fZfWC+Mw
Pqjv1LtTn35M6oE/K+bh2mP4XlF7qFAW/CbX5MjwmHtOK7+9oo7pM5/111cNhSev
qRsIS34PTE2nI4X4A0LAX7BdzEwU+aTv7n5LdsTSWPznRMIzPg/wRBs7ORoPKjX7
I+gysRkBmr/BTp4hfbCbgo3F0gxIcugKj7DMxuSXi95WPEUt6lsqgiBPDLouYJrO
vDUDLKkNYFHOTj2+wTuHcAk2fslzMx3I/w5XhQpqblEN2oCyqjVynTwFnrC8NtpZ
OmYz4P+iIHP50FoEa7jbeDssIq7yzletZmRrT87CMvtawQYIm6sW/8L34vJmoHYk
UbcoRvl0AfWwk3R4x/AUGo8k61FG8gk9rgJN0R0wm621GfyqVNgZiBRkGY9csxWc
vryMwKRLsQVyZ4lDfrkl76gvRCpROLxtqpbRKco01l6v/R4T5Njoc1yIOz/P0mnU
t196Zm2/b5WHdRj2fPjlvicF7h8h0eCdElmQjBhQDlZroxm43GD2VF90ojSOMya3
rLzNXmp7gHSQ3FiVSBbbX56BpxQLeiTjwNyn5yYO2D0N7kX5mKHSiDlS5we8MX4d
uL1IyWkE4riZ1xKmJPEIB8aJVjzDKP0ftQF6fdPTmwQTppTDb460RBY5dkxvoUr0
j98CucJJQRpULWdDP2/WHbfCuwk9vcTPKSHq4ZkUDpf38Lbw0luusosoUJc9IJt2
sFrT1gWSszVLT+NgDlqUPRHXKuQVxlhtD+svKYtqHqRfQP2aGGQMQ7PBQyAM9yHt
jQdfvGwriMLdp/IovC0lDnKnQh0O3VuDveQ5UblhZ1Ds0mFEJrRmqRhnXCwYGgO3
3T79dxb7Yt8ECfne090cdO0wC3aYjBHiiZX8VV2K8TWFeCSPskWncyKF4Opy5h6w
gXiSzXUypU3Ij0rxv/r4J7orEq5afzSUJhsYlepSKvay56AwnSOEpaMp4tlDz01a
Tt4Z2jpgNK0+G4PysVgKOyytPRFRtsjFxR8dxFvuL1YwBa5/DlsIztcrkCWSRGyA
H/jwpW8OwlK4lwRzoCZNJrlquO3k8E/JCOEYs4gm3yLMwSH5dZ/xZVX13Hahe5iu
5aiP7jj6YRMGqclPV+p6kg5wq9BXbd0ja+cZLwDxbpGAgoF59qZlWmixFTJfNbth
nfcZT4E6/wHNCVsU8N9yzohSmEtFnrJRN8j0jxgCO2wGD6/AzLsQ6R7MQKuHKdaP
2eLp+XT7IXEsYnzDh5v4XKvQHnwFbTzecmITvUnXtFxEEfGsBMpOJsUxK+XY91A0
6zIfQ9EOn4LmaHsKXM9Eu6NE9w7XtC76MMshYBAP57H/XhjRo5+w6uIya3MeNX8I
3sXD8pvuQPpWv5vYe6IRf5FCJJ47+WSvAT0TlbiPfp+tGFBdXpZZI8bgCrdUSsWw
p4sgC32GP61ZzUJWQjpODvOYOrpX6zt6FtoSEi33O4sbsiOsrdduqARLTuyXFyBY
9jtj8/DH1RwfQbSmqpDOeEDgUIUK7Gv2ZUu86GubOPRg+tiKOhgXDltIotAi3uqU
OV9Rs46btTEFlXGQbjvvENLO7ENhc4nJ2eInH7Z+HIMENYxW3egP2dm25NB+lv4m
G7mbiSCLcAhynFdvQQPcbgykDI2WIZqi8E5rPpltysR83w0F6UjcMEo78Cyh827A
GMyHLKh8TtnXh95J4twVppI5Au2cU/ikYNPDw5ayDaZ8IiHl2wAcN8wLwpmXPyBD
HLukCyH7Gu1ZilXsmu5Eh/14t7Q9MHsb8PufH4PCb16MaFc4/qpKB00vSHjFRH0F
IUZ80LJmpC7cEEZApiFE679tFbjZm8E9Dmr7rvphXeDac1JTjr6IUGspDHN19Nde
rZT0ZS++3dMqiix3dxIFHAK69Ryls/o6RHo5eh7EFAhW3koGQo/GQYnqigBYuNJ9
FVGZ/OfWwS7uvyYpHSS2jtM24IvQX7J5qgbwBhOPHE8s9G3wd+y1Iuo5Qi8xm8Hj
AojqKtVcPBWB7ZTUeWIkdEsTCCDP4TRIWkXFvKSm/huiTqgtY+4DTNGaQUiMf7YB
O3gaXoRP0QNvz2CY58lwnY3eHJl0S7bHm7XHgeB0Fdbw7bq+TKOhh8j14k6sGZyv
WevnGBPk4/vbZAiW1sXxXIu2deggxDKdnL8XB1OiQHsfpf0AzKz1qoTHGFQGTP4g
LWtzt3jyB1YqOh1IQyxRWQ/n1+oR7NqcNVbEZbAWPByM+DeGVJkexL0xlyfN68tY
9Avyx/zuj/n79jyuz8KpHt0PMtRmM1Nf5Ehnhu/YZGqlsEQNiPvPrfrsz4RCfL4U
YbXCQbMX6jycjSdi2y8UAdgYavIMMbPq0VdSKb0oCbnFDRpYank5YDiOfVTAXtS6
1YlmlRy/Mt3ebIse623MUQhSxL5nVVmv6IZPBhQJ3pTgrm9F5AWvzbeDqAIrYba2
UZr7IXRsxPVSiQgV1R2cbUR09gAqTqrMdRGIwPiJmSgcCzXDCw2tSXs5IGL89uL+
9bvcScdn71A0gniMO0FXFeJusSbXb0cPWvo3vB+TmCyFeDtqNcYaMe4x24eDKQ+7
p+kY7LCzt+boV57lrd+ozVNmjfmyo15dY5F9DNpWIsvZwYr4H4GSFnOjwKv19UVn
bd9O7HxZATcODOld7v7Pm7Y8hdf6e5iuPytIbdElJSVGCtX3x0z2A799m2lgW9Hz
vXO4SMWMZXL/vHit5w2vwCL0LI67f14g85N9iev82/MACW6cNGmoAI0bNaUZybSR
DEYVPYkgHHdAUvE0re9PiQ70hAaeD//uHoPkCvlRh0sxj9X+UXh/b+SvBvIM2KFV
AMGEYlU0K4RsevFkrP4scXSHuqeqLrqr1pY0RGMpfILoNtPH0qx3G4+v/XznXEPG
WWAI5q2FCTV/KnU6gEWWafTOkY+VR/+ffZIlVE34Qgto3r5ypg0m8Hn/z6HOi23U
RjljE/8vE7Ug7A/wYwYjMgB4y9ydKpErc7IpmWtdY2iZLxXttMhULkt1igVQtf7S
23YiwBIquJnbqjQVnPOn1GsSzaMW3GN+SL3ivRuKMo5mOcBeim3Amo6JThOe1Bp7
QUkD95FBem2HUlmB+mw8MpKpH9/cysfAgt29z2028rA=
`protect end_protected