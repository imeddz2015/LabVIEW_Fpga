`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 12576 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/9huKRhRMtvnNqb3Z+UU7TahEoHV+T8U3P3ufru7l1O
3DlgtZzb9QxCbOjthp9+wDkjygH0eUfDrEl1ovhZG6075wh2Iyq59Q9wxW6zM3qa
klGcngXNCFUmK+xvDRMroIz8hsfOWlxJn06OgZ4gqVDoVzOEgj5voha+eZZ0UPDj
lNQb2Fc+KIzWBk4/ooshvmuI4bgylUNFKkUHNhY8Y/OlXXlWBSxuUl71k0SX+oUw
7Y7y8PtWePkrZnClv2khKx1Od+gBQ9zybFIAdLTFMiq+qAkKkQQIOhK4cojjTsLd
gIiCSmvzdNLida931xOMK2/aTnzMY34fUxdXWzk+0dH05lievotAbxWi+H3XMTIQ
wAXD0OJd3U4fW/tLysG8CzQ9Lu9NOrSIPTD3tLi80fYIJbf/QcQ7g2ICo3+WaX/w
cJqShItQl0pYB1KIHwBdc0L1eZ4iZza9VzCVlTQJgYUKyQ9ralBKeK4vbabBB7Sf
Evj+NaIOU0nqgq0ZoTwabc4jvcRUY5Xz9k7VqbD1eUs4QnM6d7D2lmttA3uXyxfa
lTGRo8EI0WDnI2yN4g06EKZwtUdRPdE/Y3uXXzLSkG0whFAsq80zZ/BYbAjffU0Z
86KKUikNiY0yqqtbFzbS/1prKVUf5v78yj7Wh4v/Mj4XmQkDxu043ovMSDhifOUu
9FfjkA7DN+Fnl64dcknL4yw3GsyLjviMMlJ5QGpg/ZQhQxMdmlvJKfWp4c73Q5Bf
OpRJvv1iVpo5ZFDn0Pc5f++ySnKFxT8QeQdsSxDTg9Qq6FHtpb67PTcs+R9gt3nG
2KRpIHGafPG1BA8aqv32X72VLHZ3aVxwzuUscLqn7GciNa3u2mavDi6f4gXTJedw
LR0pSvQ26NbvWheqhRp59mu/gHKCEZYUIFlcrwjEws3x1PSLVNgCUANAFcQv6SPh
vk96+29/VTj6wCemI6yuPZqAfL+fpGpbSxRN0wjGQ7zGcL32v/yTxgX6LRXNSj/f
MSyHzNvxF3c0QJoamnHR4n7OC5vEVkyFHu7y4D4ThA4bRuaU10C7PJ/VHWE94+At
qCaVFLWc/CkAmqSptCKJ3mh9ms8FqEZREp7qeQLqDrg96+D9wEERi9DAPWbMwSKg
E4B6/sFKCfsXWUZ13BNR1bPrcthoWL5gp+cj0qafcyPXTgsjOs8a3CeH1P7AIoQu
7k3Ivn+WBzig07zQDb8Kq9F587BghQHkglaOl/oILQW1tHElPvS9XIxTyjTb60kr
I99qQmLReTxMH0YtJlv/hMxC4jJVH+8xCofqflKAKea7iIFE1Ow1MjwfZdubKW4a
AFCDOe5CeBsZwRx6nUNxFpWRIpLMhELom11jzjbsPI2FIYtDueMBdxs+e0toO96E
akFxOTp/RNQ8Dfbx3cp2/YUmNMVBk1EXv8a6P2soUkfMt3wxoz8PHuFP/TeY15Vm
DUsD9dCh4z0Bl9ecqQTn7jrpAcz9jDOkBXzUTW/GZBtBqIjm0I9TNlJnBPPtxqFU
SQtu5lIn6uEMYhCSiVNsRYklKCmTPwfHYmwW9rfOgFHVZISmAFDt7umSZvoOHMwD
SPQzZJ/We1NLRqVmGdRmZgf2uTYulIAXMRHFQEuhZTqM1iPXxWYHbuEEndgJva1A
unftCDR+1Wng9p8q2ODU9IcXYGxxuCGmhEDApicnmKDj1UXiYz1XCJknHPXsk9wC
8PdBRYUz5hlHwiZdbjDSDOzYZwvEYvhne+jx36GwTrutCEtKpVq9YRjPQSM7im4S
42e6NeJQ3lIj5xW9r9HEV+e77WreQsz7rFcaGMHkayH3AFdX5rDN7qvPr1dmGtKG
mbzbTIJLnVpWhMeMhl5R6Pa2cy6RMwE9ZosBsFXJJExGBqfwSivu9amblkN19Wu/
4FS3Snk4389soqOC/TbhBaU6wJ2SBatVbFFML7Z/sY/5+88U6Hmh9GPljendo5m4
L7MaKuY42z8RURwyZXAvW+1jJhpayKbEzVG15iKraXXsvD5nrWylOkGDhWL5zUxi
JOl/5yGXFB/2xMyl6+VRefTiQh5wPk2PAN/Hn/RQVmFRSfa7+QOHzIlt02v6+exn
RgZlNrThgHS2JvChLppjK4TRImORGKM87PotvnTO6q47Fl/E0mjeXBN20kq7UVno
wM04aZwhYPfXhPYVpyEHvH23zWgjJiI1ka6rWonH6uBWWBzFL9SOa0t3L6wIm+c1
33vFTJ0DSp9lC9xDvzVkyH1Cu5RjUObSaxtWTZjil8h/dqLa1tV6rHFV5J0dYkjG
QlcKZZ3ZLXzVDtteAppHeDz/ZWDhPUbFN4TJ9663K86TyNCcf6SQfj+fne9iE4+n
iH6WvSq75kKJoxMCz+vDraVHHYjDto27vuQKgpWgFVfyUeKBpBTfYofCCqriWHUd
nNncZUHF1ZUuhhWXUlsFwQ86DDAbgXkYJCAiM7Zj5hIaPZvdlDtjDP5DrEFBUw0K
XcqQfjQ+ihpdlFyQPqT5twmJ1yD9CewLF837955bS6btLw3NXbCjNR8ikja5lj34
u+cwFBKyFR77JMU4X/YkQWRN9liXDqxisO5yNwF2am+10u4K5Rfy8sbHa9j5t/wn
QpBR5pSFmMiWF0j0WD4YEyAXUeDZkmjvnP/6GlsER3A/F0sxe1KXefC7Pisz7CcB
zCC//ZuYGMf0aJe3WKwE4AWkUGBRBTPJ8MpSsvOgWj9GOHo+WR9YJ5S4DAL4DyPH
TX1sKg7cMwSUWs4YeEWGEK4pxxoSAG9itmlnQLgQQc660pPF5rKSxu/KoTh5kPil
V3/TMwJe9lQyNVyWCNnMe6Rudc29GfpOJKVBmeEb/cTYgtk/qThfT1ZPsp5mOWCh
SvGXAZmwtP9MBAW3jf7FO2pXfv7QcFC2fRzfVR6j/aTjMCAgFiG7d95hepucqz0C
fXx6f4tfufyW/ye1gX3soxovXzH3yNSRmGmiHR7SRYYkTmFokibIOmpbCe3vyF64
oEWCYtRVqMBPEab7x5BiKLidNumet8RzemFLmjiQ3c2kfbeiQzGJNIoy+2jBXnCO
AE7CKePHeUa7k//G0V1XIwq/0XLhUlTXRLLiVzyEAmE243zqwe7pGj0dseN/WmV0
PTwlX8reRtMKU4KdVqOmitj4fQ2j5zNCFyoP8khNgUDMRKKhp0qxpZZDK5cjmBtc
rDptWCKYm8+Vyo6dbB0RjBXoBLpmS0E0owvm/SH5fs8Uqtz2P6SYPcu/9qk0tkFh
T6dgPbe4eO9meEAchFaO3b2SdqN5ELm3bKufggQa6aqvQZX88MRvIk6dsdZwZk6p
mq7gK8amu3Hv3qX9K2HJDgWq90AIsEvv3PftCC/a9idLCu5X2ZfrS4kflryOGT+t
f+lhILTne8d1gEQyVCq9uVeQcRj8xZptAEeWnYhbms4ZN9MrpAC+DpimOxtzpDsz
nj8e47zQik4qgvG/xdywpsVM7/ur9nAtNg2iMP9XQNaDlH6gECO4EMAUg/ff4DT4
BNJQyB4+SEc2vN7gQ/NMdZOGXHmFgjFVO7RdKgU8SeE8ILavr2BO/Uybu4laQ9J6
4fIW8068DTWqh9n1pbk24SkuUqJFPd7azxJYB6kp92+8N4fA7qnXw+DUXBfn443k
4VS2mSXm+78VKXYMBCgpGv0OUi0zCRt6bULDqTRWeX7biOhfPl/nH8l/J2mGhZnw
TCACnvkvD2AZt5sG8nm4v/NQ8jD04BpbXCyQTGXN7ScBRgKSGtQhlvcDoot31rEU
wvtJIc0rmpjR96Z/Xt/NVmWOaaygXMKjmdQRs2mIstrXcyXLBDAvzgVptJY3h/ul
NBWrs1xkmixWJr393wwwz4SaMj/DbGvCX5eVX6gWd0f/nj7deVYbXiTEZMWwyGJW
YGLYHZYTmUurnCJAdbGoeW1htsTqV5CZW3yZ11xA3u8gi6ryWh7My+BLKNvPV+HH
Ype8rzgZDwBIV2jV6pn/D4l1MdwOddBvzxikpfO2umb4juiehHHecv0w34RgDy1a
Rhc8WxsnP5esxrXmjvdJ8THdQAll/GvYhb006NoflMFDCzAwdxEAz59ODq4zcarf
3iCAF9pYmprHKmCgzNH8m//zRyuSVDiVv8dXdKfYJ6dHnsEQEMoQvClWbGmraIUY
UEX4MsNcjzlECY+U+Y8FpYQ8GrTGAtPUPFMF1C1XGPBt31REZeTqd6qZnM3DXOKy
s7rYuQHZ+NRIW6wn/hRbAmu0ES9JHlIujY5tpSl/B0Anmh1mtUICfOEajf+3kpxt
Q2/6gaFh4T6mdngb+9GHRuNwjVLod/OO8QoVR8drd4mgM78SIn0LKMJyFx94skvB
lgo8eFZJWoPQjUSorAhG/OFmR7HHTgMrXleRc/9Ky8qIiNMWULlv13m4YCXBeWar
3XwYBYDodOBhZqaB5K8qMBQ4xNSF6h+XUw/qE0RnU1yD1d/Kt/WYazbCoonqTEC9
qTZGX5NqZltJTS9Bb7/tyPjkoqSJpo7ZYWuTBJt94gBB5uGp/wAI+qjWIDPzQIe7
cFjRig/GGd9L5zezyQxSGS01VnV8TaIe2cnd3yfb7h4Airkpa1fPSo6Ekfti8QL+
zXxv0OsQl1DqE2xoViiuNnwLpNOJbB+0BKoMCfnGULKxgMsHbS0MY3MsPRITkJEE
FklVW+qiH2aYU6hfvHuh6shjiAGDYz4yTrTJJva2ygbIoJbmuxqBXuGdfmatSJyf
4nxbNzTMA2dPC367r3ALKywHJGFsZ3c97LH9H4ogqnNqo4tJ8lWogwgGtapdvVO4
oxESdH6TD0dEKlDDloPtZ5HP/0htmR9WHidxq/rP7EgGTfpmkjZ2i6Y5K390g3Fj
l55cPN2MC+9UsQpnpsY3RRk0x58pDhSWKh2aTe4jpA81F0MRihjisUBGNBpjdSu/
d+rSV1ti212QT1AXU1c98AMVRmPqJ88VWaaGHZzaTgyGhBLfchmXbTGMdzJpHzPA
NGGKAmz2zP2Gr8tblt+xN4w2ezLBjfTmlzKkO4aJ5aQ/cxD18GhctjIQ7DadYvjm
MXLX8iwPkv7e+Km8qMoiOHtCjkOWm5SHkEgkHiIqkTNCZe+XFFhHI0ViLEtZm2xG
RHVkd/6WPhg2ZL8tj3/inBAfwuYwO9jZUxyIjsaQjRvg45C8gMDVCYpnGYj1SuoL
hIJIJdhy8gWMkIa/HLSmmtFBz4O63VWjDsNd/FBwuJYvCErv2N/1YujX3PDR+KSQ
im5CymFPo8CwZvm+8/a6Bk9E5JHfENUjnI1hHyQjx02lafxbIlgPiLWwy6p0JF1c
D0jwJQKk/Bsov/7I/szlLxgPUyRCSSY9iJJTzH40K6+AAb0AeLLFiYztWgAs2+nG
s2p3p7l2coLccs8L6+ZDR8V4Kcgg3LK24mxN4NYLllVghVCVTbQhhobGl9EFQCXo
LJvMw4d8fkx+952H4oaInkTRpSWnFGPPCOpZvrYgY+aGiwg0rUh8tr7Z2hWJo9PF
bdVHNZK2+Cjmq0FatcVmNu/giMy2l64oMYBlf1UUinqrPFYu5MfXPao/JqeRS2mO
IHPQmCoC/boxgDQ/p75hZXrkN1DofRBYegCu9MQ2L2tvgn48AGUhDSBKoacBS3cs
tCJslT+pT2+KpPtIsKvL9ixhL9gBpENwFE56weINkzgdIWzbTRABVFzy3MySLAiZ
xpOT3Drf0olD8sJ/rtNGPzlfZkxY8oO/AnXFezC2QSSd/gShOk/1uNaW38EFMR9M
Y0tAFb1oB7xoptHhPLTPsepnDx9mf+t8Cx93SLsE3CzI9ue3vbhPxdmEgGU9RtOP
jWt+dlur80ZFILAcxY7vPEmJqf7QgxEYJ4/m1WRxwAv6YHpaDq0tu1pMO8IKHII8
zk6Qs6KJagJ26NSfnt6gQj5gwv86upUb1eGxWdQPL3CcfIatNiD1PJ6SzZzXAVCI
GFW15Ympc4ffqxlwGv6ujUJyDjK7AyOdVzCh5mQ/zDTCij2I79xF3gZ2BEE91JfM
nkufzzGK7aoK31bZLHnyR3i+MgYL5Vdeb6q3a4VunhzlxAnTh13QA3y6OR51nfF3
UmUYyonrY6MqI5z47Us4Gjs4RcE2ODfsF/0pvRGdvYYAUMDFGiMwm1zmrfMmfEgZ
1z7OcV0kSt8gZ2E7/txQyifrcKiGL2SQqXDQIGrkylktnLD7dGb+R3mwFqllz4LJ
JEm4l66/YeZ5YhmllPYWng7gkExVdiIK8dYqYIP4bMdLx9njrC434JGqJ/sBwK/t
zW/J20LN5Apaziak7Tb/gByg0sURie+IgZeGE4vVEb1S0bZOOEQIbgfH8S7oCebM
+jH9SZ3s13UjvVXX3W/1aYU28QeWhJ7DBoYLPnmSaIaK3d8snEss9WqL3pTrR8oo
aTK3MEKBRPz5yOfEYKCZsejXYEPJZ/14V8UXJHT6/C13wHvbXI3tj2F4oTsT9EeG
8QZSKvcpJ6H7pgkgf52re1EStJhWFhC+QXdGWPmtExVBVCQkuS4y+S50z/ZL29Es
JAClSOZXT4QAKcAUdpsztu/RUmIrVJIWsvpfDYE849S7ys4nwZSG18xMmd0EXCRt
u3Z4HZiKsZHRfsnzfT3jJldmWIeLRuJH9UKcjvWm09A78LpXZrFgl6vn2kUi2akr
tbFueV65P9rqSwPGca7H9eQZwWz8tiPhzLhnFgvx+T9XPnphEjRqf7rHVHxc4oYv
BrtRTzaniLeOi7nxjOJNf3m/saUssLUuX6i31pavDYkUN3lR2XiSbAn98Nr/S0mb
4n3+pVAGeE7RsC0IK7Qg35+ALfEWodSHhRxzZdOb/sfh6Z9E3cSeO9AKCQNx5GwV
Xgfn6WM7jwUvny6ouDvFcDtIAd9FnJghj+XXcOqm7EaCILtJAwiUjFXdMNSRRzPU
KVHSOqtjCIIXv8ldWsjriI+kX/Plz+Q5o6cBc3jl6DBX3Mr4+5XPw5kiKDA+8Pvw
XdnLW9hjLalpMIEBlnJm4dZEPvZV/LZcs4SvPPsokauUFXo4iKaHqs7plAdYGb9h
O/tlElawjEpC+upCPhzcgBs/O0l/AIMbYY2x5yS9XUPU93YNwNCSBjkSyJzyDn0P
tn7JAYNVybJLnFftrSdZ7TTdDJcEyOX3zox8rOoU6e50auiUnuGBOjmdVp2KfEvs
aEwOOC4gKL80+zSL6a1b9d/q2FzU2gm71cIUl3bd46pl9esWnipAmjch9GVH0WxY
HSHt1bNsK55pP35Zd8Q7yAjYiZwEcpa3zhwh477H52Dgws8AGGKL/igUIxM4Y+Fa
5GYm81AgcBI3I6MClPHQrel3R9sq+5IoBwB3vG8gD8z6O2a8fxxxsv460z4M4l38
ksd08GqbeLEiKFYql27lFRpr7T/KdrnEfK8z6lLJE+ZOFrDPqPe74ha17W8/kOqm
h2elnTJ8GJwlQsZ8BILuI8rbl9Qu5RjQxMh7hNuOcIv6X21FyZPJr0FwpQj4W8M+
MCopx7ZL8GUbiFmMcqtSZA92NAwMVowkhAVEQR6LyEr4VJjzfAGsW6dz74A6wz27
V3XArdoraTxmMR5cPcIdySA0V0nSrrsy5DxbOJBvseZNBuE6xM3Rc9mR1nuSAPBL
Onz9y4C3e4eWJP8r8mplRMz1b+neBHHEkD1BKA5Yxcwu/EQ0l7SMOkrdhOt8WVGD
Lv2mhS+J1q0Rm8owMckHz77hCphaSJYfUzC4uyNqyMYgSWpvgo24Azpe1+npjw5z
e4NpE91o1R9n+OFu43yuu6nuoT7zLZQyXnJBN4/pAY78wwGe4ZMCki1muTLx2AUZ
9GP8ZE0PHvrmTcyIeoL7SWdEYARRnEyYQ0X1NOgN0yvy0fqnvDPod3hCq0Z9mNhQ
/JCIEX6O0hg2EZtUINWzqt07pj/r0+nMfht93mBhw5QL0wy5SQUO/jldcfDZKv3Q
sk1ks85zDsoDHisi3d+Nq9DyU2+NTqEnl0gaiGJQnlw8BhNoMpzH4WE9cZtSKIub
7OERRS4YcFVNfL51Zx3UcISZay+oyNbqfcW7glbWnRgIZnBosIi43vp/CZf4sbt3
6I/62yqgskvX2G3wxs/XnzonUNY4IFJu/mUB6QI6NT/NyXlDQjE9/LJNWKn8AxKg
HfIVL6Ugd2SE+LCCXZaRsCHcDPikKNXn771P4jKj6Xaf0vtwfBPg+ffrdg0OzaJ4
DPy9w5cU5fangmFdTDYkva11t5gXyYfNdnrayMQ2kgkzddvO2eqsMDyrhzw6vyNn
QB68qmLmTGSalCLXa55MK9Z6rqyI7XdsbmtAzR8KP1CpTviiV/PM91o9gFq0apPM
D6PLm+Q6qKyK91RGLEV4gLzvXamA0zemaYUp0GG2PQ/tLPs1PLv0j7jvpLc8cvst
L6kbYFGu206eKNYH17MmAPTD/LxBiwCdP9ajMqEf58963Odl4vQnkGtcIhcl9F+m
TDYR28FMu2/JZf3qDNXEhqrewzc+pipw4dwAWgp3dwAXbX2VX0yoLPKeTpzDzGq5
yxWj/6RZhoHKjKT6hsDwLJE3EbhOzh612V4rL6vMQpXyNP6jV/8Wnazh+JU5Xbs8
F+bJxH/SEXii9zYILaOYnd6DPkLyWs6WPZk7/svULzSM/OZp6Ng2z5HmqQZd9dBU
x3oLnDmeFLZlQbRHnN96caF4Y46RGg1590u8afv18AsYQa9u8JWBjxrviMlbz7dU
h3kIRWxbJ+layv2Z0z64RROyG99S/EFNT6UTWi5eD15secBT9FEDc00dw2bugIt7
t7Gu3x02UBpF+o+v89shPqROQ2aYyXtvWo8HNxshJCNUFF7pxaLJnGdWu1KYumD4
Z5JXpX51NT/p248/URDjVkuyzsFAaYTgntoAftC2sKRG/eeXB+DL/BA4eW4ohMDy
bZRcwQfvywGTXOysLTKEloOHncS9t8NohjOq07HNDqD6QLgkFPb4FSZxpMvVeyOR
bJ3r46u75teuI18zyHe1o+p/JaffHeLYJrKAp0qKPfCMJqMt8mpR9utlRPa3fIkc
0aJ4wy7wtGCZ6yAFgd93dxVXNt57R1yyQ6SjDroXxTzhNmhUpDp2DH0GaG5yNj8v
e4d6nMBNR2Jyxkbexmtv2HG5FVYCID5io0jEa5xTDDF19EHPuVZFBiwvN4616j9H
5hp5dg/qlgkMp7CAGt6islgoAvdhOBWk1QXsycuFVaT9P2qqoF+q/OGIbZJPzC0w
51ToawtBK+ZSbjw41qe+zKqTL/5gVzZOE1SixaF7pfwBR6DPlnysiXPdZ1Bv2J/q
nuL3Mtqz/Xpgc+SKsdpPS9PGL9Mo+3Ld3P2zL2SeuB55mYMm0lc3oZa0uprkKt+j
Unihx6pFYgApzQUSVpKWuJXfXhag6g1NCU23HnVW/02OHjQR0mL5eBc9r2s4izbm
wI2FhkF9lX6/Y0EBjBn7PjbwjdopbMtvSd8LF1MsP72SvGgBpYzj+njykSRsVGDX
CcrB1gyLTzLeyzYo5pBCSjf6JZ017pKpxSk9g/fXi5KjBMxNDMFkb7TswGaM7rXC
JFwiUhLN8hs01KFphDQMKNZi9SSGiLrA2fnvxZMlM4N00pNmrx4FFBtTJvbc/ex+
xaZcv8uDlkwmCmPKJll0ipvjb0AoHxgFkJAtMdzrsyv1d7t8pXBG7Azg0ckgr80v
gkQevHPDc3Cm6SAoi6NzugDNyspAETI4A/uEZXxO770soSQ/iOECot//IL0KLRfT
nOvqcaC0hvzLSWKCT0+U2jBqJ3TPLGQBO/50cbGKDln0U0pXjKh8k9ZwOWUY/cca
e8TJVKw/ThGJCoXTB/A5oSBA1Zs0vuN2D4O+TbaRi74Sn+LGVtbh4t9hAs5wfhfN
VWzDBBpO1vp+5J1QvXEVuvQu0Jp92Cbk06N1UV70hIK+3IkTCihZoqB/PF7ilCm5
az5Grshnch6fo6KUaoRLDAFll/776vXQyw2W7Xj6KWLn12ToIjQppnNT9NDZC+oM
ijfnfe0qZtwcFi6Uro2zyqsS1lQ0Sdy0iGkXYi53erEAnUY2pr/k8jEqz5S2wRZg
Jd4JcPfwOqJ/IgzHq96jwKOAw/qHUnVLUDzhUi8wgmH7JWPy+91dH8W1EUgwpA0Z
P5bsYLSlSB6jg2EjXlRIvAZmQ8Vtk3voeP99jfZteKTt5zGXDJA2Shtnfw0ffBUD
A1n+bvSfUPSKTOLRo7+uiFCqi1h84ocXD+z5ZU87iuVY6+pUU1kgGXv5NJ4R+/nl
bmjaL0L0wT2UuYnyreu1zbFKggghcxTh/2/yJvZBJpFbhEsIyeEPLPvu5LodGxX0
KG9DVxcZ1PMTsb7McoCwzEbYclFrkE6V4T7acfmrdesA3o9esDwhEPyEsuZI2Bbb
lcE/DlGBD7HGPr8jYPB5lbDeBrDHl19QXDyNA3pXbp8fmcV8ni+dblYH6aGi/Z9M
G1NCg3mWrf8YUGOFnZj9RO2fg1CdOcs7STnbH15qbKj6CTestbo4P8o1jqO4oJ7B
cANJvCz+DJvRes9WgjX7wrWUudVVxTwm03ltLpgJGpT6H878i0mODe+dq7dvYwZM
CjqFPYyYhMzWZpJvJNon/KmM7XjJj8/EWJgsbC3c9QFmiHJYBh2XS+EQzbXfMDff
3qEqpTvXypYjjhLlZZ1CgA8ntTq5GuCo9XPGX0cgQSV8rswCgNLuwl0jd8uMpdIn
x9jOwc19k4/qpxN5vHjXCSm//RjQFMGqg6EnraSiuniZf4CeZjDVvg0qANwtXKWP
tX7RD7m5v088I/VIfVAopLhH420ROSiq/XikeOQEHnPEQd93tU41evqQgM0VB6PN
QTLLGzIcxfI0ztOldW7rqBkiv3TqoABKi+MIakDx5MX0w/ybVieJDDPS9aobq986
pJA26v637UZ7qlVuB7NK97pYGPLPW04xyedl16D0X9oLn2mAVH2/mACktGWOAz9l
L0hlTiGGThKChe2PyyWidfWM0uTTph9pUKAo4v4EhU4oa21m+tQvQYBVznwhKj5l
6WkU/vOncdrraT8a0jsbTdiRAp9x2U0lLKsbTFzoFOPobVcvWyqKgIjmhLLmZ0Fa
eqNWB4fQBrAQJnNE0aPv4KnXB/MOfbfhBg2KtSIiKhXpVMe+O3pjzKdlv/rXasL1
EubwsXyBn1K9tO37UypQVfwi5bdlVwp57fslK3RuS/YYh4tLnl4BFvM7Dj4eOszE
uJRbsZQvNl9W+A/mNkv2UzAUZchhjz2vlxH9MUDu25QzliOkbEu9al72Za943w2l
qYJMC3YKJYT3/MvA0vA/vbomM02hZg4gNkziBMGCfuuQcaqGbmhPUYHAwNuj6QOE
cHHImM0vw23ib5wMqH4HCLf1s8/Y4EE0ulaBr9HcEihlFTGhr1hEsFOqMb/ARiZU
5bkNC+nwc4jrxNTxLkxaXm5OHQ4gBCDO1OS4l/y3C1iOzoDS1siFPLHXURpkI83J
WQIIUmoC2JkGGW2knoLJ6px/Srj1616ouSK3ydLqJJrbpxp2LXTbMtPnoMOxfgYY
3Y4t4tUGw3wDnkp9m6Qy1C5hMl6M42PCxAvqXbwWjO2F1aT2pI1HHH7/VJDhEfU1
9Z02ApQditN5c16576eji4Ca11cldR9Zy7aAwZXpoWIq7gNzkntsigHe5DL7BKY+
352AdiQ5nV/zGpWJGak1+5Q4ZWNzUFZvDcvSCIHkwRR+OczDVLAN+r1TL+sORDhe
xhXeM1yV0OEZg9osTZglEb5/dhIWkHY2f2X8wEc1MAa6ZUQSPLDpxg/OE1tJloAn
S+wrcW3ole1sGjhVovJnID31A9DbkJ0J1XSgYvqBgk/YxcwI3MyAe5NDsERnlPmP
IBMywKEufrFXFiR43AGNl1sxGDdiUmFLmYWbAiG9/dN0wrXlKkn979JD+8uhNk3i
EXilGvJet267pnyCVnJeL029r+co9nDI3dMke5uCQDSNfM+ZxzJ3Nkd3Sk/jVHA/
4sXJhsMsB2HAnpp7WKId5TWX+q8gkxYNqBJ4yQASxdrpAv0y/REReSJVwfqytfg8
DnXKwq2Njg9sof7ZUZLvzg6eHvm6efTECColQKHTNe3/Fgn898UWwiZV4X3wMXe+
bdMI8RVn4meQqI0HDZuTVNntOc9mD0elOSz0UcSBofmsi/JO9S6ISfGjb8x8/Mlj
H+LEYIaTJgWDxJKCNEX3i4JMD14Peiabs73yk+waUEJVuUXUZ9/1D6Py/cfMCFJh
1ueLtEEpe09lsGOYcJa3vJROKoEf2psTmWc2E4cKqzjp6RP9Hi5v9rc6RV1H+QsI
i69fqMzIzxl9PIjN6btUofAdW9UpR/EgKLyR+xUK2jqa3hOACkn/ZKZxIawCqmFf
gkhf330M8ZEmemF9nJSDbPUvBGbf4JMYyu22EjPLAPNusxA7eCWnm2nhz6Ztua3V
oo7Prvcdqp06zY114Z781WojwU2Y8MGbpatOoxmB4ehPA7PnlYaHkE+FS6hiQ/RI
DmF4TmM3zxwyLdaedDJzJd9wv63TqykJHuyYya2pBeQcdv45I5xBXZzKTnho/YK4
zpvtQUOWkRm+b/5lGQrfi+WLC4iTgOAlODwv7KZJp9RxA1DF/h3m615FY7g56VG0
ekQOL3Hsy3y5hDreREQbqeyK2vqGuqMPqOAS9w3be2xKx0kauDbRD93Xdt49wWoK
0zblFkjbRRW/fYtPiqbOkTbP/IV/SEmaiLF2icqrYpJvrq4332QvW+uRumDpdGA0
zvG7THmHn1YYV9eG4QMVWsX1Pqdc6Jcrpj3fh/mgz9QmbUfiiMzn1WygtquUvyQO
fuxhSlLCGureGN6pPanLwXL8VIKjjUgoFKgPnWWqKWDjG5ZkI+3uzrzVEtodNOC+
wyJOVZJfs+tL4L8QuEn4Mu4MCbu/dmFd4gQu1Ud8B5uMgzPry/RBNXq6zccaCDqs
dobTLX87+ISrwd7gScm2urmmnmoltrr9vFVZXfxvyWecw3Y3elamswsNal2RfiBs
W5frU191k4QmOlWqDI886oUhbeOQrmWeMhx1EkHayq/Nn/HsdFxcuFTs2y6XQMJg
iigrVbLmj9Xifjw04D/UZYzy+5oyf0t0e9D/wwaebzMan4p64WX8B7SmnhT1bmM9
tLVS/tGqKUDE3P1CK7S/9iSx93w/lryjwBm9SsHSHtexonnle2EJAqeFdzCuuzFs
qFNyizeceXB0mlwpYV8HyaISlLO6FE7amCZ+cDYtMKMrSr4WfaUPSmoG1FAfms0I
T3uym77S/cH7nPSNmLFC8NJ5LSWHX5aDowy9eTJkMbos+3GO9WgriIgLCyjvGiBh
170ub4ZMco6MHFeaGzHeDco/hap5YOqgeZS33WEmHF48rBFg+cR2RkayeekDamD7
rtjYn0uvKR+vka6yO3KlvY58Lga9MwMeNj7V4kEy7CPCsjjizjbluvMau3XYDrhG
1u11pyw0woEbL/mYulT+b3P68OKAxnMyDmnUqm4ddU/FYD8QA3q4or3hCOpUSOhP
9drwS6vx5UnkJGssy452Zj0WpazW1mSG1oji0x9gcW/GvpJM6fVJEMR2MaBSSMlC
Np7TUkuUHYYidNlh98L7jx0sl8rnhE/2OVDbFpoQA+D9+rhnpPJZjagDsfpVV0Rr
LIp2yUr4ZZiJQa19spF8JrRy9lfkxQFuStvvQHfWiXIq/ozxZBVH/dj69TzGibLp
L9bMRMpoB1xaCZUB045Gs3nz9RmkEhvhIeFBZyAt7ykRk7IYBH3gVQ//IGKfx4l9
QNAY1rxN5GMdKlNJrrdSl5NbXnVkwJ5roqivBKaqcevo93pfIajkPuxafpHdtjbE
fCSbEHyhgLCM3uqQCeD3v1zMP+TOEjNF8K/EHcklRxwvBzhhUfGP0y7bswDJRfdq
41dWim1I9dBFMY4KvA6kH1pqEvlu0jr0FnkYFEQJjEEY/PWpij/CJr0Y2utpQLsk
MWt7EjOGZcdRr7F+NekMelnbO90GISP+WlGMbWMfAHM6rlhZuIog7U7VIQL1p4YK
Y9iuZWzYFSErDi3jzTq7f+JWSovN/dvB7xSI9TmoBc22H7KpsGBWR2KVGzBQV34o
Dd0g4Hf3hhdNrvK1DTP13INytEEiB6G7JkaZJzGX/RGLNUe82J79OtOf1n+6seHT
W9nKCc2EoQUZl3BItWyL85K3kSF7s84WRNtjHuPJmSw/izUslZVpZy298HRL+kBP
iRwW2BROFiogo6TBeeI3tJD5O/yUdm5wioAOBND+CjzzEl5L5jj8PTc6nyDaOCG8
J0mxWPBzJzgDCAEZ2XsTMho8h6SpGzOICqukOCiDYh1Msz9ana1kRu2gjYQWqwWc
blOFLMo+ukQHPYO+elcr9+J6GChFiC6b0pcJtiEcytjR1N34RvK67v4RFxi+yiKr
Gc70WdJqurz+F/dM5n2MXAXnytD5HIXOXq1Fr5F7N0pFO8zaKV+37MekvJE1rJzi
0NHs3SgjxHfEdbxmiDZh3sA8/xUjP+h4JowCFENFs20pvDvE1Zo2JNErDPrcz6gx
LGZcv3N6s9Z16dZlFfXAGDvvXRiCLvi0leP8gcGLk3vw3Og05IS96KL96OmLrlfu
re2TklhOHuxnJ9pp4tKJmexCehE1nxeuZ66bOdiWPpB1cC/WNrXw5N4jpavnldR+
8XoyrT58v3QDsGr6fMnlUFsZ4LGS40ss+KxUevNLRfBKUBl1YjIJJbb7V2vv1lte
3+HIGRCbZ2nLokqngcvDvDSx3QCn2AinbL5cti3g0/36Z1aOSckVK+NYHMRjv95V
SqHMRXXRpRevwGogdSX0xz0fcnPtatPEL3YABomsb6Jzq6DjtofdN1JxkiZY5UIL
Gk0O1xhuJ3J4Jmm1L5sOQaXp0iWnKMzYsF/j1M7PxInvXsL9yvyxTOwaLpyh/JUW
6xkJLhBkMrPkfdDlCqHg6fQNtzNjXIJvgu3NS82w2kh34+pPy1YSni7kfXHTgfh4
ZLHH0CShM8EDXC98VbPMcjXh4mrm5cTPCuzDosU6w7XlWSAoaxi2KO35TknwZSId
/+WtvyAff0Hty7fHUJJjBR90pZTr8jp0YWTEhECg3e0vW+lrAnGI6zLCx9Zzikuk
khTk+qWbdgn5NQMsz7f4Mx2qRTtsvwa2UWmUhip0Rq7DSnlTvg2r6LAZnC98agl8
ml3crtQzVVQngRzeZtqo1AxQ39xrFylTyB6HwRaerrrw0TjFIOA3daNHk8LM+7PJ
0lZM7+cGPwrBU3re0dryuSpnXor/kTEo61zZaP/VAkkCha97cJI1fFI/d7MF4j4G
MbbDRQBW4kNSfM7MiOk35Ph889Lgf6CxbTgQ+SXpsJ4Ae5lZ5F6xSvjgkCQvjK9M
a1HzcoGAaQ/rKHLPklWvLh8RKqQPqecgmb4II8/w+DjbainXFJi8fjtCA1hkFT4U
hvGuxqd478P1xBxJKCRrTxXAeK1ThEdz2cNOJ6DIsHLbqNRb6ltmssd7QmtFyv24
FQINm9PeywwnHfJzldilL8TvQTT4EAOnbkOz8GJhR82fEfr/YGxqeV9sEnZlXnt4
Ui2ohKTv11qE+9vxSSeZyn0J9L+qT4Ldb3J7YRo8FHLX/TfQDHkjmxYFWgrjL81F
UFZVwrv+N7MSjaviKhVqFT3MEt1ad7NsTaJ+mxW13vcLudQ5+J5oWygfRORGXkQk
MOqHPzKSRORbFW10QK5bmKI+LO7gI4AdqZtnU+CXZr/0pDMPzVjGxsydkoavV2LC
33+xr1Wg0mjm9312VxTVOog0IJhotPvqNGKUYFCK1iF66OP6FysjY8kwauzr7/B5
aufWxg2VASwVSB2j+frIgrlPDZ5X4zB866rHUaGKBKfXz1rDgKiyZXJ99YZeF07k
yI1o2pKIj6fTPK9N/6KbqZDnEqA9vMl7Yk0Z+ZZmPiM9lnVjLXHy0V7jLP7r0I2E
lOxno70Hr/IXJlAAliLABEqIdvBPwGxIwTtKCR5+hXgtlpg5CkFEIO3e+3Mz61uP
P2mbttz46rrfXYj+Bu3sk+5UHX95W8qiN3m6KsNfMu6jHKQErOLMCpL750ARhhWJ
wCcr9QY2xZzrKK/MhrbNOHrBT7EsuFx4Jb28TKi7i9h/Azh8dNcaFmmAGENZcgiF
o9M1M8k7S45YjaQmOJzl3Zn3AUEkMUECDSv4hZJ/WuIyjZ6Kq0VgA4ZyDhm6Ec+/
X8JKp2lb5+19OfT3FTdM96WfNX90sdVfOVl1MDmwmiP73+4Uu5OsSFj8jXRBI+jK
oIsd9qnWov1vYh+D8Z94j/gkGqwNXvY+aQPaXkG3CRIMxGGGGV8an6Ckuuj9IRDb
dWRWouiY7Kvwgc5cYiV3/TDfRTh//EL5ONbR4NnhxdpSMKcInFPXCadSvDp87cyQ
Y5NnkLiFzgXTwLV7OBfRhfHSL/6IdWTi8u52MX3M0BZPwRkxe7s50Ww3pDRf82g2
0pWf8kWiXzGD9woA0J2kjJaTI14jInNQ5826IkxVZ9vNBFwA1EzlIUGt2TcPECLB
GFxY1XfBoGUh1le/lJWA0/Ey/2duGG85DeqK3ckH00/YexILg82O/Wl2w/CCHq8+
3Mr+5YJ9Fs8Tx5JeyAX4hco1Td6o8bsKZln9u9uwmhtLw7bJ0ungkyNO3SDCsjg5
zZmNV4wmS8RRcMYtbQRmhCSlWyJjxQ/ol9IXgKHXZtCCmo4qdZlv33eLBYM9Xd5d
sW/NWsxtDRvGp1qS4w81vXEnv45haK8lc1V7C+fCywF7Cik8bj0jQir3q8r7OCne
`protect end_protected