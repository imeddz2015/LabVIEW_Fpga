`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 53984 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/9huKRhRMtvnNqb3Z+UU7TahEoHV+T8U3P3ufru7l1O
3DlgtZzb9QxCbOjthp9+wDkjygH0eUfDrEl1ovhZG631oDlpzLEajTtY3bJ2d1do
4/m9WXxV45j7c8PbUG2F8EjER4dKHLcx3MX7lxUBCC+uF4mJbdFhYQBBwaRkZM70
OrRZysP4R7o+Ru/f5WlwCSzHsZX5yWHRzP0mowwA4YE8PLL1ugXlBbHMS8ONrdrF
WDZW2hEWjA6UwrhqMeQkH8jCBt6+AomLjNY/MBySDS4b/jYbJJd+x0H7mbzQXM3D
yM7fOQzw5/skKf0u8TLaA2I9BVv6I9/tqyBu7UVYYPLWOo6etoIlXOybLFzHb4Pj
TRBpc9pmTqVt6Cg9ooS4Bqq27LJqVN1V6uCce6QxzAs8zDgdfH08SwGo0xGLhD0/
oO4qFPsrRRCA2plRZFSYtzPWlYbnMMcuNqCSesVi8q17Q6/Cu+VrsB+aSF5gP1r4
1yxMZtikfUMKpHfPilIFMvKkvR8txjzBhm5IdRxsl3d+3ccGFmQMxA9TWS7HfXRU
9N2fVNzB/YohhfFYeScyxfkkpQgXIdJZNbsv6uC5pHRWoSHYu33AvtUKxzbt6zFQ
n6VdZjnHwL3yXqfeCadtUWtwg+lu0wkuNrxJWgG6ycoUVkm27F3fvRE++qmGKAs0
CTogbG8ZXUPpKDwVZwFn4gCThn4Fz7h8bvhnKErbkgKe5pFC2114IMmevksOZA2c
SqS9n5xC92m/5g0Ep81Xwko9Epe3VqS7rWpk9+0UH5a6ioFG2r4Ezb9xJ5bdE0YR
YkTgsVKtC4Stdp4M8q80jaox98gDI1ACb2RRBo3g8Rp3hVEQZMhqLFc0J2VGRWvk
6/TeEWRzx3H+2Kcdq66YZl/cVSYxVtINDb7qoV/Yf6IEJ1MFQE40QUFVQbxz697c
Khdp2Myy7xtcQBXNqPA2LpztziRSBa9M2t2Caod/cefMWLfm+pzDyXsD7BqrFds+
HutFZItqRrXPIdUXgJ+d8lDd6vtK5bZI6w4AP57Rp5dg112qPnHKu6CYG2uqmbai
nwArGDw8nqskYbzed+/KAeBdUGFj9PR0nhKguxJNBBJXUju4b7nchDeL+hIiEgbc
7u+f4Ew85QmO7IpRm0J6cYhtwqS7X31+NV3EZFtVkPuRlP5KX4rajT46z3HdWvu+
OsGSWI1fBw4WoeqnbJURbUzj5stciQods+f7JtEyprm6b55nGsTqXXRJFRTfUuwj
gzAB9tMvmrRZ0E1UvmR+hMtcr7hvL12X0hKyubsTA7ylrjx/amivNnyrv7OMyH73
CxzMSiaamYkhPKPoBGXi85Eg3vQKu4o+xdR8NtxMiVyNLQMzZYo++16Ld/klOXHe
hvpzQKwXxctBzNwqkFwMQvh74lMKfhEA6a8pozlh+f3SSo4sIwtHMfucPs1vG7zG
LV6YtjWAXh8nt4KDJWfT6zW3Wc64JfvTMCiHwfRPhIb3wl4Vtwgjc4C+UOpmYTVX
asZdMpYZW4+ORzPsqt1tAySj65huTayOyp3NtLZTkUT8WgH/BVQ/+sFAyyBY76Z9
hj4WzvvwytCUbOOUR7WLAyAG7ZKxpr+QhOaQ6/DMzlLj7B0cM4oSBgI+u1mDQ20g
V3mBdIiMnFrNdFLpL8UcF71BiWqktp/ZgjurvfXhbR1ndZAW71EcFCbfwU6cVicL
zskr78XIGruUJpzKF1Aonc9KcxXZ46EnG4ZZY1K2bhG2gheOSkB4mK1MBkNvzz9r
mDPb+CzCkn9IKZrn8WhpX27ORAZ+foygi4PVf+NZRg7Lo9fhMm7gGLHqBXvZFQNJ
y+joLke6v0497v/sLFLqJiARtNWDGvSFp8cn6v+cSjuOaXseJIPtkBQwz0DFkkmA
8vGSCXyxH20myulH9gJlsNvZ9fdeu06nhUl3m5Al0kcIxNp90wileQpatWVKpLfT
IOZc7+GqTqZk9Maq3Vy7fAVgZGQI5mFmBUsvLREQTEQWMn8CzeNsf2ttqq3LSY7j
kP2PzRGnyKbilWKc2/CtVtINdYdT7yoS9UINHTbzin77sP3czKAt/qZ6MUVKG5fv
Iwt0/OpFCI6bU4pDTTnWqXDvD/Ql+HShT/TGXICwRQbvVIse+0tb4HMcqwZKU55L
XNJTbYK2N1GCQ9o/eztwMDO6JqZ+Fi0jgtYGiB5T6dhX7y0pBqT63MA9Mpl9nNTY
URuZTx14hwyhv2SLm8D8hwTIM6O0QRQBV95o2w6c/Oa77RntO756ji56iY9a1jD4
07sFeijzoX4T80rg+sT6/W1a5pBVq3yf0yXQMztygyqmi8kZV5YUH92BueXuLG1Y
UzMh/KWw6/2+g8/ZKrhopkO7voMcBdFq9RRDaecxYFc9wyGNbjuuYocRMhsPFfWE
r2ZvcrT6zMEJNvT/t1f2YwZJmzhJGsPr01GyzRsxH1pWKVHBi1Lh61REsrdYiro0
QAuneSuH3jrMRRmZBnlo6GV0eHyQqQ00NDWnoHPqEW4U0JObKAT/KKILusqK+zK4
QDaaWGaEswS0MHds5lFITyy8pyyiJXi6p8+jlT3yZxEb42a4bW+8vRj78DRSYwtw
0Wuq7T1mJ7jIjASjGS3SZVT5pN7927T6vYBiU/BSJWxioh1fkIYQ1Vjx4rkBPjLF
FQaLBsBcvMKlkQlwGvvNQSGR7wtRFOjbKCgfyMD5LkTu/Pt8eOKAB07fJ4MsTEMa
20jkcG6b0tNMBvXUvHig6PgVcbNu7uXtL8idcw6gbQ5DgrhiDxf5iUyGn8Zl3mVq
0TCOzfyQtJnYiLGXeQRPrEWH8VbAgaPtN/ycpyVtRMDqPplmiz904nuA3Gv9rl3h
rlx/Epie21U82FNOAScU64+9yl2TdDH1LLiz5M+eV0hkMQXWvDUZvDNtcrZ1Kn7w
gxDM8SZduYGZ4YeyAS3nsrARM9s20/p3dSMfCabny5IzIpdlRR3dc+RVGroI0xu2
rwRssxpAKZX0NnuEeZfPyEA6abI2GW3inKXqDjljTVG7YvkXtk/uAJCciRrWYXiG
hdRQ80EvhhlMcXKQYreyntZfJX8iKlRPQKcPd2KIHvWVkd+xub/R87sYq+j8vR0t
xHJgPAbnbxCOb6GDCAZF9au9xYo7GauZ7svC0XoMwvIqOw7mjyaafI85oZx4HNXp
8B0wdqXOUlAgh2knkF2hWCkivSupW1M7qaJVsSGMuF14Rjawm8raYK7Zcv1TiRcW
fsFFZ40mnDKgspnskabMYll5LGm7io8WX+Ulw/VK12NePNx0ZlCVDY16oLp0WxWi
jQmphaTp3v7w2EPQ74clZlN9wMGdc39RPbJMZ4hVap3cn5LrhfZaxgZk91wbzh4T
JVZo5DdTJC2n77wa92L2f+IvzASt9Mq+DCjbAMZv3lvJL1yuq2HZa/H7o/GLj47K
ivPYeHFE5vSRFwfcFm7+VJvqUZx8TDKd09c7FxyGr9TM9FzdPIRRF77JE8SMY9Z6
SgSzwvOasTZQH4e2AWLQwaec81oQE163JOSiY1bKikLc5T469vFKlAICLib+k0uF
3nysWwT4p1EAETlcQLOaGPqUS9LfVPW1tbeEpUI1kgIl12RGmQebyS2N/DWFmLsL
OXX1B0Wpx5pewtzN2VleM0X+V0fo3CSUcQq9MDNG52EnX3UlRFgHnh+WkJ8tWV3h
Axmk+fj9D2IwRO65Jj4qnymcWtLYE5NVwHgr0zls2Lrk4zlJoGjqfzyij7B0tADG
+cjAn1kShRu/w77EMTEsDrLH393JZGrVwTRqeJDzTqCUhCA7iNJLhPlyBwX0cHYO
5hmWeoc/hRfC6Cog8oaBlKzDzhdUzMNg7dhS8/B6ODLKGSnEFm8b+rC+X6BEKwCj
+t9WQSnnZDZY4EkUjpOkbZ1kou4ySfdf5x/HRIeI08Gl1IEJ/2o626r9wT0z90zl
NUUtjjHtodqba0RUFMmbYpqZaPxRIMeJCBYs+A7ekGnyqasDvT0h/QWv+xmV/GGF
91LXARbkP9iESkZ4rys9vAZYy7c2gw6TIbPAMD0OuNbFPmteTWCLxIM07YZJmIgN
z34njYPSMVAN/c10pbh14TPZYA1uHdiewLv47rp2wndIIfAoURHRMMyt3FK163s+
sv2WtuGI1Wme8Kiejh4PoxoqxHr6SV4RSnDVpFsFu8ghYsCDLr4H1FrG+NlhA3+Y
0CW6wEp0CZXuj15jbilaiCqDLw0mAb1pvvHQlDPsQNJ0yKHBaOlSPtrGvZY2NZKk
rh4qE2nvcj8a73CwymEKmKQUSMrlAtTiWw/JnOhFFwFxlA7iJaM9POOrUdix6J+g
/FZ35o12w3PtVvRV55eZduT7qLp7pOS2MYGZvehxCw4NI1WpGWaeeB277uxXYHA2
BR3VW83LSOOknqKiQgnitbWtofELu0JbhneRzaGrzt5eIxRj+G1bo7qbwF8Ey8QZ
lcXLrgOF1NKHTB3rzpPvwhr2u++dKQFAR7eHzj9wXFyt4zTBMTrd8Ly6i3XfFFBX
DR8JkfbtU6b2VZZIrSGbEHYp77buP5LYQ47ssu2e1IPF+XKOzuvuq0APrxulDXCy
L2K/g5luWWRiVXZ+ArhkacB0IU54G0bpOsQXUO+zkHkqhL/oixVDDU0uVBCu++X/
eO3vRcMc0lA1OVQ1rbK5Sn6v5kwfequGOCUc2j154lrfFGY+KGAYJbyia3hxGNJ6
YTEsb6kOl5uvy3f/os+GdhF9r4zpVV5C/SESUdpaLZImLlc3Rk6Cb55PuJXXBKsO
7koG4HvNSXUmDb05yuNAanmfl9G14BVKIExOQwDzJ4sMu8v0Gm1/t1N6Ra5pkeDF
dJGiI4vNUVdew5F/p6qXxreg1AibvVrIc3vjU6TjLMfF1XYOWrJzLNdbPyAJwBef
1oV/IjJQHcrF+7YFan8RydmZUzCfSRXU7uFnVoogSupRA4Q6+38gtUvCDzsu/Uil
b3ScU4wBvYswbqSwGjf5SLgIpnDPyOLIIlQPczJCqQbOimJybYRHf0qdhtPGX6Ap
0R6oBNiKLnF6HjGxWXYpWSeIGKP4cIshaAFie6Nc2hv19d4RdxP86eoRuGx5+Rcd
aqTX8imbHkoapbanzkZVa5pBnBsTj5ObrRnOuZkd0MFXW8DLDjYNdXfAx06M/QJS
u1nMLo0rFyl3kzYvzzO3Z9GbAPNhIUSZ/WxCh1F+FecsRLbVuzWvlLrbqOqxVPev
Rf0zB+dcB0Pb7xi0Pw1kqRbSymal31snSx6ttd2RvS8aJdJaLusJph0eYsm7MPuK
zHbgP46TqMuyKWHeeTSMiRip+1uJsvemlP6yTYOKl0tkQm3HQS8nYDc0Q3QOrUkp
/H2LHxd8brmMdT/BICFDzE8JmiIvEQVp2o9hHs/DzEwSga5VkJvzdPjh7RGj+b3r
pqicghhiFWaPsePBpWoPR4t4eLRpumuWXli7hhBF9ahFAHQ9LNvIJ/e5SHunr/0W
+MZZ+wocMPyr8sc/lPa3GZXf667xovH9PX53jCiGS8n4SdcPUnzAx1Pqv9c5M2RI
751DWSxvxmmKhDF1fju2JFlidqrtvGYRHRFAFn0/K604jLLohLeGDIaJlNBIfAW9
oS08hWU21ekDvQKYbSkFtJLZUkA8V9Dt31ecrv2zAIAPkDxt0KHmUBQ9mfkZa6aw
UkG0vhEjVDXCtxuVBQb60j2Z3iGwU5+3ddEUk3y0/GdjQImA58kF6IQ0K5VgvHSu
muF/wB+L/r5IifhL+cmZ1f4COnw5ou1JjxOzbUkXlEEiU+u/RgUJFlIHrepL4m+6
tA68pgkDFg6xLBekXmNIafeRSVTsDB++f1/YVy5C6K6SFSNYo8Slt5Rj5kdf13tH
sgU897bq6Uq/CZadBGSWywddQ/Fv4s2FeV0G70wf7KHpz1WMn4aTUwPZQAIMvjiM
UdY0DSNSwTb9YzKD2zYmDd6RYIy+2FF9Kc53kbOqsKtjUE3B0WoEW7yIBRIKekZQ
1ooWW/rHcWmkxpEPKLKOqXXEJze2PPeAAqpOamTHv67+Hyu4Ef7G/+pGq4UL+dEk
fBvDUkJ8lyqQuKsy3jBhYlB7DkWfpHMyjWpERR6d3tXs+Iy3xXXV/zSeNO8Goms1
JbYxJN/nl16wIS+GdUHzLVVl5Xl6bgpjz6K6X/UzadGlsg8EnyYk4lgGRfYGqTzu
Td+Zr9fXKLX3COWMlL3vLC2P45XWwhCm5TtPcpDjiwBn/lLG6alfhYzZipNMfWsv
uJ8VFreGDBXmD3+SYhL64Lcbh0OrBBu+SsoIIJYH/1v6n4I8DMcpODjF/+iZkYh2
rMg+z27qmUBTyqjjwfFyTZELytGavBUoEF3dyvoDrXopaFSExXOb7gFcUjInrwSm
iDfHs93rqymm8ImbUnMO0LZiKORQhImPkrRqfkZATwF8BW1m2g0l4YtC+/1PyQwj
obEwRIEMxJbRI8ArJlIBbdvadh77liuWSWu4v8i3Asgju3bKQZ9ZMjCIPDoCJuFg
vJz2CVSjd+V0C27Svm3LORvCaflmC2MwQ06zHWyps4P1Bl/jo9UKMZirxkc23CwY
/q75vQT5hl7CpnbJty6jnh9xIoqDvX8vpaGZOqi0QN/dKNKzh7k6G7gdIWSga3sC
qLMSyHZ3xrIZW7aI6Idfqp7eImmdqACldWOydUIGqkh36T47x6ZF855Osp8LpJph
9fT01XWYxghrDeAPusLcXtwA8J03/7O5iGa7l0xX9cQNSCAcRLNOV+2PttVey+Bj
9Ta4GdU/tA1HVutuX44P9tLm2OGueaqiO9CY74MslKUPU8yRTFzb2AtMgGRsAn2a
/qc4m/R/P/ateVP8qLkZiNCeG6urmmwTrVx+p1jOwYk2j0sglIcIIe+3kmOLvDPP
WUlbYqvm4e/TI3qKKbNT/TzdE2Wrp+iTlSVGSGN1eGtv1m8I4GHUIqvhFx7UEVtg
2KDAuPwM33aAvJD+cV6JqJ706gX6kIz5iJY62LzTPLrJhXkJUp2j6WrUBgig9DZ1
6E5vj1/vEMYI2xi1hNJ8IeoUlX3QImmAMVUmeD7fvg5CE5KiNlgbpi20cv4uSkzA
vuQS7V97tTVv3AalopSronGK7p4cEFugmc7qZsy1uIdC0WpIhVavLi7jawMVVsd/
QFWrQBm1wSH6wf8aPkER+UZcbM0YT6R0E/I5JNafloz7LZevkGTA5Qe+ZFR1VKUY
H/LlJrVknFts7tpIYqOHds0LfQgcYud9ESLoLZlXxR5mVOUG/7uFioHmGoR5FsU/
X4JODRslxvCiod2r7wCa5QsOtm+mKwUTbh13tzpjKN9XNKBOa1HDD4AChxnXc7/g
AgNL+Q2inAuCZ+kEND8PTDWuB0n8C0cXwzM48zWC0xH0mCJ+IJZsF7tWWGTDU8s5
aJov7OMkNKviLtX5N1PURxNCiP3i0gCSZp7FYntBZZjtTWTIKc0aMATWwWuMgKZX
Fi7/ZlmKFaG71We+XaZ77goakfQdXqi5BoAV8RpCzzIE+pa3k70dJDYPm6Tn6eLF
IUkyiYxfj7sDiUyPpad/Aaxs4xUNkaDpaY2h/6uayOs2VImMvKcDG54ILoSm9z54
TusAA66tuGERSG8HKqU8JDQ+ifugpmh4aWomjOqsFGLMDTxzqPOb15y4NHf3snd8
2XST0jP9pzuBb+MJM0EQK204GSuI7BBB3yQnyUv6nF3A5sm9gIjSD1LAN57wQ/3H
W+4wo8hb+7vXE6otazlaU8brZM+ikE8E7ECSs8vBZDthQxisd7CFEvg5I4AXNfaG
Huz0dGf16pdJgkOiozgaVZP++r4skf6cQk3tYg9gMGgECpdcQosemEKvxR4024EN
wz/sUsRAPYRr0xF8HO5nai54vurXvHvDzXlaIlVUj2Bxu8bIWdy9b7e6aWW9k9oN
xqIpwuBH2efMK6q2w8yD7eMx9DRYsiK2JVxmpQUAmWEMV61WE/N04DurP6iLj/R3
AVFXmjaUU4CEm2YNf5oeZMxUw/owGLAGCXMnlYz0+D+HWPzi5uXCjSthejv/bU8g
IShB68B3FMzin0Wpt7rbjcojtp8s8B7k9AifZktB7TIcVdsy4tL5d9l5xfmEFhhv
GYrhWg9/3EbxH5SfTiTL0d+8Posd0O05hbsTxPHPeMxamaXDNVap63PQ2CTrsNQM
l5TjkN0fCt0G/aNfNrYHluY8dJXC3JDI2CMU3Ti5MnZ63iim8f7Vn3KQ7uHMfhzD
h41Vkp8WtYOomoE+trNhI3k6uGGHkq53qCoxTY59oSYLW0WzKlmadaSae4o9bDVN
1lMMarvU9uiUveibhPugT5pS9KbYrNRt1tWEE9uSjsI9HvHm6BHH1dX2JPDTbLHn
D0tNFnUBI0PVuK5ownPLlCA53lnTE1LtY1hcXI2elvwKaV0GIWLCVBe1yTzFgrUM
wr01W8eUwJqyATyTFOlTchBRUlaOhTmv1Mhz5fqP92nfM/PhgCJi+gLPszt8QTyp
aWhdwjx9t0APVxmkL3I85waQd/mARF4okT+j/4qxkuFnXj0srKVhFv/UakEMXOSR
zjDqoy79sVOCWQBrn/QLcqxlVPdL3pQJZuoguK0ONM9Ak5GrrMi/H8+Y/t43tpzX
6MgBfilBkuKucBBuG1NJEVPEHw2Q4IkZBzqrNshqGFHNyFCOft0xeFzQ+rV0sNsZ
MpvejLb0XsiCpYm057fzsgGoMAoTAtP3EfkG98E800LUMmfcjuqZYpX811aJ5SYm
m8qiww+B9MwtpVEOzuREVODHhuzcyWqMIxoff+VlszLjqMRAjNELIpJN6z37FXdM
waPAI8FdgJOT4gkqovOT/PG7QupItmgGyIcUgedV1SHj6J5Th7XVNKmh8ln9TDFC
Rku6lVvbtpXbhgMGabZvSaCPez+4FAhOr6OnVhUjUYVJiY3TbrKLsghfmcepa8nX
hDLJSWA8tS3c07T+KxrmwCo16g9pLfFYhxBBNmFsBIqYxo/9kA3voXyBhLJYFlhl
dg0/IBdQz51robGPGHVMBX6NjyKWGCxr9MHkALfH5GY886USzmR6BGtJ+lwNUJ0S
vgDGEXJtEUBZGX5ejCTfdFSgZdZ3sfDzmFx4fs0USa+9ybcJnJ79UYk01QTZK8Rr
umyYsD8XdQDq4rL04IWmDhZKq/QsMKV3kV+ySRxM8xpxitej+mUEOnNS9K/CXgql
reU5LMFSDw/KWr4HIHElvdVlKpqqth5gx7ZN8NQ33E/0gpsnCBQNeDlSTjbPkWLu
3pJrzR13Cb3IxMCfBYx2mD2mPZhdMjqiU8DYZWXHv9na76W5xjVsLlGklWvVAUeJ
Zh4SN3GqUrAXqNeUrpk67D3J6s74uJsRM9eVvUHsi33H/gz7w/VQA+TTTLekjfo2
nYck3LD3RsYwfx4VtpoLpmyG9Z9cOv2dIEJLfLkgOU9hZ4Ir1/JSxlK3Ql2UKClC
nyewKyzJS3H+jxX2T8TC5IYMEqK2gZn9W/DFiR7LF3ekGy5Nu1WFxt2moGPx5E1F
WZ+nfsKdp36XMYc2mxZy+N+KZvIXz2mbG6GHg4CkfYHXr+FtANKoMLwy4BXqJfVz
3AhDzcWKGKXfLz/55S90Zk/8vM679hugLafe8aYTu2jSpKUTQf91QkK/EMm8wMyx
iya3FdRcH7JCX9Q4c827+B7MFBqSY2yyOAtOdCc28nGpkHdhiB6NxG0Sc9DdiF0m
sXRsxbS5dzVM8x8pOruk9ifnHX94T0QFnjUcvBchnkFKwdGDPqBPg7byE+2ewKJe
L4Dp2nARQqj8m0aS4Bsn4jfkSs4pCrYvGt8XPsSgJvdMOA9ruumaYxHj7gM6tvQ5
DTv+wivnhrjV5fa10QmJQFRMu3cr8zgzu5xrkldLiZLhuNc9x0kICs+dlYDXmOjT
JHwMchgAgEAOAl72dU9wUyxlF2xYjPQwvQR9lyXCTgC7gN2UYUxIPjXoqBfN5yx2
wJ7fxNFsqLZUTgrzFJjjoDHtvCL0pxITMZ5DFEuq+bh5VU/gMjg0LLQiJt/GzsFt
bk6bIEE9x/yPlf9tx0yJCL0A8WJjUl1fsA99nscoPGy5u1KvneXlA+4jQVicq8ye
mdCPKCHNeL135FrALMRqZrLtGlQHxrOFNhspdusvhLy6WfvOxcf88jQXW52xUST+
GhL93OSCO5pEnuV/ATyFKAtABU3dv4OuUkmNZx47UkStNVmWIqhV96umIP6wrxw5
PyelztGdJQ+v9kGo0zLBwQdo8AHnVj8K+GLj3MtC5DGUMEbMno2uW6VVGHC+BrqF
CReFS9FO1qcCad8XhSmuuavR//Xpbb2hrEmirO9BMb1p8zqKemaausTYM51atSXq
X7i8cSwnSC0ShipygJWndxGL9SET1f+EsrXMMTOpv9cPlaBGixiSeKHRl6nMUmrY
AHU9zcnaDI4UR8Vwt/rlw+MCb88/1NlQz0DzMIbHQaMmOvcXPG8hsBFAs+u7h77K
WMj6CTz1ZBaWCVVbchIr3YyIDv37z6CRaMOXehYndko6t/2rX7ZAl2/RrC73+zwM
7hUJI7sTGT2xnMuUSSQh33HS0kdzFOpLv+D2fWmFDUpB3IRe4PnzbHapa2tivmDs
v7wCSFpcLZZffnhylOba3Rz86Ph8uD9kvftY5i9Bytv9s3l7B8onkXSULhDl3EQi
HxawKcim1tqlfeXwSj7uAQmeloK9P9W9KILer5HSaocux7GE4Y3snhN3wa/3iV1f
+kg+EBqaak6zkB8UR7BVFHQfWXELnL3e3rryesRw9Bm/wTnoWkXVzQhuW3XwJCfe
6pzEqgwOdyWE+FsGYnhDYuDiiUFAmpND20sBEFv+AQB6Fq6C+pHgvXQ07u+im6fd
Xzj7F0ogg4U9EMVBXA0dxwlQ6n+OatO6Dn+bqbspRyhF/08wh7k+JRBYwcRhrvaL
0ITCbWWm4u/2d2wkai/uKw0quPfPg4UBtd7GEEviYxVW/i+ZBYS+m3CibWp+OWAY
sUyw7y3D11J9afPf0zfZmC9E/ThusGOo8jvzGvPSKRg7DggZN4utVvcH5XEHpEjv
UagU2XtKqZMGbtMKCJnsL0pPSfBWk1/b1V7bKPmOj9ESdvTCzLC4FjOiz6zBncjt
AAmQQkftKUpaHXo/VWZFUSsuhZJoEsO+5kxd/a1HaRvUooLXYFaW3Udg6UdKkqh2
EfytRTUww7vZZD3Bt+mBx7Rk5uusmNO63QPfUI2SvCXXtM0ckn1PJrbn6VSyLLEj
UMRxBFP33pcVQw7vpGhHy054vhUjVeuAx7BjkpAKobamPPZyL1Ei7TqrG95BxTLA
7O2BHpz/yOtjI9ZQBoLVB32/LdlkUO41E2SaHuHKcAMcOd0SJUT6Mw5Rw6RRyJHw
fEK6aKqX4NsG4+OQsw0fekNGnxmvnKIXU46rSAbGygjUHugzAdFNQbPA5GyMWGQb
gTwj9hukwtGbgznBLdzuJeXWilv1XnR1N8Pf8N+fETFEt1I8cQgHpLLqL+gljPqe
VPQTSRhWp8pWwDxFJ/J+iraeoNGqUDWmZmp56pxZESyi5zrrFn1bHo4lBLfXI1XB
FoeYa+5huOWuUe/zOhAmnPmR2eBbtlPj+0Fup/SX9woi+727yuD2VEVqbGqz0Iky
FSXl5CVnbCsgP7B+ARCgvpV5AnEjGvrBoXmB2W4gPBUPvzrocYt4F3T01HazCtam
xmR2GCIOFdNrtVKreyiA9FN6zOeofqARxuhpD6tW0H+RAm7PkxKJKJ4g6qsv/Mq/
Y13VNfXnyR/2Cwykg9dOHSU2ougmVlw82PJfXXkfJOdsmOhXKlAj9Q0sGOMUw5xY
F8Hr05H3xTBWBAKkBW0HJ/Y8Ucp2pXpLEI/1mQhL6KKsn9mk/nPafBnzbozijwaC
tOCyChsRmIyjiYnUlbwWLpLXykJn5w+h6FD9bIDIqo8ObCzkDh5V4FU3RCbnMTHB
tVVEWmjVSNJP2Af5FlLxlsE1BYRZIzDPhNCyPi0X9H7QiTodPQa0EMlb9MlsSj/B
OCWb29HcyMUPBK6Beqev9SH3/OIWP5ssAf8jAq7xg0c1yYRxNp/Ad2gJmLWReTCA
0RTiOt9atnLHU5lit0zeJsg2npdLmfthup4S5pUvYFWql1SDSwYIm4ZS8MPm2off
FirPrYYwHH08wniwbamNlfQnwmmhDIyCIWCZEb58rlmY5lo5xDnx9QDYZch9R7Hd
mhorI7X1TVvEvpxJjoQDflH+iR+PiJj4cde2Rj4NUvdVI8DUS62ajuD26meBOznu
miS6Ba4e/A6Isg3RN+zGJPXz3c850wB3Zcchqrj3dubCKpVc2YOa2+lCev9J9bCt
l6cdNP6CKiEMl3nvYUTUyiQwL3diS1f62EJWujghKs1kSL/NGPzgJfbCq9lGGprg
aE4gdgnP8T7+hp0/b+CR/x8sekyFGB0Cc4T3JUWCxAvHM+YrQMeScB4TigHTpFVA
2qLxTFbRC8/WnjAJ6+OrJA2tyih15f4V2I5YoxQdPpE1n55ckokbLZ5XVinQDno7
W7AwXgwKjDkzzWHWnaSy6o9BGTh4eD+Hltu6fja4bVVn9O4ZE0sUYKaINFzt6+dV
zuuw3fNOPXGzrznJ5Gii2epCa7AsGLB53kgXbO0Vg3OgA+6Nbww67O9HiLKf8UME
FPoHvaqr9e3JiH7SpuQBuJiiXlG8EEqb1AnMVy/zRtdC0bmuJ1TVkbCJ1indsMRf
XF9bUBVKuHhjsbZMvU9Tl0frv93KjaOBLtGlxvaKxww9DEcMCnYCYzqQOPyBuOI7
s5joKH/d09y5n7jQTlwl5wQMSlemksXRJH0iVeb9hReDd85Xa4cBIgEjSwXN/wyG
hQuwmYbKVvoinEtPP+aUVMabdxrbE6NXh4kFed2CSRXIEnRmoCXBpmm1c9+pZMsN
uL1UNUUS7UT6xRxsQ+EWwaXPQBiSyIzMawy8f9itIWTH9L9PvQ9QbyNVoL7p1f/0
yDueavL8gfFuaOkq+/dfy9FuAJ9EVxRQOhrZRHq8r6qnPkLSvSXccDyQJZhaKFhF
nwVqvobP6R6suf6wjcWkyQZYymsNKz0Zx7NyZK5K31kH5zxTT2HGivBHgc+DzbjK
0+f8HWtu4wJ4rJ/7ORhuPBla7E3XyEuZfe0b1sn79Q5R6tQSLj2qa1G0wdHFMUW2
Jq6gpPMY3Bvqwsyp9ZFOiHIr6PyTkL/U8S4hDIHnzHipg9A3lCGmS/BNRodYJboo
X0y/WD8yFOJqqTjTfOw6wA+jtpAwTxu/E9iLQUZ5CyX5E9c4VyvoHrH28GCL5Jib
qgFbUYrmWgtVzzTyXA2BzxlvjkuZzT/NWuFIsgSUVurr9BxsJoEpufbJycYz0t/m
W3pxA5qAnpfgaQ72GUBZiBfjE47TFwQMRWKdE1BqaLXXcfhW4KuxljlYnrrmU4bv
64mdJk7A2zGeU/uxH4IDovsNksmzbFTKaBZ3HU7tUNGRNlg8C85QvQBlNJ0gREWG
GOQAAs4DzwdfDHw4AnG1LPu9qHDK7xLSmiPUNOT5nVjAomnvcqmCCEqxIXLznbyb
XketEiVc4c4WAqXX0kCPXkUQMCLL/TuhEi9G1YfSE6L6kpilgIm+Ep0KNqJzd6EP
KKSkbCt38qOS0jkX9+k19/QYSr3WH9ZmXPf2umMSHbpbd4CNg3ZK9AoQeQhpywS1
p1YPnrDU5ekRRFMRbrxjZNEk1TfVbLgIsgOTd0bfTTAyawyzyrmaVdVFkL6ATjLC
Kgc9nHEi19XYaT+Hi/z2v4wtT/baSbMs8Ub9BN0wBo/xyNL67nz1R/fGNE5OKTz5
M8wU9PTNxpEkLcD1NJxueeK2z3perEI25pRIzwHU+t4VF57/v0f25TX0I9n94MZM
+77JO4OJCOhrNRbGrR1XGkqr/vc8ez+LV1AEXj6ehzb6ptcFpYXPBmetZHeI52wW
1fnOycOPNIpfNQsSjYOXvG2JaiwcBO6Suse0ohd+wE+1inekoNgPxO/OsbtqRz3o
e3fQGfj/6CTYE3fXm0quXTbcsC46E6ic+9zRD/RM3fIDY35U0+l6agOBK95eorOR
SugQk4H7xNUaG+d3+HXIdDe3DuXjZeI1KFgpY1v3QhCeKL+EAUmYPkgt2PA1mawG
mM+l53EqQQQsi70ccKZ6GejSqaEC1QKiopksiRUtRSwkNN1UqPJlz60G0UmWvvQi
E2I+a1oGzIu3Kz8kIQsOTKj9r4bPZ9/vWqFHzUX81LHTdPW8XGQimENQWoHt2u0A
s4nSphub90xtp9J1B3LKbRrRUAwzTc6M+VSCzx07MFJBEUs6r9SLN+Y+5JmTPs+Q
6bcavhAy3YE8KrYFRoWfQHiL+lMhHCy5HU7xfjiECGb/GA9BdauQKnYxPsTUgTbT
JSi3DgQIGdo/Yl/ahd2h6S4rfiPS2QQ+WjtTXJjY2jgVvgxx99xJUZGBTqDl/ooK
uXhKMsDt6DkuGvS6Xoz8BLZCCyAq02I0P9FlpQLtMqudI3fSsrVbzPqKeFQock95
qhvC0bjQIkooXbw2hAl8+ja0VODdbms8YgfTy7mCukO1T84uDmpGEZFd9U1TJz6a
wfOyTS+eCbNtdSveNHWLPc2mRXgs4fnvh70bY7IGyO2RluKsJLCcTYw94cMDi1iZ
8YceUgKOvt8TPIlFhdSjPgPPxIYgJ0VuERHQSKA3Sh8MUXPj5Fs31AjoJBZm47XR
P/Tlq7ZqzPrpaKsmRPkwF/kkm/+Qc+kxFIgeL5sg77cRoPSJJSnG0QZGXzqIK6gs
IFaeQopfwaFDAtX7JfygVZENjlJZ5Gcwyntflclg3auBCrf4xqAR2q0iINWC3jdO
otpB+eAIVSfENVMXFPaQojVgO/2GjKJjUX5PXz5uMjeliYDLCUOz4ETI+SUSc54U
dAebPABnU/qRY0UX6m295DDMe0UkAWe+cFXrpIOrlIcjWRgdpi++O6eIPvWINAEg
FJPbB9WaJsJRPhC5W/KkVcctM1Q613YEPg7bYTNo8hWPeCJ+40IFTHAVc/HcbEUs
9fId0RaAXCDKki+v+7IZsmDbY60aXKNAk9/gIqfaY/U0blSYTfJYbRHodlqb/5Ug
smZw+mC61yN9oKbxa7FS6r7ODPpPdfcJWw3AdXwsRhPBF0ODHDhEolt+IRoyaeW5
SOrU/pdaQr+4Cy8gS1CuTcqx95un5JIPorwlBnXodv+xb4BcXHast+E74/fB7Ey+
TSDp9N0wrdowTsUefKvgv0mrHP8p/yPHII7EjWvW9Ir6iaQp/Mh05fuBuVlIEHKZ
jUBD6IBNPJDrrF/A+ZlAHS0ZLC2fTbx9poSc8/Vqnl5ZA/jqfw9bLjDkTkYQM0+B
0dQzvYQMocFj9jmI99dWhFN4QkTTWsxnyOekoG+qAX8Ahft71gAxL/YZ61fciGLm
ipnLMz6YXFOCVgamu4nKRp1pwyMjA5jTCEWqHvW0shyPLI0Tiax9pvWhoB72xskq
RnX3RMgSbIsvcBosBJnVdT6SPq7CqMAqxKFJmuVsGwWcvDJ7drHkp4Zh32IOmfks
NXypRFcF77sMdtc93p890yXUNMQ86QdRM232zSXkrRi7zGvQvbrnh078qhGQFEBe
KD3SXkTepetZzdnPoySgfTLwBdhQ2othxyJaWyqhYeFbMV9FQnQe8X3HAjlKSCSn
q4hm/OwOtz4+zbciDmsxieiRVYcQarXkQFXm8abKpRHcWJ7B1daa0avnN2FdCHYQ
fPmhFBQ12zgbWRtlSmXaSSdPLXwqzvmz8QqUm3D6VXOGpvRpDbfoa2CDiUn1aN0/
u7CIe6Bf8i4VsxBJM15DvxkdYhe9ruAeoEPQoJQCxfCjcdLC3CU4G2NxHaqpwO/N
HTJf3clUiJXaHeox4QdRy3yL5PfIqg5jVXwxf4bBSxthEKrTgnYghw4I+++2mhg8
lIj6mJIyyUVF++lylymvI9pKOgs9Eh6UQckZpAhZptra5Y3IoR3wO01WiG4aRxIa
V4DxrA7YUknUpwuwwkaAaWHsLjk7xthYB8hUfU2aLwbvyUTP33/3ilVREqV8VORl
2OHnXKDHv/BHeknu9UQPS0RXtFjZLeWbMxLv0wTt4Wegc93sEwn/H5WB/z2d5qiW
0CWKZb8ZIA0EBK/6SDgWqMy1CTz3k+/DoY29ZeJq9Qo3cEzmy6Scq3xo9xTg/Am4
eTJFmcZqW6oDcoNsDIWX02diAAzOxbinGdSlPUUJyrnD6rWgrqKbta+zwIEq4yUn
b7gL93LcFU7oyr9/Jvb7OEH4UxiUhXE0eT2HNGuLFbAOB4UwBIgLqbcKSpdPecgb
xxD2rzupVrozENZWZUT5kFKoCuO+avRAWMO9PsUKaZzGL3mHzQjpyr72S1kY5dRg
k2oC+hrMKZ6R+peTFI9BQEPWVTJA9DvGSlKWrhRstr1Dtym05kWc+Y2f8Gjb9dxC
BjCgMTulBGK/T+wiNIZueadtKyuAxjNa6ay46q3N/brSJVENm1HSN+CTh0notel1
/DLQsQSVCtgPvTXrLnbx8oQ8HhoBS5SBCBuGh0k5VgytBAS2lUu1OjYrGom13TRK
iJ/Z4U5SanztvotfI/JhlcAuspY0etY/dMiWvDIdxtvHyOLqp/kYHuWnWzwEHJFt
PUM3MfaM01+yftEdOGbu/1zSEf0OttOtN+9s2JeSWeX+HJ1J5q1YNkM2KSRAv11x
i4muCi+iWJu7RYZs5ZsLQ5mQ7m4ofzIY9GfDge6nInDWM2LDA0Bd7zWchLDbrQwl
qPiLXvEKtsVMT2byu/5/FqlVrL8HGOk0p7JPZrsepGVLGRR8Ber2euQCfqbzopu/
SV055rgR5S957YGB0uW0EOm9F/+DxOoQCL6HEQkwl4o91XoWWdTKhLekPpkSZhQD
x/+3+th7TWchWJtbdfp0dQ37qBmm3Od05QaWeNPMVTaoXf0v9u5chvr3JpH+760F
pMcq4z6tKOgNoznsze/44f81KjyqJto9OsP38iCpWFZOiy3JSPiAeTFuW4OkGjyy
AEQGEcfC8tsBEI+jBRigGZItsWjfZPLVtgDdfvCGwyW1Lvr4jAiA9CEwRTNKgGfw
1pshpQylSerb26fzW1qrcKddlSEBC3YPGHgfQIPc0E0ge3ogGucCRegqMdleE4IP
xn1LlPvDbjxt7EEJ4uUkIV/bjH92f6gKbIM+2g+AFPXeH40I9YmzmQGeUdp8pKqK
i1QDUH6KMzgr4nIDZFmR1KiknB0eTXSsj11n25P3EYp/36zAxj+f6L+f3lIFbO8Q
Mrk9YIpB7O2/yV0oOxpdsu47s8tPv0MwULzLs02mQocRQ7BiSsjx1tfqs5yVe9PR
FpWw/oWkNU2CPht50bcpqJZTob04wTH2/W4bSQKOUV0MGJ7xxLqNGQKmpxOOQjzv
qi8aQq2Rwm4ljqCy0STCRNNugJHszC7wjzqm5zx7gxUxPwRvMzl9VXtj2dz1pEyd
/N/krNWWiki02GONkjrTHBSPY45qUz94nxF2NSeSLJyAqC+ib0Zeaz97WzvviMtU
2buvnB6L5EBN1tubIjkwaeLiaLcmVDZ4Z5Zsls/UveB3IOVtMbIrh+768nd39OQq
biwqRjslX0XFJT2m/+xn8r/glQwjoylvNtBem/s384KzJ9LLqr6IZCqQguUWcejQ
s4J36OfHyPBVC64v9n90YQE+WTy48g8vQ5KXZ7BkLS5kQSWm7siNYEnye5pKhDZf
WJeGe1SIkGERCtVywCcs80ZDVfT1aetmFw7jzFCTU/yp0lGmMQbCf7eyQhb/2F2z
bvYwkuTZ7tGrR1q5rNW0JSmXqwlnfnCV7LcCZ5kAqvuRz5AyW/XqSuQKriOI5cLD
WrM24802fAfi5uVUNRukP7R4zFTeR0yz9dXHusi4Yu3x/lry1QYIgiKYAqtF4Gfm
pkz2f/6iAGWYucSbDzdPpUg9gRzacCQnPbBBlveA3qGoVAQ1UIg5DWnH7NY24Umw
kDCwfRaMt5I0h2dN4oj9Og8Nv+fYiHp4sQ+EuaQ4RDBZs6fi1RyDix8tspOLFiA4
gOFrIGghXlgrNHqkuchdY4W77Z4txeS73d/CP6lM1DHfFEsUVK23lnxEMTKbekt5
Q75r201AZPaenAeJZ5GQpu2frcJwOMkfZphuO2mDcYD8a25I6gMw5vPLHs8xMm8y
l7WSxbf49w9XvTAMYnIORxMBUOGfl64+qNfOR48PimWaaMVxCHsCZAoxJTclhyIW
7HQqkZFRm5/K9UaRGeAnDfXdTWRhHXfiZxTy7ZnaRcmnEekE7Jmd4jJMlP9z5t5w
jO7IkINMh5vEJkV5EBrp8G8TmkEiK/nFVvmN6FPrbEf8vN5fU4BKmZWFNnJ9A0al
+pZqjISbuzAmfMDuLRcI1VfUE6oyjkLQQadgDX1DifwKAOSOXJNa0+eIvNYA2VEz
Hd15KF5VN9rbwD4j0a1NLq595f0QIEl857jIRyInZPH8H9r3fDQnKIsCDX3CB84+
KQ2oLCzRU2BOvmBXhbVtqAB4dSzPur9yrKAPxhlNlX/H8vq69/iaAj8pnveoYFZ9
rNAmMWiLV8AkOVFbgPZD4L4viN5rWye0mL8xRy474vs94hu7nmzhad2AXCrYaOY4
2Er4P8hX7k+XKZqfVXvlbRsgkB84J2RUMlMnPUBWMFSfVpfkOM9JmKifUhhfeEZB
X0q+wczD3ibOEFQaKpmOLB54GOvoFxWaqzrlLjZzJbHUgupEgUAenquXtjnjGYZk
Rxkt3qsTJHNV1jSFYli2BP8Y+ASv2fKqCAYCntoNnSailQDPnGI60gWkapvOywxj
xldg1yjm71S+7c0bEVeYEQaUahHob4ZnGDV0VQ2ANfj9Uj+mzNd72DX6bJ362SFq
Nzvc32oGF4Cc6ck4dshQHz0srk27Tv6AkcbMDtH3IAF0CbxOuJiEdez3HI3NlpUo
wFigzU2v6P7JK8nhYD1Jw+6VPhpADmO29+ImHVe2sQxhWc9op9//XNmkXAmOZHGu
Wi5oh5t0EAONLC0R6iR1BOAN0tAl3cw76fFPsryus/Fj5IomeGtKkXb5Ga5ROZFp
+GPK1xV+0bUdRie7gKq5r+f1SB+mFnl9v1/2uD0fbCJgJ6KP/87o6kLghU3r7fB+
dHJVPPBEIpvN03EasVzHgJUxBW8I5165L1Y8odURtzUhLrF4fD8RrX8U6bt9DbJH
iYMccG8XCUNAOkcX8gZvA2jDGCizH1lUlEsaVwiabQ5JAH39hcoo2hjRzJ7Vqv6H
AhO1F+5nILyMn1n6GDbcmUIHVMcz4aXTBja8Z26RWCy59wBkSSdv4VxVk41HAQa/
2L2nr4rpHHuw9WIAGXG2PjTheOHUknyRlylnYi6yKgv9ROt+jfjgMGdbISwmvCWN
2MVC4EqMyhV/NlsEO0WVva0PwiEsLjfipQuQwAFMG9hKpPfVHLrXM0EBfpc4UrG0
kHyddjzMmJ8R0qjyvYxLnuBBKNOCQ+7O1JQJ+6bQqBqU5AarQkOsTTBWtp1kV1Bz
2Ba1i61LwwSGNQ67PqtVqF72DXRLCbeJVdVPvYn64lWonldaLOE4FDeJdWRXs97W
mmiBJuJUjuxFbq32+fF+B7CBwTGKfuvfDIKz1JpeK/FMMxMmrGKi8L45jrp0Y+ZY
mkRC5bhREDUgknni24g9XrykDa1EtG/e9Qf+lsVs/ldrZ4XTNzYJDmrdoqcSZX1C
PVgKzFIRBB9DuEVmttv5siWJ3MUsGfVYY5qDU95/TfOwe70LJ03629ZnwykP+p8I
rXvxue6VxXliHZ6xWECBiVdyz5tyZLsJOi95CjOiJX+qwId//IIXvg1pRnXR+R4y
rF33/mMyyPWw+dCU+jXdvk/jtHuOreNTD8y1+zNcLDxqVAVmBSywyE9DdBanablf
BZ/krng/yH5F0TZrrs/b3sBZQBJGizuPl4Fg4CYfx6X1UaUOwjiIUyDqxW9XUHuU
g5gmO4w/pOiS5dnDws61x+/zJCWsyXjxhNuOpJavv96pfeKvvzypEAxOpArlPHGI
Uuns6kTCdOC3TYtUeK3NHMB/IwL0hqEEwEr37hK1RI6i0A6IM1SOMadjY+aizYQA
L1Ip8JOB8OQ+KABj2nmSA2cPPjNJJ+gRPpoz7djcr6Q/Bv+1/esGQ4OZ7o38a61I
JZ94zA7xmANg48cm6XAggsPcJuH2JfhSkMddlCv67DNCQ38eklkF6Rf7Sc14nfVV
/lNjkdnFeKGozaAh2KHY3pZVkNcRZ3lD8WIYdXDM+5UwDjV+8nVsCNYFl4NDjSKC
1eLKeplNvgyxlGXPo5/TAPtE5MPxwiElZx0AlBq0FxczGVfcp+i2BxLTzMUCECX7
4NiSqk+sBR6r/dX20oY9gT+/faWYdFwDX5gFaSNdU4cYUFkXXAel5LwPVp0yJMWU
H8B/A26nfS8P4RjJdSlDB78a5tFNPXQhNSznf1tQdAmU6nWPwoMG/SgEbVbn9Smg
slX0mGgA16SxrCsj8pQDAlHrrNBRvCbN+ISKI4vT1ButU1m8shfX4wZAs/2qhCWj
T9mxuopyygmtMKeaCKyoIC2P5iiiviDT6qJyYGqQsYSrELTVU05HcyAbk9z56Zax
BVI8n1hefte3Y1vdj+VypWk543HEXJ9MvWhdRih5cDdf3mOSeIISV0tW4/wwha0p
gVS/dog4D+85X2vqtlGQJePxIxV772qrfC552ILL8WsoZR6ByjO9uuv9J99e8hEf
10mgkBw3/UtlomkzDA4AvmlgYgxr4RmBOybPmW0RiDBPgoh0DFx+GzC+lucYljRh
ezbK+lsUz2iPGoldA0IxoN3dzCaPqdyuAiN2ruOv+VQWqxRQE9pF9FqTmlRlxN/L
Id0mkT6srZIEbS5PU5lxLjxAXNPbBl35RxeZTyU089GtXKJGoLV9uhzzYnD+sZa5
UoDxR0jwLH/7bMPhvZ6YxPfPdfyV7+qzRcq7WvZi1qz29UvDqblbEQ6SqUaknGS1
m4irzH5IYTUArQ9GfuN0RJHT3rA4/nJRQz6cCSXxhnf3I7ZdrGZcQevw+Iw85+kg
OXhlcuC74oDUYlXvlYJAxcBoskXXuZVFdIkjNKLwN+5UxZUMv5rCMSFbXGk3I8aq
8gyyf5gAMG4xGYnEYS5A4dqArTj4piW2+EBmPW2cwo9GdG+Vsdq9N0cTz3edS6FO
b5CyleZWEjJy/eMHncPnjpmb98LBRaYB9rFvRyh5RBdLgsOZHNTkzkJJ/FmYNAFJ
/inRtLxoBbhQDy4xWoFX/f+A+863SKIHEDrbcJNedwjcVGO4iVjb0zcgvkNGHO7W
bFsfJBMF2n9Bti/W7HbxwyaDgAi0QPZIJfJdRbNuIIq35zgjirWsqwP350NvUQVf
G8sN0iJcf2vMTa5YR1E+PLnXUEN0aNDnIv+jOBfAM6T/RX/CF7nKjXpSd3uV+IgS
dam8kIr0zqZzrmUQDmsEJfsTDzP677sejW+JDrvnG4qLCEUN1zXwudaWgXLWfFes
La5qTZAUDIgvKUkXzAcw2SuzzyObs9NZTEyKohEav5ApVKuQwSZbfrih9DXr+lBc
UGfzTu8iFeKRi2YUFn8er2x3nLR/f/w8ziB04I0kA6dxRjvO57E617JDW2VA70G0
sVH/V6AWKgsarmXOgP+VErUwGUbzOXvpxzq65rn8qR84nzt+vVfL6TBN3LMSz5Tv
0LziKzdYuwLAWQ5CF0YiDtO3kcfd1HWJug80gZaJXfwlDu8q0twm4CizUoHUTiSY
VP0pmrYtdQeHXiSf4fSadgk3OocYDakvWUOQqdZBvFF76cBcDxKmc4+RETeeCAOj
eYFFyC4Wx4Qub7W++coo6vblTfXFOGHS19x3KIBmKllo8vt8muIJMvwawE+HlDzl
Ww/iMUIT/UM82q67z+bvibSMIbiyGMqKMd8dP8UBj0Ngk4ZsYt9kvNb6f+V1jG4R
ISW4ypXfEduc+nDABVtJgsgjp3ENQAk3P6yoU/SBt3+3JmriyOd0UtLoda6wvVd/
OCYA6T0zLBDXiGD2CZmEVyD7Xf9A48Gy1m2HAKTC+XDpGl50sTAZ0sWXD+fChDv8
Tm1LAVxWd5zC4zpnh2s4fD3YYqus27RyFOMnXIf8NowopArNhHqEyN8Wr+ZCRwLO
+J6n+fxWX08n3zD0RGORztCQf6E/56IMj7NtLT0FoNCJ2mYGsBAOJxgIbzqTL2ZR
TzsxXaj5IEx1zKiIaN8J80qIG3+snrHSBSXG10nLsnc3wU9cgvNoTdXMnae+aWb+
OvNntKREOnwUSbi5/OngKWEaAnYGX8jTxXoxMamvGWFGugCtaDHWLn0HGMpiz8Ii
wUNhy4XW13Qll++WsWA2tf+ubcDc1cWzjh/OS7fgCDfnrMDjy490HY5S7lQ8LEkp
nfV9V1PWj1uczp9wNFrR6hO8Ct+Le4ioGIs+GVWgYrfjQ3suIy4m7TZyfzWztW8U
LB6tyc4BdwGaNiHAwl4hZ3hqGCfR8/BNPGYIBgfQnsH6eFhFP8rQOxXKLhVIUv/o
VdAdr8M98G//yrtcO2oPxSzvKdouLAoj0obd9XPKhXp9Yum/1osJ83Xh+zqjh/C7
HU0seQ/iVW/327xNXpaabY4TPagKJMAG4fa6Spvsqf/aUO6N9Eoz+aFATmK8idq7
qglRcX7ukmtTf7LIa4xSxMTtg2Ekm8VcEx1r0QdVNXY5Hv1ACTrestzpmGwBJM2k
8aMzl6GKiDpdgpkSa4h/mU1DhSGFVPVBRlhuvddTzIqr3UTi/C6xqg2CZtf3yI36
Rl/VrGKesZXrt9ng0SXf8XawgcLzL/7d1T1ww21v13eNejKt1bi0d3He3ZvhUG75
YKRligiFEkCUENJmIPlW4Yb0eM6tMn71ENZcINLgl0Hi3PLOZkOAJuNTbdRTqabO
lV2GB5xbHJ0i6/TVKyZHcVZuZchSVyqF0YtxpCmgGcE4zcAA8GjvqeAywcR9Za35
6Y/q8natw6xhg2tKh34Jr55JJT15XVGLlxPY6A+ACZuhQdsgJJ29cQi/ne1SNcW3
hrWk+XaIoHVcDe/IC5OHDYY3/lAjRFUPehWGwoD4lAdPLAxCjmlf47b61Td6gKmj
DFHWKuZ3P1P12kGjZ+3SdHdsnINffzNw1pCXzdw4MYISAgJyPUr4Lz3v7MsrANda
BsMJt4ceNF7xil9hqlhoIIMBWSumdxQy9KcXDTB568I/4+Gb/TvkOc1NOtDDSWQz
gsiWULiWvBhbWyQaTuct7UsDqjjGGoJ2X5n0QJvh/S64XHUm+1Jw0LYZv0sJmACP
UYYwEcNp8PF2G5LznH2zt6dwb02y1gZZQBwE//N0ETl8S4YGf2mHR7qP54ESWdJD
rMk/a7wtPw8iDQDIKQp7eIfws6xfV//Uk7tv69G0uScPlWJsvUjYCk2TIl2geIZ9
6IHifJaSMvvRabY/gjzpaKhQxVklxYMADRzPTnUi2fboarNPGHis0Th57C0qbhGi
Qf2zIMChhmLBICb3fvR/tRqWQvJtZDWsXeOTmWTAnYR2dKdffzBglTGi/XYSS1Gd
cS1W2SxXCqwtsNPZkgifaquLsViY8oow7veSf8aolx2/pC8AxumKNUpEoZTXmP8B
HKwO1/sir4Ig6Cejx7Unc8WIIH0juXQLb467N0t3YjsGEDwRHZBiuVY9L6WLEwQB
D4dUJpD/uZ/e7NO/dlKGB/bhxF/5Gzpa8ZEMQJRMGYfzlzDEuqeC7pLLFGdTnjTk
F1C8YQk8mJ2SdaUDSLA6UpnW2rkCSQvqfMyZ3pWV26oQv7eREeiyiRX//mmwBO+T
uE9HOxR9OXHSbayPps4BYjGzSk7xXnhvVipsfXWyshxVJDoKYqp8n01Sn2+LB8bz
IWDVRpKhEkZ4cm2tMo61istyRSN2URigXARR85uyVHob1XSLQcr4Iloq4dRDvyon
qzeGCE7eJpqlOM8lyIteQDeXwk0knjjfoorIp0DSzZliaTBBTmqSYKg2X+ChxbmK
0+O/KnT/z7Qj6bCyWvXTcbCYN1wRGUR5s99OzLyONaDVk/rXW2JD+1DsrSr/VvIG
0uYuDA40ngl+kjxRa8ks7gfedlgS+CAu7vweEmo5LZL9fgdQ+zYvqekBaZlXYd8L
PNgwVs/iDt8Yqt1jZlpK1427gIC7BJVtWXEe3PnQMU4uq3Zw4vb48KtMCz8MJ3uB
JaMNHfuj684QlS9p7bh932rskU05790OoQd0rhw/zNUQN1HFO9SWij/FfeypEemG
BRAPN/AW/BO5r2S2LTTqhs6dh/eFA/K+thR2jbGJrrqNn/BxdwhCuOOwsQLfUt6g
NF6yEUU/I6/hLVu60r+2Y8pCKLbMCSeFxbrT58j4G57IJiLfyyLzh52dU97a9Jd6
Z+fMUF8rdH+/pYoCySQs/yrmbNtjqH2SLRJNaAcqjsC/osuUOlbedUDnGuFMbM2V
B6N3HxgvQRNoWRbfn4va5sUaLAIjvnuxZAa76oDQje5ISiijsu1Gh5uIAZ7onIva
t0wINnVA86seVJxKkJ/xRgVtenYd2Z5KG5xxmbynwgG1E0kGOqqGkvamkM1PE6oP
5iEm2GVKqKAUcx5YuHFA+MOHUptvShv5iTtbchQJd6Ie99ZjgvVqdksXO/V/fP7w
0EMpAGtvQ2CScYc8ywhlMV7t7y0p4QUEbXZn7nAR/Z0fLekCc3kEm1yj5kKpLq6r
73i+ga2u/yk7XD/6sCBHWMU9UePZiTrpPdl2GqlphubNVtxwUyKXdMM+K0n0L3Ek
m3DsC4gtvCIVzICROaslmXhpq/gG1lk58KT+BGzqG7yOhKDBJh7jgXKIXN++++VV
KF+4HlTfglCtbbAPUjwxxQr4+YVFuxW+cvLUP3Uago7KOdbUNtCvsN+ypKWJlsr8
oFTwzS9537sQa9DASmN96mJ3y5I+BUiowd17aV0RZbWiovxfEhp/5Ew3noTJ24D3
JChaDUEk3NZVfPy5gyb9PCqVIqz7Qat2++WKeRdU8ZlX2qIOPfjWSXfCuKVIt4Ve
tiZIjC4pt5Re/q4jKfnLouy8u9m1SR5YD2fXYrNNrYpYHNowBY1kyXkshxR1z4n3
pzD+OJ1FBaLNXz2Xjr+bzoVFEe/KptZtam3BaOZ1dlORgslxPhQR8oJ0lhL0sqSc
HDG4RJbcPkSerqcpS4jyZtWEeAVfjUkBowQFCFVcS5w+3Q+gHnWsTdZY+J/XVbO0
Wexx2+HT2XbW4DQ/BElgkduTlRAJM99pSapDYJ+hfCQbfTHxOtJrg/yAvEergsr8
wlM8Xnd9zjzj0ugfvO/wc9ZqboZ+vzCUkHrUbbADssQvGvr/8qVdf6C7tiyIVa7D
4GPHvqm3D916MCGNwRu8Ca5HNL/Rp8xwUeXEWr+6kd0U3xgOee01R6KwWp02j8V6
SMH5HQ8ioTcBBTPjqINgEhNiXjUbgFJIJhhLEuZw68X+Cx6z+aPRaOHdBEOuY7wV
ms+phCVh3KmJyteEgQYn4/0y+rXa/gjGZXTNN2IJnANX4sZH5QYV7SkT0NjEKVqC
o+sTU1YLOZEcWEd8Wr7S14/iX2/xdEfsBlXuVDsnzs2AS6j4xcIT4wq/BGyZCSyZ
yEKVncLNzT9YYSKciTRt8rax/CuuTvchUVhsGFgjZIVP+hKbthCttcRJrKINb/Rq
4NUQop/zPavYMX05RXpsfM1nU6RSTE6kQICT2JdtSTw1hremeovrxXyjVYlVmek9
Xyyu91iQO/Z3TKG0qk043ZmjEwBFL3+O0unzfeds6AwWy2L25kp8RTEmYOHOw9qz
yGTeK7mvQQowuL/NRXyvTKNqAd/KinqGC7e3pnfFqpqJ98/njn6xBE6OUHdq0R1I
wwcPUF8g8TdChASXFxgGJbLK1nddGHNdnXwTWcpdVLmwJ30CN7YVLMiuy0X2ln01
IGuq+7zqbDFMxXFz/FolMifQu0L+/JXoujwnWNxTZSmV+Jg83XF5nGVA5jHaPs4l
7LXbM63AYDRKRGkH92TwtbdKFjyVhNWv4T2vuMkgzdViAjMBMqE/EhW8Pfuyrhqd
EaWCAh183/YIvunpD5NBLyCUbrMtx6rg8AJqkoEGbZUIoiVeY67UDyykcqL2F3Pg
2W4gjyOFzXyIWmbatmgf7EE39wgP1rBnqkHK9x6bvgkOKc0fhQoKdb97rxQ5eWKQ
Xup6mVYn65t/fcNc/JT5wCM82qzJbio9b7IgHf+Jxc3ILi4me/iNDxzy2waKuSRt
XSiU1JLmlpEFwfYE9to1p0Tq/J0XXMZs+d+7AbbS41HRmXm0DZopZVRfd7TtTZZN
zi43S0PlghNVGu4gswudvqVt36UyMJ7TOyT+njVHsLh43SVMxqrgjmC8l0l/AdMz
sbd9W5uoStkjdIbZu0VJYtAW6YOQKg8VPdysKsZfN3zELHZUS/tdcst7fPqkeLVQ
Jpveuz1x0vdNM8Oe56mNifue5QwJCQmsf1rr1nyXDohRcpCNMFufd3XepuOZqEcM
f7hJduT2eLfdC2LTAa4pyDqfblZMVnkgKL5j2i+yTOyn5km22+QH3tuDFTyx2uTU
LHi/PRigLfX/2tzJM2M/xGDXFTBjd5/wyJwRRV4oPSsKUkN4KjWOvfDocuvvM7Qu
PayuV3yk6TtNCSbn2upHcNeV8qh3Q/2sllNoNYe7pDLxlZqlVBlfs8P3+UxtGTWg
ER/y7lBVWQJCwbiwdTNN1Ea1T5lJbe3tb+m1I4jp37b9b47Z5bQy7IwZ3Dsc00Y3
EIYbBZbHfS9koSecuzEJSDhzGhcDE1EMX58DJiy3c6qns+20FqhtRMzVnk+KygiA
fitElhcIfKbnUyyzckNR0LX85e3E6Y7FBKdjhFYd5XiwDRLa0L9U4YNP4vriaMkj
u8Sop1QwN/mR/edrXR7aUCnzSkI7PpYUSkn+qCAbRxKlbHdFYXwY/bTKKS7x8Bdw
BYAOqxarvsuH/8lsca6RRo+xp5Fh3eQ6pN6jNaUnrZazNqZul4EqAuKvwxpmWEry
6DYcxwyW2tTsgxN8GYqiSdsjgGayvDJVaJxYab7MlFb31m+l0vzmS8ctTsPU/9Qj
DvjWJzHB0Ca5+ZjHQQsR7MZ/BsjqC07Iq08j4zMYek2sMmYjf4SOStsqPa4NxGJj
Prk4MJsyUyZbssJKTCedA+LGxXkul5QgcRXuENg0yA7S32CmD9YUhMUiWgCzvzMo
voIzDkstBDSIoMnUc0/WLHffTkFUyZvEXqRyHNm8aVGGDQUH2g4aRNjGCVWWDiNx
zJVgNCaqnDk2y6QaRIbeVESW5UL1Uzsi9HhYWBA9E+LxON3uaNih0Yx9+StOMUCk
2tHKVvkvzzagXKny1FO8rnFNiBn/leM9dovadv6Afai+vd34CTUNkdUo5owHEWqL
p4mDQQQyIfpLikYmYgYXu/qEnAfoZ4IRxdByiTHHXIM8S0cRTBdVNuxWpXZFNLrG
ANxXP30s0py9PhTzEpungiVVEHUxorLrAd2MGOwfA5AmEeJvyEgri4fH/1vsV0mB
8qH+0JIPrtnR369SD01/S1GN9Jy8tIZlGAwTf5f9fOgILqC7C76uGYMuWW4PfWDN
cN0jXR5IGuAipciVYhIKHNwISAHIckiL1XFypb2adENPGUeYmj54WSUHPVBXIu4r
3mrmAKSoZ3R7n/JU3nMl/EqK05SVpinKdG7UCJqATxI14RJhBtwJ3kMeVNvlfDyu
DUU2YkZOy80qx3AEX53uzoNBld+PR06OwLKT6i3w/HH7k39a4DUkmu8f7RR+zF9K
zISEMpXU6ui0e6TghT9c77aIiHOuvFv/h204nlFkbP0daEGNGsqhvUELXVAKSnYG
7Uq55E8odE1clRPGDwHh5SR5RuYSkd3gbGwulT3jBrt7AqL5slN6JmYUZ+XprkjS
il4fwoDOeI66qXb5Mq58FL5SY+obOO+nU5hsifvg+OG7F6nRSwZUgYMEtax6mwHD
kDZ8bmCO/5vMjLooRMTK788r4QCgE2S4572+pG+UnCXuv71BVQWC+OLV9dGn2566
6SH2VetUTmRbagdr1hzqQ/H/7u4lKXCOUh9c/Nghu7FxCnWGqd/N47ZYWKoQG2HL
IhTGuHEwIfAE4+g6vGRRiYxqjK53/uiOMzXpFd6nht3ZUTLwvn3qBGhKapT+gpaM
mdN2stZ4w1Bl2QHSDwD8nup/Pf6EKISXgDVkJy7ltQCD9NA+fGk4UzICWGCmWxzl
HkrP8RqP9SHkoRdbBo8ydp1hTe4fA6qzEVTL9A2V1QxhSVZ7eqxi4WYJWoGTZI3P
+fuynux8c2QH159rPDCvgCrCJgcQRBd9+fQ64Rod8I5BwS9BIQQ6OrNNQOCHtROH
lk2UxjJlbd8vc401SKvgfwKB6rV2A2pIiYAEJz7Axv+DDMAkGqF9qtjg+Xt3E7dZ
LHk6WCXGXQO3AtUhQ6keRlW4C5K3H2HAXoGGEmqRbWQv7gHnVfjQ9ILEb3Glqo7E
a0fBFAHYUSqDBHOm6H8DM5vhekgCobLXpvD4lK8kXV28d/nXwpbILjVJl5EXIzYb
8E9rPIZNl/6OHQFWe864jOM+dxL7PCWbZGiIy4JWoXkY8nPJPP+ycHCnq38BDtGM
FZ0jqfMKVfTo5ESvvGuf0F8nLpOAxpTrHzZg6xGjjOb8YQ6k0yIpAm5JrKt0XWK/
Y+AmMk0hWnG2NwJQqBvXTXg34Ym8YhdMZFKtjNMVgY0c0ncWqhFy9JBYGyvrBQ0x
g+ksBKM3Evo7FUPWkYS6DN7mqvO0ExgzHqUQFMrnWZ+A2B3yCnSU56fKYq0GOCy9
QngSp+kvOZe406R2U5vc2A8bf9qMHXS+TsDs2/+4zOH0lCe4nef5KBeBKC8WqwIB
3hYMk7lrJb1Gx9QnXDkDgYvo9e4oT40oec7dJNld/4q0nVBGuc8uwg3GICk2TkQ+
RtbfkgC/Yi0HUsK72mg2cQ4MgPd55tq3WKs8eaxLIEfWdRlipfsy7a4o7E2yXCBu
In4Q8VgFOf8anAxLXglf8iqLCqswXh45cPdiybIhBBHUzbvGnZVGJzVmS/Fc2icA
S8dY+uUMdBXnWyXVHiDcq9EFqspilvifhsCTp4c2uZ8u4dcz97vwfcRprksjwxor
nNUMeX+YXqicZASRlQY3BVbKfgHsUvmO9cdTAUVLYOWU2qHtC3T4zS/eN8fdtRes
tqoFFvwOZJCsSbvIHNcV8Mv0o4cvb8PBMZgJWbLCKEc923J0hIa3uAvhXfjZrA6q
hYJdqE4EhW2qcbHh4TnJEznk7jAMvl+aAJyWUloCt6mpX/PXDjxDiNqYIgS4FftT
4Z+0Ah0hnC8fQiH60Nf0m3eLF+mq2k/20UqDP2l07Lse8hBrfqrYV4yZOyfDnUob
C+t2oe0Z7rCdx83qgZydl9nTxcjw5CndmJDzorQkcjWTj0/PxKrTyOUoaBIDg2Yk
okMD2Zi2yLr8PGx3D/mKUmLUpGzHvIw1v0kT/nNmT+CIcOxiARqdr2dP4l+6glsw
kX+paIKl7GZCECMWLvUU6t290cVXHuFVmv7X3YnWFU0jyZa94UZEgBYOx/Gcl6JI
zdoFqFEzavrzysvn3g22+exGw5bi1KF14RnVHy0Uw74ljovzbDZ6CTkGMF0qHboY
pFuixuV9TMJCkhEYc1z5li5tEPZ1m4uytpap3RKQPsPlLPN1MyckFzvI3fzb1x3F
/s3PwX99GpZihow/XE/JzqyVdr1K4aHZkpa/rU4bhwoZwI/ckTBQfGfLLY1g2IQy
2Gha72RYhJWFEtIEd3pv0yobXUUEbQ2q13YfSpCSH/pmtEQHbHOE7cbd108cNG4F
rNELwH7RCSw6xV1gCHcIvxIG3X0nWdpZWk0gyRt2x9nveD6GZX1bw0/xI8OWRw/j
gIybF/Sq1S550UW+tz4zrI6VrBRlKnyc72f7gXrvFyeWBTJt/Ef0pKFWmkLsKKmU
KmV9QaiRyoCK0A2feTU2nYYQfFDxjKyv6yE3RJSR/hswB5MBkEZYjKLaUFSELZYi
a+Tjzkat2uTLxaFV6JJkl8BRxAk9wtpdmIDh3b+FL8s/0TEOeTYsP4f6u/9NtAIt
iDatYIlxFXjCS5BFaS8xwApsJha1GlD43g0EK/b1+gxm0/S1plPUW/tTRVcJlI8t
16NV62mDqqxnHs8zoQyi9W8lcu5bDYwxjfhTtNiwwd+7qDHIcSjZT8tZLN1M4llr
CHrPkTuq+qdI6OhpDM5mujhnKZBj7WaJgscTZtg78YYr+jgRmTQFm/3Eqj7ScBV9
rgJgNvFe+zmOffB5ymy9gu/nkWaPrSYT4ApscOh28KdPwRfs3dm0j1WT7ZsS5fYc
itBVZ7DfnoF4ZkJjKAzwtsfn9AHMr8QsnKlsiPGSj1g9HcrUMKCiWmhlH0YxQR9v
WZvc1ZYwxyLYsRz0NWrOpbBlI0ngdj2j7SrUutFALh5eI+HAGpUQQA0KU0j7pOLL
UbcwjnEbGCFZsAMHE25S1yss++M6ZRs3DFC+I2ECAj50pstZPVjCPy8lxcstHm7t
/MggL3zqslHBHvxx9XETOjj/zWBLiAR11nsBRG78NcLPDQYLM+U4AKjei/LbXWM5
BjscUzAJ0bic18mOiIZjJuSF6n4EnAbArVJRhK6ilhBxhUbIwSE0g7NIZVH2Jdo9
lN/BByIBW993XtHQuDVor4AnLhj8HA73RNHIDFZSelhUK7ONER/Itb/Z7l/7Gqxa
xqVi8kLukBDSf5Phx6I5VuFS623NWcLZFcf2ImuH2qH3Wnv5hPhdArlvZsJPQPJJ
FU6hmEmOkt/++nnVVtDm+j4FFNr4k9CLeiq+KmNnuIL7ycjKaog2i5tKZTgHiv5e
xL9PTBpZfu3TV6Q6Tfi5mSw8FseCNezWuwkG0aeo7lt9c4jbg5CTtNQ+fHE8ejEa
O7/zZiQLZ6gX5OJBG4dMTNEI4cBd9YZkWz60KVjiZxDY1lK+/XKmfVzBxJdtotBx
Xo9B+wxlyzFD1CP0T2nczfHZjF067VHJhaivtdmKX5ovh7RXd4CNcfTkzg30/H9O
Yuwz3MJrgNNGY/HWSsMxC8Z6InJSzBRkMilsx3BzQaURNf4TrNHWu6icrQMIFyzI
bKj9JZ67QtgDKBbeZr+5PNyKNHc+KaM00E/niYR8F/Y+igBG6kkmtvFQ/zpygO5p
+jy77CjDXdrvdFCl7iOS0tk+MiDpaCBo55CJEdYeGvo/bVlN3IE5uBhdx0yfWt8c
fqEqJv3fN8AjiDKO66u4KRP6PgwYBaw9Enxl5d6YAWkHPudHAfEu4BZI4BvJ21i0
FgHAAwMLc82rPhLEZpHEbxcRfhJxJmZ+R/VeNC76ijZ74RoQjNpAkJ3GBs/yGUpm
Ol8qnQweKg+3nKaScotIhyQMPCcmEs7vFqnC8ooJ5teV8n8TcOpA3dd7xfiOyvmr
0p9g3SxgJcQfkFyVatnoUlEqh2GwWPloNKY7S7sn4NO8jJC1NTu0IE/j4qpg1+J7
pHv7VvF+FbypK235DW/zokA5FSrFEopTvynoh0EV7Q9LzGUWsM9+YCBFhADjo5sN
ILpmFkMsk3Qfi/fQtQpNSlYMQmDUFX7Npn+O9yerZcOsMaKGRGLzdljzDc3h4ExB
5ooOmdVHtX+vqzxqEz7P2d3k9t464+nUDTM1KH1cZVQpjc4jBQiv+SV/pJrL42fV
TijqMvmL9TT697TJIvjflNHicwVFraKt2INzsJP474hMr1c0bVwHoOmedSp6W+b4
j6fgQBniRrw9K7miHlsArfZ91E/BwtjxGhXG3UhO9Mjyn1jEjr0r5wambWPzbyYZ
aM/PqrcJRy40TIqax4VhtcbzxZZBaciqwWpW7qs2UTm1E0SrgYxiWUjFZz3UXLyY
JqMtybQVxMNCF3sR/FWkveg61V2YnuVtQjUfBhXMBWkK/ko+A/F8MJp+IczAvzxA
Rzxk8SZBMNVUTII/xipblrl6u2RrxSe9LYYVjUr/HQCeek2Lg61yRA2JgYep/xyG
lf9cnpfV3AwvcwZZmFk00BsYKxgO68mZaRijxN8UY6sF6TvS1Ehv0Vf3bWGQXZAP
mfYbCF5y2JdSBblVh4rMhPRKfppGvWMWYBo5SdbsbFFceN9ifK+g+p/uTkJylCxP
smUgtNIs2VP7RzGJdxcoUXirXywZ5rbTLRI5xXSgId4CBhJ8aycS3iLeGhOdl9xU
jM336tedLXu3oDF1QmP3ea4jQda5xpBo+rd1WdZw++/7F80AQeUc7o9mBzn6df5z
fXzZL0q0PHeFU0wDYYB9niAYditHqhdfuxaZn0SGUBhzbYew0/dZVO8fKcE0HR2K
IcUbblezTEcTh5nGojW8LyIy/EUpcl56C25ZJQWCqfOBOkU6p4fqJeKr/Q6ewq57
NjnJoO+PLsfyOnE057t304g5G7sRBUozWq2BHN+j9cejpVhics7CVy7SgeUnANN0
SniAwoO5v09S9zBKSp0YBAPk0mM7OP/2tdsaTS+DJ9QJIcDRdS3XLJ+IXCSkMjvm
jieZy6AR/1uEbz+Vp110fXXiLaGt+zIwCEQcC2gq/wJ29LzuqkVVpaDrLOGukVK1
Pj3LdPou+OZr37MJD/+QGBY17NzeE7kkk2UM0xEwXpnrDHRKg6Dqsq/pMVSZRlxm
uARbjUNg2ipprZZwmiMQHzboPBL4w1Ej3ExKGO86tqW4WMUmDesTzkF3uKhH2Uze
OZd4v6cT65wql4Fgz1GkMGk4y27G+6ih/A+0eHMElW89hdRuDKtBcHnVmgHtLD41
kx9Nws0mmr6B8nfYg5eB2SyqMjjcIclikBygTuw4yjoZHryitNCGS3YG/E6Oljx/
44jfV9At8gfw1ow9hsq/ADX9FJfZOG1j1Zdnf7OX+Oky2TbnJ52HKGuV66OlqO5x
SLSgwpe1xEEKAh1uYc++1V1riLLfAEWTwi6kBuEq0cb95y0x5yKceOYBfVwAJnYM
pj/fqLAh4eKgEnR9AV5kwkGmo7wXp2jmt79F+qLueUfC/7wPbfvobc2Fn5RKto7z
jqpu2tdUZsIRWYsIMEc9lzCoMJ6dU1j2BkIvcG0v0gHePAX1N3EeE/22dVp22F7k
DRQwIqcGuE0H1gT1AcAfBYTlzzpGy94E7/2d/azpOUTwDiK55aBy8pjGyYOgO682
r0U5KCFwLfDU0ygOoqkgnjrL3fRtAygeZEhFlojcSGtSrk0Rxm2TLEr59cTHjrNE
oVYXtoYx5wLKiU7kCUmfbLofnqSata64KimKHLcc7hYWYmAY9FbRsa6kJXWIZMJ3
zA1jtzRU9zXkBHf+2gOCKmDKFtg2uCEjL67g+o7nb2uJKO4k1fzObre3UGSClY3x
vOpn90+mEZN5XXrskA88oFxv8ucZtSWBASnb1ghd45NDdsOAryaJaMQ9LawaeoXK
DciXin48a+9XvnpbcnrMCVLfVlzXO4gWIlsLFzZs0DbjYOK2OuxBmaY1SRoVbxJh
MegeaON/dGLKJI28EheYux+xSKQtL7ByS1m877LNuICepoWrB5xK0/VFYCVtewYu
GrlcNadkrn2ae/mIAIuiWvm8aTa2WK3IOal+/inPY/42zc25LYWRlwlI1RYRgdHa
SUzrXaODIpMqYES4TZ5AFfEgliDrovqQwpym4ztYMgxH5wRCzEvwHeQl2tcs51qy
4pHdDtmlOccrhOq+aI+p9RtA3zy8MIMFT56W3lUgJEJ9/4NfpDSBqrJgGrtPLYHH
mX+ep564+ttnX+Ms/M4OTrvXcvL/mmQAamVgJzIaVONcpWUJteoNm8jbiVH6KOfk
lvwihs2HQtrLP79QhGBK3nqataXk3L4pPc3QtSdeLUKlaa3f954ohLLQWql/mltu
+ArUDhFXRtCywsXMKslzpPSA7jeuo+IK4KZYoFceik92IRlwkDK6UtPubIvc3Z+A
WDRycbpthMQYy127p6cPCukzW7urwnKj4cOwrr8qeLOgSe8DFhVoTdp6yySzLAfG
DCv3hMPwI6wtyH1lFhxLFFrfMMGXPHxRmyEyXbQR4k0psMPUAeL5ZCoq8pwt5tGo
OLG6I7Oi/H3QYFXWEgMVfBGD+A1fL8MKCnUDfBUXcTjx1Jve1t4LXKCwzW3D/NbL
1AIFpf9u8Q4dE/ojmy7ZM1e8NKQvq1CpG+bxJp04hB6g6eRW8Eh21BbrCb3vBUqj
HzUnZeARY8//sPqY6JLrMHQTS/203kvU+HAzW9ExnEy6bjeFdap3zuonO24tWYZX
1yiv8xVOtHSxieqhHPyRlp8hiS4BnxsbMMMOBbOc+AciX+LJWyCtghFAF5EQZHDv
RUEl6kAeYqxGiu6UOV+f4pvY7WXESK1y/yJr+OlARGge57fDw0oddKZ/q6OXUNpV
BEV40ErKf5ZUpSaAWJ9Ey9jl/5YZKeju8nYY+WstzLvWiQ2ZYMWlYllRua2a60pA
4Vto5buIdKICK+khRBTz00JrLfamOoozXxdkyPttTwZmyTIQgf2+etmrLl1rh/QS
aAEydw5MW7yZ5IJlQnDs4uL2KX7YSIrw79YgDVNojXHS6LL1XpzBVwSPbROpUtm7
2g0Ct9nuuSVRX/XWj4os/C+R2nQl5k3EgfzcFnbkql6BBRCmHW5gJ12QUa7LjqEN
e1c24lZWYHtvDMTuM+tQ28vSlcbPID4uQsOHeeOC5HCGc/MdmNEJSx6LNpO2KjYc
6lfKMo5TveJGmBup8Mvkrt8uhCa1L/piVhoAJi9kNP19g8XBmZhkfHc4qnkXLJUf
eBYpU5OdzOQFnSlnAVOFAQR6W+FmaKxMWnwrifYvb4ZHhkiqr8q4h8pKAf28oMNd
HLcFV7Y0PjBD7P47QwbOZI05e0Q63Oi39cV/U1y2Ab9yUND98cWayd9M1maRrMpq
jJxGQiBTO1C6iRm8jhamueD228LZVZZxTksLQlTwc3UDmmTivOEHw5pPN2pyOHWh
kpnyKfML3INmJosMOXVmi8A121eCiF3LwGCKgHja/rq31zrrjcV7XUvfLlYSgwVo
uE1GUeTW7VPyaxOOaeRWv11rAEMa6srB7TRZZQGTY9wwoqofNBNP4DD3DWXQxWzS
ge/jJ4pmN39EGAeOssDc4Jwgdc340sWVeI0ZXGXSXYWoDdsqno5p9aL/Ao3/wV5o
c7fHLi45RcOZMELxb9qKpxLa425FXDDsWAGpc1IawKlPbIA94Are46hpsK1G5LCL
tNm1GmfqmoCfAl3bJTqkSG5bvdprid+6jQKqF/jlRSnhIoUTJUTqGNPukNlG1ZtV
yyV9UCqs2akup28bxSlIKhkaTrm3iXDMC9Yy3X5knGlaC1dUNZM+1xfC/0r1DFfS
a5C8daIpWis8GfXuCknUPldpiKkSFbnZ+D9NxDZNQXoKheDu3jRW/hjMVB2Vmy94
rgaMUKI6zCd47iEXq9wLr487oMFqK3TLFPwL8JZ5H8a3gX7jLj4xFwoNdzNL7ndQ
LqFEO73bX8kXe4ol8AH9ODwsGtKuB7jRoXNGMLoaZtZ66HoMGHMjGMAx90KIycvh
yde8wlBGuvnF3lQRMvmYZeR9L93ZniHzcjbO+uSEuSNlveF9feNRnh4esua8JaWA
qESo7T1/FSIhF/j0eGw7Q/pqvoa1puLI7ik2RHRVkP3yjtQWWA7zO0eA5S5BNaP7
2L+VZz0HFbVNik0yVOxBuso7EkSMTkHMZoZUEaPu+WKsgVzvlRsF9BEczXQUBJPA
7qurJT9yrMIoOxPXNPHN6ukpnuvO/SQvfVafXlyJe0h+oqc570YwSyxRosOmjjLj
xFsbGDGXOJ6HtA0Yi6ZzqYq7cacZIcHxX6eN0YJichCAPvbQIfFDrRN3K26a5dLB
G6yA/C+bLjQ8a/a7pO2haaQwHe1YhPLOecav2jDwgaPlFGvG3XATiffCDn7voe0U
8jVpqaN57/6dlcK1LT1WJFAMnvSQ7LohPRhgOs3uW7d6xj+kDfhdhFwhtQ7U00hz
DR03fl/ThwncMGcgb76P3O5E/ALRRNKwg9XOWn75GCRM/Hujlg9zy+h08YdDB0nU
8tODt68z9I5yVsQ0No4SnndfN5O6giZfqwCbWjKmfXM7uacNloqQnlf2r4301W2E
gs9zuh+G76ETp/trBEKBoL60Y1LtD8yIccGg8KlQ1d7bZ0sOWW6TcoYvSNFct/W1
FCcZR62fgkJNDbtuMCCZTbweN7n/b/HeOFmLyt760mqtWWEN/BqccRPl4QppECqT
u47fmHpnDWQOrgE0rY4o7pwU+pjJzVjpJVBw96L7hd2QDH8bGGfudBzApXCnnmlR
cpwjFichZLCIIS+xw4O9S1tsldnzrNcpYIcVmgwXnNx40dnLdSIpqqbu1u7XqOfU
qNl9s6TAbjjLGZbzrcrj411QnEBLHHyYYD894bBCsYmM68v1VGX9f0SH8xFWTYRi
aU7F86iFBIPOps24HX8KqlwF46QN7Dc/oKAY473RJaTT/o+t7I7MzUCNzhC84r3v
XV7Wow4H2lsZUO75XSqBJTqrWHWKzfxOGw+QlFocn5jVePPiWA1pPFLJ0JVY1gGS
kYYPg201zaFYgfBpnuRKFZKRVT1xHMsVoJw42KZW4fUcJkb2aZ7h23B8KTLUzPIU
PgKEHlCHfGu0Q7MtzIMeDZzN0s/gaAQAwfUzJNijdq1ZubBc7cxOMO3y5RYZxxwh
OniU2DbdgrdjMspnV4/EDgysm5zjGr1XaRFfReiSOBPlz0dM20qN3gc8sbkiDgoH
BQxIcKaU9GzX5AjJPhIShX4ZDKl0dURbNnCBEv9qJjERLFy+b1lH51W2GVCIU3eO
A0Fx9DkyMFU+ZH9bfnSviP5BKUGBX/GnTZkuJRHCD6bLJ2N/9+mwSmZ4699JC1gB
wumXGODgqciYMd9hI/IXM8Pec4UHsQVyFZpKJMZQYbBwH76CyXx9dcwUSMWckrGq
kMlnD0Z1b6tAt7M7/mLs3l4wkhcf/txNH2uoXTw8VIdaSXD0046hAk4kpl9ILqH1
g0lIOawi65gmDhZ3dQGGl/p3YbC4IdqniPRyS5IUN+LUMuYy7YRkqfdgeE46WhoW
Oi+lqhJfPrHtpJeB1L4WmP52pk0tvlHS0nn1SBFSabtKUnt9eXKhlyl8XIwQL0GX
F4SEA2JP6VxDIwA6cT9e/HlxG1W7+xQxj6r4jJ9Awfdw7k4/VjswaNwonKKAv27s
x5zGG03SdM/ZzfceHCnPHgNf8d3t5oF7bXCtaKy1oFyvMzOa+9CYg5uilso6YDwy
JKm1uu+SkyROMr3e3GoYawAVtNt7x7KyfGC0C+QwDc/I9PtaNqo7Sokeqlo94AUN
l5T0ej7yTQtAG/YRm8AH+rNwKKO/Mx194ElTpeMhYtcDRzwO9PEBEz5JX7a3/YLO
QZl6NW/TVv8pMS/CcLMCVhSl1HWWR7MHJndxueQ6D3GngElNiFJ7YhFa1QqMVZvQ
O0HUOfp8gLJdjYfZHH0tNa62dB3Q5oMBQgYyqZq0Wumvl8PQT7tJdtq5IWygSEYG
+zr/+xXqAE4J6peWI1LXr21Z03js/mce8zd407TCTmZcDl7TJECu0gF2wHx9lNBd
aRnJhEZmgO99iHa2x+omEbWerYnI/1jC33qh9oef7Dz3HW/RVMZAFOdCJa26gtTC
PucHdLdSe7w+HA5D9aQtA9fKAvRKfw7BRw0D5qLha96nifQ7A+aIzbS+nqiFegm9
+limTVIeTFOKmtMcUnleRgmdEY/wbcK34slLWn3dtwfmwN2a3SJG7mMG10kQsNp1
0YaayWG3v+v4PiXM5VcwXDyMYtphz5hsN4q9JNWiGqedyo707T95gUdI+UXFdyd1
4Y4Nau8Am4r/ZHGP55Fn0Wb0oeUwP9gQOPl+wvD14UzNSGnKlAXlF+SV7hvJFO3C
Ve71smb7d/ss81HI7vMiRFAtkktxdgY5rYDJPpC5szNXmU2EiM6BdOwhDJeBKcFy
2WH97YLeK1T79unbuKHuJSNOJ7BUlXjLJ8gADcmCfg5pjMYOb5p9xwQWw6YFfpI8
eYm7jp2sLh2K1oSby3wsPRtHOHlP6+eMmPpSX1gIW7anX4Q3prBtHBvyYgVzicR6
Xt1PhRx1/64kaehM66wejywiVO+hJyyW64OOXm0EZENW50PpbURCiexVeox+Dlg2
vwWQkOcOddFEbKDYdpCmSWATWPDpQ2Mf+I+6xZlUVmUtIT3gX11E+xX51VxvlSq4
ZiuBlq60KWNWYCMff62c60fCdBSyUgA+2vu2N9ADV5nfLrbDVW4aFHkaij9WQIjU
vHA1lPBk5286kC7KOr1kzXt3KCcm/dsCULUAJXF3gmCDgEINYNC8KBVUXrdIXVXO
k9z90cFznYaC0B48z0eeZz0JCkxOCi7kOgF8PKGBmkSw4ZL35SegtH24vENzYHW1
/yqcBYnbjOQUoDGH9raQixi0NyUXRNVPzgYq0v22ACl4to6snuOPzG1l2m/gD3jK
rsUXlLGiI2cdsF3u1bA0tQosnAakun0B+tlCL0i0BiJccoep5SKnNsFEgdcEB/aQ
ufZENPrBsrjs1jkTEszi2d1NiMMbz4Ch+zBSw+VeDhIyw4g5T8Hl13afvVKsn6sN
mTLyg/AzK4ZjyS2iE1ZjbZ2AKgVETwyXW0B+iysKsDXj5QkLv0edBZSZRBKQq1eD
z4wm8Us0/4UnXhFofixCZd5lLd7YOqdZpFayPunWGdFX+sVQCD5wvX8NDtwcn8iK
lNQQt/O1al64EPjP10nZnxCahki93I+tLEDFbmIA5DCV7KNqEsNhshjjqbkvRYjZ
ML9sf10xjF0RZ74oXewV5FNPEY+u2DkOCbYkdxDNrw1cssZn+jisqXK0kz/f7ier
XEoRxWjg+mxKRDJATYJ/gvVJoj7sZDXiws0YVBL8SfqVN3c89ac3QSkL9I+eRtzN
U8gozfW4RIMSrI90B2IoowN9KXYzjITI6TZF0p9G5muqc1Eph6lbq3e6nqF64lvM
IFxXTIQKD7lzEMh6fH8cLQoj7feR1cbLNh4CShtQ9E23LV0XOv5reseMHRsjtirx
xmubaZ2tgp5MlsDVgRNQ0nRBmQJfguTJUtpkiUr9HXydiopWt7gPGxmhUPeiPqkO
KF3T2h3aky88KxS++xVSKtp8mfy6Fu4DweyW80Z5I7/dKHD7c7wUzhSOIeMgn/d1
d0kUZvIEkz0ofqoVliElMDef/uKcCj+78bxBq5N/RX8eh5hwO59V4xoh3e9GxRAy
dP9hAKeS07jUKOwfBeIF52KEBx/3RL+vGOEDGisGtqPVu33CGNoCWdSlws5NKs2Z
EfdNNra2HN5o4Lyt2zHldziBzekUR6Kct2hJvRSCL6mAdaDgb63pP0cqrezDEWDv
0Mfh48iWgbyqi7D3tHcJIA+2qV58v7tvvH4FIaJ5Zkds/XdNbsAMiERxVLgz0PeG
bgueWKni3jGU9cWdsMF8l0t8d3mQ5NI961P+/dQNr5CkSxcDWQGKlqgwlW+Kkf2K
moBsgqes8jfurlYqV4ywj51r0pwCecV4aPDB6my9/2yELRLOq0I9rptiVSGBrP90
NMcrAg1jgJyNsczEgPpNocwmmSkO75DTmUbNMoJ1QvuIs7SZACbqKIvZfDPnJ7av
0QhoOT/Vaft3pbHqZoOmK/2zuG8DbsBf1/EAk0xvYADtpuCMIsCHWhk31ZN6tGTP
NJrLoW9kJYu2I8sT0qgMNe8YNMjm6zzsAk1fs12931NrXfB/IsXwSITYGv9qoXE/
KNTGPFYqKQQYQMI5jf9i722nLRfjNIWPDtyyXCrR38JDMqvvcuXE5pPByzrhsD10
7a+R7ZuiGbh9HF+Z0J6zxNui87jDiCzeGIT8/WdkRcbsWA5BzBrBn75VFJlBiE9D
7VyDi9Bu1QyH8SjusBhIN5tZL47NWQa09hJGsfPSKMbrl1DAInidB6/YPu0yEVx9
iuBn3N1H2I7I0xAmNXzc95iILdRS851fXuEDTrbdxZX172u/n9wRFddFZcpVP6Ay
vbE+7lhBqJLjk5PL0+/MtMJRLUWbFcoplfQg0q6sNrfr9yxeRftY+KBc6LU99GBi
Kltu+0A7Pmv+2zOwazUpJRD2se7So7AJF6APH66d0cUjErCXNAthdwaEwpSmeWX2
2Vp9Hvd/mZezGhvd33nbfMkHHkwSPnZQxJeHRmKHX0QNnChLTnR0ah2SGHW9Ibc7
WAz5F1oKBr3ASj5nZ68MtRMxaL0bKLNZQB3/lWgPemP1KjW8zzYeY/5Bh6vMSJuk
Vmm7V7sdHLJmvpip/iRWp/QAI2z+dNzmKGhxySQ063xQODRKsAmDm6Mxw4Ev7wBp
rcG6v3q+DQ9kTiiBL1wYebNXEpRoMlE+f+Y1XUKgFwoub9sRJTR4bPhi2R48aipP
HFs8Nvqow0QOKoAXdRzwkcjCYGC57vjbVSTGd3MXk9jvlHrwC2eF8EMQ41qif5ic
gtUig8W6T4Tbdy5ytz7FGKYJQQx1Y2MchX8TEvLriFxWsOpceoDIU73z8speA6m5
HZiR6VuKKsqEbz70J3lWkSKFIyTbx3LEXi0AGsJsBkKKaf329Gq9eX0z9U68hVEX
H33D+Smg0sKn4oQL6a8P9Ok4OosHUZJHB58hwEa0GbDe6uC10Tx7iB/Kv4vatYsa
rH4pCSGjhZGw9ZdYxZC7BwtHQYM/kDVm0wfNnnkQDBJx29xopKcVc1Oh98bpnLyq
/UiSuMxpKOtBNbbqgsC2TAl7qv1jZ2B6SkUsT9PfUQFb+6KhoTp6io3EqIytNIoj
qljycABiwqnWnZqRSwjHhETxM7MQrl17v1QMcFn+f/CHTv1sMxG7mh8XHRs6+G9F
395RvNaEwGFRL3bVcE5GRk28GqBWnpYPwSo/Tvm76B0rL7t1aEmQfLaOvuDhU9d4
61tN3Y34wdnDjG3+g7zAPnChfwcTwHzn+dv/2sO5u4qfb0jXnwDIZpQD3EDU/ZmA
m03vYNMzwFFp+Qxhrr30hOLJrrhpB+2wDcPotKVr2GSqntg8aUgy4Y7TPtRmkuz8
WinPIhmSB3kEFTA9VeexmNllcBGZWv/zcF+uriZBPsCoTy1Uy1ZNv84ogbWxaqCm
djSfpXSBnV/K9Het2QlwBqgZzuWoJfoxJCRwheOU2GBiwQcTjTEDS/CLvhnvTDxh
g+0jz4Wsnj/+yuhgmQD6Kbz/Yl4XL+dsv96ut/WYAyWYH1NnadKNoo3exqRTceRI
YZ0w6Alc3ImLSnTadothZZOL0Jju+JuYNxbYAxJvFqkTmGDz0EHqa65ZAJdtcQ71
YMChN/zRS1tNF9VG5p7vLYssDUgAgD3isiLyvKlBbxhBdxoMkPUgxruEmVBvpJAW
ILLunGeq9cnQmL+FxXE9LVgkRi1FbfhhUU8tJrhTpOa6cbdqEvbzQY4ggSAuUpUB
xTa5DmyrisYOAp7XHo6jrBpWKgR60zF9VDewnOUwk/lpCggkcTfUHECf/N2A/7JR
UBTJEEMdIh/yBGg3I73xb3Z9D5qtE+kAc5eM31SMe5FLoDO8IZPg4P62VgPhSHaa
HjCgQvIXe4nhjsJWd8rolBxVvKMRCylEgu9vTkCq4+UZW83/512FzayGLSbxa/xQ
eDGYVHrtutCZwq7RoiEZz9HIg1ZUzBmNaKbEqp6h9EQIEw0qeiq3srN0mZkgXo5b
g0RlZ7PYnE+r980n2bDqoSugSCWs+c0Gkf9ut4Lb5Bl43lgEZmg5dOGXjqnDd27r
SgAac+J2CO1Gbt60kfGGuMaU+vp0QtQjHFxZeea+aJYDTnaYg5gutcdnIXyp3iX7
Li9HBL706whiqXTUpG5PtIyuOnxHduDre5KFNXlhlApGcMhFjy0tMuRMcln7aTq8
orVTeju/7IbQTmRODcH8sdbaiFqbxxoNMP5JBRkyVAeA61Oy5APGuI+CD3M3wTKM
1CTFSB5f7/yz7Q3C7Ycp+590zocXA+GTvF08X66Jrkulp+9YBmAEaVMJ2hpY0LHl
0YiAwBSAW9NRFyckvaQbDsIdYexovthU5AoUTKm6jCve6ZMP3uHM/i7MxWkglMVA
o4AwGe6jTHt8ZLNOzZBnd0UaG5h8g4xaOXj/1gXIHPmL7w0TBUYnkcZiaStNnd1c
NjPQ/qlfAcbyElX/EgUia62L1E3uI9stRYL/IHjpAke0PmuI89q7Xf+sFLRNhn7o
IJkUMO80NEZB5Yb+C7UiuUMkVDVy0QHTRE/sgih0kphoiRhablThn9k5LZJggDSD
y/BJyQDI+2N2hrUiqGWKkIBIYpiZI4OffkrYS48ghx0edeGmBCXXkLlWj4RlLQIi
rDsWIQjMInQZW/gpEEupQPbNupr3pnIKQsZMvI674yeEBAmBcYREQQd9B2YQaiEX
8rau7xUdCTpX/u8wtGl5G68rkvxXGtL5yasApqAp/wwk1c42hr5jSyNLpRU984bm
HapTmLjBEys+swfNWspAPFOPGxDiGzFETq0967V474GcdwSJY2XZWvACzrTwxe4e
j0rIXPgHTO/nw2w2r5f1IKQwcL7yj6gJnZrIKD79LFrVY2xLOJus/+arZO7wPAU8
Pd0TszC65jsqtLT4DSp4TP0NYRTWuaPC04V1w/v0PKfwxDhJtoG7rrvQIMjLc+eZ
DqqR1c236DDIfSfITlVTIKT8/MJbccvPgTPC/KosQQkpPw/xBjRLhPcXsEPBrl6J
ywP4bYd+Sn/spGbDIucMrj+boEQ9nzEHGvx6qeTFCwzbAVRjfSF15dKwkuU7mMlv
DzNiKYasYALTb0+IOXonPzko6M4JMz9VlLoupeMu3r6P/YCxplOq5fK7WQ8bQheg
9xblnrLMOHdix8o6BntvQYm4Nk3k1Z7IUz5S4FwxJxCH0ycCYwTfFZXpuvAjvL3a
qOyCpdfaipCkGWgH7+94FreW4yqs5m/M0fTCl8Z1iiEN+n4gNtRsN8ctXml09l2j
nxDSsdO8DfkT99/36iOUnU6OlxvwG4Bbsp3dzVV+4dcH3vxBkxm+27MygmEsvTth
XrTSG0sAP0v3+o2Z5F/VRLvNcEuTewjq9SsFCQoQvDeut7+/0qCnkkpmBylhzw8G
q7ne04bdyf8DkjVAP0KOkmkH2CojBDSI+I3nXRxbWq7KwXKPjyHm/+c7ZgNhYf4V
s6oI5uA3RTnZ4UKyG7iInWKjeQNAYry+GFBElhoeSZZJYEBsvWCfMqyTng7jnvFo
PM+hhfAPzl1AXAXqbg4YOcsy4+KyH5od0RAfFR6rSWm+v8VcP4l7iAJC/ZZqJZCq
zsQsbnc5AKyp8y8xO9Q9MFHM89YJ6b92SMYLBfrbpegu3J0qda47+5f1UjwvttKr
z64zCFHRHtHPDaXTuLKqg/I/Dp8B4cxk4Jf79OQUNIjGDeTlFPHg5HB+doT/rb9C
V1X5JaisjHjAstdI+Opo1PPssfwyJAcO9mo7ebIsasJmH7u/Fv0QLoISpDk5mqJM
74mIV8i0oNkiBs1rWEAz9ZB344BYNerOGzPCGvtfWduEA6Y1osjccod+zn9l8XWd
nAIXyJ2ABrAFb+BGY6aHRHoCiyEFIUS4ttpBnGtWHSXhFvJioDpScH8NPflwWGb8
IigY/zCmEK5r8KSEZSJXcwbrEHEKtYCufLrpqf/guhOrnH2xV1rOBuq/A+fyg1Yh
uC2x1P/fm498t4nvFt9YZkImrWiKp4TBaVygYdD/PW2VAwCqvWmkoW9Izcfb30iv
FPPKKIrM8Kwk+u1lNNut+NGdMbh/kYXAGRyTt29ld7QyvX8nUYzdVVtDJy00FeYU
4wjxQXrS1qMNUn8zBuuUcFc/FzCQ79qSb3S2flmWXov7JNlZriJs2oLmxa0nzAgJ
DRiennHLVE1PPxIukkRtgEoxjd1TOxIfi8zTCJTL7zs503uptlR96GLxMjsQSO5E
FL2f+aafuTxK94yOG0gLhSE7/Vip4MQdXiJXH3TaNRKi0K7nxw9sKxBsjVc4+lU9
vlve2Ngz+Q5xPay3InIADOzT7K3fHpmYf/aZLL778lqrtNX4bBuTKB0bjdhZYt0b
BLHu+8ZpQSrKzlG5M2iI+pMUnIbJUdK7KMopvXG9PbVDttosz80YzY6KCV+Casng
Mq/a5+8Ke9rVRuAYXs5tiu8exibBDx6B6bIEDyJqEth3eCnBxcRbokW2EIzWdb68
HwKC3ZVQlIyMIo3nnqZIK0ndHqMgruKy1P5zX6OgwKCFQxtSpaG4Gwcz43ySbvgP
b9rSKGJcpMDyRUCKSZJpC292q1YsUOki2zliddBo4FzYlkncskewFWILXgBJwtwP
rZi75NOIVASaelIvjJ87Zq+EXjxW+ewmi/Mp7eSPMuC9c7jQnoiNRVSekkaa3t2Z
Vj9Ytgse2b5U4O9tp17eaKyFAu2MKRoNI3tccBL/UCG0K4K8V7bVZhHbt/+JIeJY
9aOef3iBr9YxMH0rkFBoUnBvDDSZSaRJsws+/DaFhaGz4kn0LT4GjxE184DOiasn
hdrj1YY2T5UavT3Jj/vw9LABfIkbPY0SnZHPrkoraxUYpihSFjwj+hCm1TfHfZxY
vu56DsxMrnT12obiCI7nuR90g/L78mJVg4Izan/Njiy5Qrzp045lZ5CVQoI5nwsY
sW2wFRp7Gsy77EBd3AsVVlwl8SauDq8sABw5sJw+nj3B66iUcldEPgx0Y6PZN+Nn
iLHKVrxPbxCh09CCn2E7PkATTS4P7fY5AWpDhlkNZ/44pp6CmEuNqfyxcof5oIQs
9StDpS7umwOGE2IOTtfiL8kYdwfIi2Qv2SS8Mzful3KHrXjUwSeqCoj3PqA2yRK5
pLPREMF9l0UMcRb7TxVnz0r4JTghX4U1GxtOS0HiBNoY07B60Zk6viIrpReH759u
drl96rI/+eNMf/t+i/4WJeklu1D2w1LRZqq00ogBPjx/mbvVkg+XUHGL/9xAizqt
/saq173JoOt3d4mPMCBYIK2+T75YwB5muOAn3EnUul93lo3cWi4wvD0Sd9Yt+HOr
AoD4TFXVtSGw32KD1GhVA4fERZ/rgNvYzhz3f7gJ2Htom6EvfFJssIaOvBHZRZmY
u8JTH1LJ796MXNkwzklDaI43qE58+yb3AIhiVOAXc3C7xDzjiim2qnOD1urfO4ZS
URJxgSv0lGCFSbV/JWxfLGnw0QJQlZShELOZuvBdZZhyWVdeBlXvxV9Ph8A8yYKi
id1LvoCkUXSsk4Rbsf8/+BAE2t+g8XvLJ965vJ9NQmvUln5dcJt4XEBBMWjxiMuc
F4hMPTT37iJ9ZpXDamI+AfqEIM9rM3XpPWSv2rh+tLaOD0Xd7cAnNlAq8aPlq0l5
riYuxAdm96Q2o0Dm+ojZ27XCCvCl46DWi4nQVFsO+OsSDhQeBbf4VBhYdHvZJcOF
zRW+vlrFouhJxoDpUBCyw/ELHoepAOcbvmvejIauiUeAqzkgY5KqaTaKDDwlkeSB
I3H/a+6SxHExs6GQBWKmlqg4MNGEGUhIvZn2FZC7VsH1KtTW0tpLT8EnjxY+ezak
DdXjnhaTBQyDdo5ygCW7coL5pg+X8qEiuw/LQjn7UjczHz73Dut4BPp9UoKyP0jf
MfZCJYWS3Pfyzop7/ETslZslZ0pyHogNIv3RQ1KaDnO6a8kqlTrRzyNXBhhCIRIk
WbTnpuUAb+wO5DSSrG62j7+MtArhNpCYGTYYVRIUb1R3U1q7xIxZNR32Eu0hgIQX
PkujLj0AIQds9czjX7P3E3j2Mgm7Kizh1MHGfSvHlEzS14RKhsO0bZ6YyxHIjZ3M
A2XLq56tirr50ow5eWiQY93Lvqnh20djidTv2byOQTZazev+9bC/wArzj7YijUhb
mJRS09tcVxz4xEcnPGj+7WpZDT4lAxLEK/mkJLeouNPITSALqEMWUbPOg/JlNIPz
FP8SLsZNTP+mnaIjwr/k2PeOksZC2im57Cf5gZsyDFRjgXDyfG83lE/DAWkmtwxV
CgmG7DjYq7rJs0S74eQ1S6PW+V3SB2v2Whg8C90dkY2YgPQksJuTUCszbAizvpU6
xHqioofYaHd/JV5hqoRmjCuZvJgJ9vzh4WQVqNdxcrOqIsZZwcs4+N1sVJRs6pM5
Phu66Ryj41VGporwk8ItUaCRXSMVZhsNiH+tyBm8v9Q/dLjAIe8x9Vbtptzmeaje
gd2lLyiZkJsfKqMF+lACaydh+8P4wKuFtRvZdEDmQiLA94oII8Dd2EP2tNYZUvCE
zxqO1+4lxL1BAMbhlwn/koOEytaGCcDW92wdzAc+PyYPyJEhtPvBUvPuVwIaCWDx
H5u7CdqVQj/RImA5ruoal9vqDnYcAUvUsbM6uSp4TiHWNFUbknaotZLICprTxOpa
n82h5YVsv8V73bOV+avL/HEQIeWk31ETnasE9mWcv4VYb8jKlOZSW+2iGjUm3KPy
1kE+PJM5afVyK4YJ1/7A76UdKZBFxSNhrTXKZXgfzVSAohuJSqzkVQdjmZc8NlLj
9E0SoZHqgKn9613WbGtpUz+EGhWwbworZUpBL/fJ7ijpDPohJMgIR5YzgaK6UFPy
kIpcRbsoHwR6d/YHYC3UJDdlPfE/1shTErQebyXKMRp7FHpLzO+FrAVNGTjVehUn
FWCawL7XFjBOcN5cO73lgi/IzqVMuxsfs0Tx9BQyCCzobUsh9ImauZ6xPoky2yyf
K1kusICbYtXz8weczUXGG8IsxJQS7jKpWEJNtpyY9XbJjG4toXpLeH+EE8gQzTrp
TQvJLuPjfbZTpwI1RbCVeZPOWCXESG/XfqdSEEoFcdcOzRC7szHuFh/zOqMX8Xi2
i9Im488oGNrtTtT6h5cpIDaV29YYvCHuQtOuHo26UiveGW5lBnNypqOi98/Yo3p2
T1SaaLIYvx1dJk4RPDGSf49OGs+bEFmaGfMCknpImp9ySjEI8vJeafHB1BJQZb8t
f82mlC++aiURzxll/1WPSvOrpeA79G91V1G5x/weCdb3O5Q0Vi4gD4hZiV4Wrgom
JMaiCWaXWqUm8kQDljseXn4JssMhXcD19Iqvh7/VcqmBo44l8vr4BK+1jts2d8og
DVGL1h3mT1h4jCOOBFh5EHOTb7dZnoain5jVIfKV4drfbj8WKPfC7+MLD2aSbj0f
NzrmibspPlgxxiL//gcft72nGr6sumo12z1tfox3dxBhoCWZWJyBkMMn9KkR2NGj
AFpltnl8CZONkLIeLwqI6SYM/hiTRTkLHMgK+Rpc6KB2QxT2kcZB/QVnrqAGO2KR
HSjH5SdtXEi11NtY+PO/Ohwmcc2z6LVzULFuwHfP2Ro8yrZ5mSxCSw3l+e4ZIaoL
/WUnXh3AlYK7n3SWZgxNo4lFISLJDEQ+qbVGFKi3XLNhHvd/Kr3wc2H9/bP717Uj
nuGOf5laFh6WapDfqRTaBeyqwGQHJh3UB2MkNiVp7ORfUPGpJLHP4j0wYbBsXCZn
DwmKjyqSAPbp/FMaANJUIBfKvvpvBM/OtAZA7vISSiD5JwDeonOUdXAqTB/QFxwI
4pF4ixpWohlrUXaNoc6hUusj9uavtOWex3rAVWf0moTBjGS4l8egcasGoHa5xBWM
ijgpNPdKqLllPhW8whJBrF5Wxe/lOeW6riMVJRDLwJtDShNOfm8pmaM1clv2vZVD
cYHY/x+YOozYORrqX0l1Hz9mJc9xtIEWCkkKYn666AZ60NzvfFy8cBVy+33eJf3C
B+dY4ncfBrcNhZrmHnGLEuNGsVufxkfT4nZhySuvVRRXDAvkh/RRcsfeZdoQe/bh
RYJdejHItquUR0xYb4lcmk9rELsydLN036FIs3sXXF6EGzI9exHz9/vbcTQNpsUW
hh477I78Ca+ElDHcoAujQFAK/X9PzsIHCH0v5ncaQGkwYHKYPiB7pO4V41x8Xfv2
BIYTMnyXUsG7Msspgy7q7D7GiisNtI7Gs2xxzs+W4zl5wd8A2UwxtWNl8f8aAuQN
HCuxas+Bgk3wlWWtatTq8fKhKJIFUJu8zWtvjfixUvgb3LhhpMorL3XvlO9+CWc3
DySk5GG31eYj92dRSYSt0FRqgYuuDeHH2Ui9hK1aJy8O/OACmmjgy3CQ2lEVPwZh
cXE9DP8trZS4br9TY2InmvU9k5EUB1MDN+oZApygGBbbShymMHE57v/JTiLuHIas
St7GAMCFmK7CDs4k27TRjM665DoUcBUvpnXdYFgd3t+mttLMapi87Vh7HtP+87Ux
05WkmhgiP3bfVv/ua6ZE3BSdoN/zUN8aKL6potKqPs6HYewkTA17paV//xyUFdne
vD5usr2wpdITqzcgtiBwdHsx4H/eccIhS59zk3Q+a1cNEjA7V/5cGLGIby+qN4vY
eDOR99CTN358S5lr1JKuApPjHpgQGE2S/YI+UY7squ19DbCudxZNzW+dUfklUDM6
zinGTXXrE9zMN2SvHsPQeqh0iVC19GZG0J9xo30phVLiAOXp+/nxutNPyg/UUs5T
gKveC+7IUVWBrp/WzrNgqM9Z7VG6yckiBGRBiMgqmhNsv5hzBV8aeLIAa7SSL7nn
aBrOSElBAejsVaLN6BYwN9x0frZkaAz3Uxq3shLVYolZe44+B8uGSw9W+ZXLBLwM
Pt7iairvN7aZSbakCHAX1ycJmAswpBfrbRC7QmFRLl04w46Y3x5wXyoV7ITE9tCL
lbLoTSRAYSYbnJVc/Z5YmRB50Rl5P+2P5dfCpvsGgq+bTgYmY7gt3grwktSPlPff
QHN3My6MSARNHkrmlsqOn3ouFNv81RVwtiKpbNpoGj6rXD8aZbu/COQmRmv6D23u
OeBTLoVLjmwMM1H365LR8xUkGF94sVZIopqTLmCyTfvCdFP0Mp8f9NzLlsQ0OpVV
pdZZbtfomKJLScBEFnhejSP8t2HyvZKbG9ZF01YnM9s15FTJ6IOOA3AQEYAUYOMg
dgk1CktWCR0rgrmub240SifXpVBZPlbHS+GeAzqi9dweunLw16CoNI6Mogk/Q83f
mVIV7zhS9DMC/ZffgTyMr46QT2cJBcLHaea2WDEAUTc/mX9joGPkKgFzzoaJjxBz
AH/xvGQuB781T7Vl5x7unc5YjbNO3BrEPS5efRFLD8jTCeuylN0GNa0r48j/iSQr
wJc94/r5h8fGRJ6zPG0vqYl1XziyswgB+ciz3p0RPiDfG7/AEuiUEoEVWX8AjI+H
fWw7o/NnBy8cnlTx5YXEUcNHlbF0l/FZvfpF6IO2MYsZcNuIPEU4WZ9KMmqNZPOH
CQxli7Je8btsuzWXSCmtg2X4lPH7Gp2e7EJW916B3RDstIz7x8BKIR0GqwbBXc7u
zwhHL1VOMYJj0JJttUO0H6e50WqbgR8zfUGRetXYGyQoIX1AK4a/ezv6G/Rb+Tlw
MqE01olTlk44kN9CYP4B+TftV75eGAOHSydj+34jlN3dQHgzq4YmnKrtZhc9U+JX
6sJGi9AJaZcCxW6qJTuh//W+Sn5tyHWC5UV4YTYwQcwzuwUlsOyyS7O9zFDyZVW2
jci+SlC832Y5yZZszUhoGybezmfXUkn91VbSiOVFze/sh1rPI1v7PmIpx3IMmJfv
shd6bg8nv8QW4Y5g61CPvOtbFoXZrk7Kbxk/SfUsTnVtF0cvVEyiMTUxZTjFr449
mSnlONbte00S1HrclkCWgMnOhLnyLt+rGGlxXesp7OwRTT3MzGobCP2OAvhY7ELU
obCV3P3dJbL/e7bhKV8KpZHWmUDZXadeyLAVWXSWZcbhNafQ2QLs3QIEH8q1zk21
V8Xn3yCflI7gAwk8OKD4FuoYiQSQa7kTrIiOZenLmf0zwdAd5gCeBjwjxRWza3t9
clMIQ05N8+yIBN0VSiJVfBdrJKF/Kl1p/1BRMOP9bO3uft/7X8CFF4MUSLQm5GNR
aStSuj3Qx3/FCl1dbv0ZnAfR25N3MVjQviaBAsRZomDH2+JxzyIlR1hkDOBvIcip
NOAo2fgmLd4cOH2gyxvNpIX8QcmuDTr/rkTiYOx6f6tVbYSxW4RzNXf4DsvQIdPX
RK5SGzIXFvBI2jnb+yGSP+ew5SBi2vkxReyQ38iJFtRmZEXbaTwU3IhmHGpshSBC
WUwK5TrTFoGfxSSOAGdUJAIQJUk3ZtvZtE9RAdndSID9PtFTMJFgUBHy+PbhX+gG
+GrmPTiQjb418rQ2mk0+bYV07gW4hohXzKEp1Ng+kVtkb0zlIIIHtyBqw6P+tSc9
8Ka43X/+9kD7HjwNRk3hauAcDuvcWOh783kMFc0S0WsJbUB8vm1+HRL5j1GwDYxr
VIKCYNbCVecRGIEVcXDqx90xrIOLXlM95cs9weiP6heOkqWAc21ko3ni/uwYSWdt
Nny+YbBNDSj8tkP9TtN2lbB4OhxKH+AfaObQueYW4qg8kZm+UxtXmDd3iPFCs7+1
oIgDG3CJsDqBbfyVQJy9u/c426edB72FuaBlukkqmZ8+7LGTQc9YGV9dcwNI7Wcd
zMYkH/eDXzDbl6SfiY/znqzABn5dO4Qz23nJSpDJdGG1Eqd6l9D4oRHMgmq/HAj+
I53dbPOxNZ9CSUASYeViODbiRp35PBN2cM57S1Oan9pX30ldiezyWGVFO/uEKOq2
GyaDHyDDqsQnTCPeKKGGAQkCcVgyMtZmu1mtmv20+VP+eBih3in4oVCPVUkeKIZZ
4ZNqgCrJbXJPZq7xoRx/xHlz+GqcDw4eXPeDjfgI7rZ46CxKvxXuAYuw5hudPcOK
3jGWd5mOdo+MN2hRsQ6zr3YFz9w8CLqK+Hbys7zY4AP7uyV9816lY98h1LAb94Wf
GMes+VbKGUdKR7kE+tte/DF0NOoZ2pggl+Jwxm7mEXVePGrrKi99L01pnVgs/f95
ZukVmKymEYuXHpXmrfASgeBqXo262fITczMhVyt50IdxdVf20mr5ZEr13sP/6+sw
p/1CjDcB3mlrL8ueacNOpTUWyRdN/D7LuOXRPfUceqafGlf3Cwzdhxh5bjEWcsh9
QqMhzMcj4n8V9n8Hxk1jCxcL7RdEqAebHb3PKsbDdO+U//TBabj6ZE6UAToQl6ER
KTJGtl5Q0qGYNbEYXWOXQxohADqHSZtNkRibH6q1H0lDLa2RSHIiy67duZmfp/Mu
IG/Jmesvh1wpp0E5TasGYCO+d02IkEJLCvlL1i++BQoZESaoqIEATRy4tgiBiBIC
44j4dTkhAQJxIDsikIxh4v1SoYKyJ1AD2ebpc+xq4i7hrmy4jJYorEy3vnmDkcWL
svPLnxBEuN4K0NNftGIB382bX/xLx37Qk8AFjnB8pbcil/D7q0ECZvKH2pKL4rv9
O3W+JG0qcip+fifwT49odRkdLpeuApxFmx1PKWbmOxKcRm84ITJ2rCYN11auPalO
oWxZ17DCyUsLPMd0qcTZLwnyA/Zw6aVKSG0F1QX9RJBgY4q6j6viagL29KLjAGJS
qFOXhpIJGRbp3Awswrtn/BgfK2VWi6+3b2KeYtP5JP0pLN4esyrV8sRknHbSi+EO
Q1qx6IZM7tZojbOfYpo7f+AeaLq8BwQUJUmT71Rxt2sHvbtvlpG+tAVlrrAJrFAH
7BF+0riPbg2/tevHrNYQrcku7aKtc37Ona+1M//ZTLSjhOkzTYqJZ5Qh0zzlRock
hHAhDmLkGJfvkdMnKrIeZalkl5BxfjrMN7S8rN8xHEmbO+hsIQYOb0J6mm9jQPs2
SrziVbUZyDpHAOvJ1MAUAQ4oomNzgJHq5oJ2QG1nyyXxznfp47CeLf2CwpBfKnPu
djj0FgGmdyrswcEStuEklI97KaiHQj3pgX2oGTLk2OWi0ocaRWFxHO5KnD5mzgcZ
k4EzxuGAiBuKPsBm15geLf+DejeCDFMrt4YVFNHG0reMNi0W6BIWOmPF+iJ79d3L
5HuyfbudrOHgq85MysjuAPefxmRKyLDpqTNKfPmwlxGcvz0GASR8UpdATymGOzw3
GrP8aWNousOIKXerEcsINxKiQqrRnAYVnKcmXi2zRNyuhDbLapFQCpWlyhPZ3Z2D
a428EQrJVhhs3R5d5h+zzA0B+bOFpXX4dT0tNCefkrk3KZ6eNoFQHbQG9yTmKHE+
R4xjr7EY6NI6rH2hr49OG2ACIS+mxLR6tLY9h0tRjNkMnSu+DG9UU8WoxxmJfLDE
XNFpy0jrtAghGMQWHjYDyrADTvQKPSaeqbd4rC2IkcI6qd4Uh7m6r5jwEzZjVczU
ETvTRWPWq0ZeJL0ygRCQMMnv34Xsi20lscdXMHrg4wgw6qP3Qy6UwSeQsWbO76qI
/lLNerIOSk8c4nFJt79kJn3cKrs99D6bK5AHb7TQM3BY6HzPZEhxyivy7ercwfs8
ujnJtXIfQ4RGySFkEwN5eGwgdBsEHlLicpvJmD8qpvcxeruziHOYiHASoeGcBk8X
rXGiGCZyZoR3X6y2kgcET8ZePqYkSQcJ8hosah2ATIe45zg47wMuIkzZqmVcwlt3
7klq9iaYqR1CJVRE31GoCv6PiYM/HrFNQi6WASqGxXo3KI0+rZSyB+VkmhqYrXih
enFn2kOtBZy8K8sihzxa3NQFSolrOkWcsSEO4gZ6VQl6wfZjv1Tsj24BP6iB/v5g
V5bmNuwZd51c+LJfqr9xjF+aBavxbOFCYG/xlaYXHHyqWQ+Gt9MlQKIgp2h/Nb16
Uydcz7C1KJgPK7xetrWRz2QbXnYgzdBCEXQKZYhr1QcHfeQniiqZWVsgyijlyw3u
hoSgxH9nHEqP3H6l31/zJRgOGMaNjlCdloY/AiNhmzPcEJs2QMoM0XK/N82f8jhL
fJ/rxEII703tw76cyhZmKBI7ZtimupnqsjBjzemIfn3vuAVG5drfNUcE0YBvEnF/
FH2sL6a24s1xC7J5rSBhVOUdqEYrE0rGB4N9eijKrVS88f/XnP1WGj2xCdh4a3Ol
mjfVedzJYbMauH8xLNP/6Tt2oNRoW77O5a5HavA9REIXRBRAMVQnNSaFySt+RxbI
5bLmxe2ptjZaMEvpeoxh4KVakkVe0Qdvo0cxyW+5p/RwdPc9adUKP+p022XBppBu
wlgdRaOtnR+Lmx4WO/PSmSZAmIeHQGn/4DR+NFJZw1vXNpllNFK0c0nJkZnenOnk
UDFAIzx8cpiifRK+8jIWIq9IPnMiUxA79OqKkVQYtHmen7jBcLqc7UPllxHcK5jz
PennRZ5Z5H37ZAMF7QmDIZ5PKUJIshVxvoh1kzZkgi8QjVmAf1ZoFpfvGp0QQZdg
9CdvJqY/wqAJwgfun6/aUBl2PddJJT2JigwNrZHDFar+PDJN7++DT9ngxPUzzJBP
Qa/lVBYIeX8Dy4fWT/CT0xFfTS3un9cIdKtv+1W3qtlF9EruBg3sMS+Ov3xCqmDi
TglSv+nne20HQe+GSDBz+UPfrgM/pXsvVDKXejUzIrYSYm8BgdBQV+hyWfEsABaD
aAZp6GTwsDC75HP5Kes/6GRuFTQGNdnSpuOdOVqITTEg5DJHeFyCBojzyZ+S4yAg
6y9Or/AH6C/KSxE0/fdbBqpxTU02B+CsNWnW3mY1vh4se+BgJZltzlMZ6lk7UozD
5CVC2FvOPkTL21D6FG4cUxhNVCruoGBPuKFJkk6khDiePdTJ5Z3Cjm37Ryau7Tgz
lok+BN7bGpRVcmcA4/Join4eDbSbQ5XgI71swJ67EYMsGdFMAuk2a8riWlsEPTeb
5WuwdrwBZbpdqXkoV2fLQIyCSO10rYPS47MIgxHFkTKGZS6wJERPvjXBOvUw1BNx
b3uWtyQzGsoShjlrHmQvh7DfmFRKlCtoW97fC/HKSUeu4N6yC4RbfA5r5tGSk2ti
hWziL29rEjLaVN3B8zpPPYigexMv874PEWn1L0RcJKP+7pGyZIpnRSw7DCBBxkyl
sjncMiHH6viU4Fj8V2xp3twU6x4UP4hbeT0gbMgYCkvNUqCMJgIW6Y8DnMGDr6JC
RZUMONyhvSiXdKBiAHMfelEeTkPk9kNvGwJVbc4Eqoghowii1Iu0FZjw2U8CoKFr
KDYtRd++owTPmgg2aG/ahJhelgGmj3wZhr5KGtzfZjdqUarHfjhHJpmq+m+pM3jZ
beYMqYeUID5TL52HgS7399MhcpGGPOuUliwg2Q4HTCy/jL6buNkUHVtkpJujHaCm
u/JUVIbeMsDo/CP/zQyeBVZUt4+IYGxd376vx5OxVRXeIGK3/yzPtIte9aBfyUHj
UURv+zY8q7gTOWS2enLNA0jOuDCT4sZ0//HyEpCP6zQI20Xu1S1SNx4UElSGRBrX
YX38P4U/8TczA7EvbNBu5ZsK6GQENK5dBs+DH4Hnz4A3rN0/pyFAw5b7ewHE2v8y
fCFVsjje8keK8r8nEpBskSgZVqtBodbssVcEr1hIuFlejLrzsJU4viOXd6E7LKy4
sr7avOJjc4NCK0wWsePQ/a2zXT7CQFzUaQpSUlnPf7sK7+2qFCmn83MenzQ1Woep
MK/RPLN9N1NzN/TJMMYaOQNOcVbKKdzzroYXnNpmPqaOsBEvOrzNX+9Vf7gOWFP8
2sn28YxgNlCMnuWNd3QBOd0sZAVn8FRgCj6hh1becrRbsivvOyEW8DRFC7YmHKER
tHQy15RiaapklP2R1dXj1VjxXdJenOPzTIQUT2TesaqWNncot9nSz6MozCnnbOYh
H0JJJDZzJVSO/vIQrUzWwKoHQ03uX+ipBoVjE6Dy/X+06iSL3F41hKY9NSSOIe9P
Xd3yRGXIHsUFfYXr5MpS9hoEg7oJV67hK8E4Q/pd1J0Ho5/Di7qzbWe74a0B+XiK
dpUSbiaflFdqpyP3kLQnH0OPdAIe4pydiO6ccx+Q7XwyPaavy0wLIogSmOhy+Y+X
0qV0TtxmvQmPnHRFr51QiQXZXmmnzGRWbSmnntmrLt4+WiwFrShVPgbFlgjl7lLO
CVhM4i4hgfL07upM4heIRHGxZQN8OOVpXIq3BTJVALp3MiUGvJg0mTmnMIsBY/Km
4bSntRQxHNle7VVDZGfLTQL/2MMIR8aQrXpZTjgp2Y4CSNibdlxS8vbbvyYEdk9s
mnt1F1qMpluY6VNhjXHq9M6khsFtpyVuhsQeYIjEZa7rrx+p9R4iLx6ZH6PtYGH2
Dkbk13v0X/IAvB69U6Wgjoa4xVmMV/XJv3EmxqCHdP0cTzTH9NApntdmZieGPUb0
H6xP8xHDSBADfK2/gsYNTFjV56SKFoTBoqXgOWxE1PtAb3RWJ9B8RkCTB27COUQs
YfLpbW8+L11oykebljR+lNWi/tDpeIZPkjRd0YtxkgJkjRMmFNLm5bTbEap/knj/
yUNdKUv/rYgqS8JoCVd+WvOjfu+FqMJNnFOSpo8iK4+Nv5FUsyOn5i+0asn2aAzq
3O9EN4Sv++OyBNq9zNFAt+kDYiPCFM8ojdwuzXK8oORzy4W1tGQLJ0B+eZdAKKZT
JLGfy+RBcUaMvZo4vnRIYTxCKKnoN8R4co3UpuNYmjSHTWKxi1X7hFvdL2Km5XaO
n27JKkPuSfGedDq0RaR/ct5AZx/RmF5jpgd08drMUf6luzxXMt94WSJC6jdF7p65
k5869PNrJ9+uOyiY0LO43s85hjeuJBMRbrhKWW5qq/IksCjhAy0xBI0PTflEapgM
TlQfAXTqxoS75QiP76uNQRh1PP+fmwR44aN/j5z3wQpz4WNXycrVo06LGmXKXwwz
6Eii7UJv6GrxENb3397UIXpw34j+f711lyr5X9021Uq5DSnHTHyrqP3Y465Mv5+L
ULhBTnREgwUkTcQIxbh7Mv+cEIZbpTBf9n2QIBokPEgaEZpWe793CNjaKozmnNvB
wLID243gsomelohyxy4uTN/AktabGjCS1RWdjE2E4WZoV63R5LRqNAQxDCNGn8z9
lX/x5h/Ub6xih5wzarXTA4MpDFag661CmLzdu09kxbWFElSIUQ/X7VLQNpUdCtpb
LHlLaio2kxJLzb7GMMxgqJA8tR3rDOe7TDB4wRTu5cNdosmQdT1RA4MDJZXXxt6A
xCLsRyiUnGefw+eyJGrChMOiKBe1exVfumKH1hX3CmLkW+lmNiKmESZYiaWoX9jk
JMPsRi22Civ6fgQVkpjH6M3sJyeqxeV3tUVUnue+74pfdnJUz/aduEjTeUZen0s5
RdxcWvdZdlbzEKWOW2Qp5Xw+fELwUi5fRhT5GFVICqXxdzeR+q9eIYecI/G7jD4j
PE4trJUaywy/Ho1LJVMCxztVQRw5r+WnvM6EbT9oxmwagx0OtHI5fL5F0WoYXuWt
U2dA/5GEp52Ou6C+wgYnlJ2iF1DHO/fUm3timxy7oh8qjlA4pjpaFGyJ6OiRjr6q
s/9OZSm8IttkGisXJ9m3yU/AKf1Kaq4Ux6EJ9+omZFEEygr17mBsR/34Q+UPokLQ
Y3rDY4Fv516vQJmKBk0YziabUkosKkqhpg/3n2tHoS7P6J2eDfRmHnXtgBpGEZ2f
j5pYVZld04PVlM3X+sIiH7WpGkJHUY2bdbDtu0QFFFhu3okwuJ+tMNlPY8xifvH8
zLwCE0B5r+6VHh6Ffil7Uk2kvlE6zsp08ekcerikhvSj7wb6jbwfiHerGao19ILl
W9gEHizuU45Ej/7tTbGPZO+3jNwafciDb86q8XZRwjN9dQRXFoabXE799oIy/yX5
Yz8/rUfUChlKWR84i/zqnzcU367JctelEFzGRC4yBJZGeB+a5rVw4+gH7jyvtufn
C558pBXKRcr/0ILgSRjGhTFH4C4nHhwNPvy2Ytyg3Hh/WesXB/cGawgJOWzqt/+l
Ts/D+uYTU6ejrIEf5uXzuzkhUmUVX1XuY9gWLMD7UPEqPpcspRl+IcM4tfWgGrK5
ioji9NpEnuSvvZCTp/a/xtjbxjSLLOqZyWSE2gkq3t3+u3AXyK1toSPlwPUItMtI
hsTtHNUk78/7vmQ+JwAryuIDJGCvpKDE0/ARrTKt3BkFwxtOB8NTBylpVYWuZddU
lFZgx93HzYncSJEaY3UtSUiD0gIAQol0OV2O0gCuGyRKZw+QxintogxnTkOP1I1t
tWf6P76OPAJzunxlAniLkolPsSQM2ShqPS8P7LP1pNgDEMLddCLGuPpSkOplTiCW
Sij8j622YU1yUDMryk+62rpVdXAYvDb4RKPG4W0sG+SSaeyocTxEPvzfV7OERBbg
pAY6S1k7cQ7nNRuxEcs9o7pBmuxlRPZTrkfYM1FOZQXwDH4ljvCGPZxkhPuGfM5f
Sjf0vZ+258Y1yUoOqvtBbqhBn+ZHChA5xA5I83v3vUeyoL0jckMj8EhQnNe7X2Sm
PkxOaVFjhUIN27A+V46MGf4NUZkU+Hb0C1zG6on2xdhcqwMdssTdqW4k9HUXSEQ8
2N8I6VYk7pUH9dZ2vP1a/gpTg3E3medQaExJ5aMkE1WR2DBbY2Obk59QOAlZq+g8
4yieTZZFZhnUGio3cQbFW7yvBpiKlZ3HukEOATT1Xq5vfzHmHeVJ2BSX7JXNnenk
eJOcx9YA5ieLKbmyhb3N/pRXmYrkbJGs8S1/0dRhRcOyInaLaWs5O86tHD5GZWiV
zLnLKSkQ691Ol28VsMDTBiRSgvFg8JR7+oVtvfcE+0NMINdknVqepnbFQEZuD+mq
vXiYkXh7oWXLE1zqTU1kk3vCHTha6lgGAg38vqTktJE4e6+AlMBk1hNt3kYrY+VA
oZBvKVg71bSS8kcxJ7gvf1vXMF9ROgzEBX+XgEMXMMniS60zH5/+b0Qt+X03SFXG
UG9N+ySAOXMuU4w2Qsylp7XskjGyifSAn9YximAU7zTCi/w+sCzFT8PUPdDPIWZd
FDw7lhlnDNDZRJUe4+t/hjyx0101yXRltOHkpuzv3kddT2XYAHF5/UulBHVMfXfb
Zz+y8IGaZbmW9QIhfN+61OD9Uim0GMGj3IrNmjY8zacasQ7zww8fCwVkOQGjMa3B
5lgRfQwsUF/0tr1pMYAvemr/oNTHGiS4x6/eakkDJkBc79IjqmXQqZTU03zupEJL
l2jEeZ47QiDJZPqF5u+GFbh1uJW8kCfqqg71G7QFX/Tl/RmbQNhzKLPcmD1mZXOc
ISRAs+dUGX0QAO545djBsIeY2AOAmyTSJG9Ral9ygzlatpK2DXuwmRbezJQzXVJV
ZNseOH1G65UPEaKdpPMRwqzNBNeXcyQOBQHY/NcIcwMRhTstAjZ9EfbYMDZKjY/M
DdPdGkH6dAZ+kRS4BzQdQ3emoXf90KGEqR76UsI36bLFU0inhIlHaOAufAfyFelM
vRz2O6pGt66WA3IWbknt55F6rb66n0qupk2j9nbEN0w9OpTCaKFx7flZ6QoO8zaw
OGJP1nz/jN0izzsMXn0K2zonxkgtLOxANEHE808UK1WF+TqLW/GyAPW5+HGjInBN
3C14dlhzzFxR4w/dx/dCLgXkILXX7YRGmA+6joTjlmc2L4Qjpc5nwOWbLZ63imST
hr7Shla051mrAxJTVvjlwlDyjzuxyXoEgXlG6pnzLNbtv3VluHlDAQI2kWtqUN+v
B/g4hM4gc1Jkvsn63auBJ6DXZMkU1MODXLrBEK5dCV1uMMFqbom/3W5Y1oiXmtlW
h1cp9m180L9WR1L+SUoK24XhB7UkjIfD8DE8f1KALGJomHhs+pXVROptTsz8rrQ6
TAqiPf0GFMyUrJBZcFO6TUgK3Sztm3mAxgz7MWM+RtsyNjvGNPDfVDsy2hrC8hdM
CY8uB93cpMXRsfmMJVjoPrD2WgoJH+aUUMRMDwY6jaORdzKgNqYVJGZT/g7BPZpf
kqki6dEC8iYSKqR/k9wcb1cfleg5X/mBxtMfo0l5ZYhoq4crT74o5G8BjltKID15
C+Qv76yOifCiQ7jefG94/2OwahdIwNltVJGAd1L/+kL7lS1Mk3GIOWwBoUR0gQqy
rnX4BotzlXRSQ0I6dVxHbwPjz+gHa09oSHq/bfB/HDLXGQKtf5Wwys3FJ3FSQbEL
SlWirQoJIJ0qbPjl7lF2MNUaBky1DWqplpJenXFzowfINPxWgEAwDwz8o2vmg2Uk
P17X2mWnPwZT/EbSOV+jcekh/+TDwAhYd5Tmib3J8K0EIwHXTxIQIc5j/csFEra8
XsTBZhGr7pOZ2zjb9jHVCKtTxYmBvraVDbJEJirTFx3qHMEtWaaZx5KTjvz6UsvD
qZfieIn3qb+42U7CZ/yhK2bCHv+bbnLpiT3Ay01xfUzOROJ2svFhffu2vlNF8A/x
z4ggZ3he8NbPZFpKhPJYtI5vFw95S7kzgstmJf7VGvXdRZ62aC0RETzZpaH6sZbS
8w2eBo57rXHPSlIqOKPaAraROPrZEnGy2CbQca7k3utdMaOUB8wAWF2W6xVTra/k
2KNBmdAHfDh+8TK0RrLnjlV5aIQM9a8PXTOPq+jWVWywPRqHZMfAmziACjJbl4rL
LHHOaVsKaQfzAvAf4w2DYKYoFqKEFZB28MsheuzulkCatC2fWZQu2L+kHlfFivPA
cHT+WQtLBoNUfQUMWiJWiJNUGZe90hJAVJx0TcM14n66DFZOXd994Rn6WE8tqNYN
hSd4LP+2i2jGEF2MH4IT253CUmRg8gT5kMUIMwpXhCpNTSj+pkrlpo5t738f7BsN
pNiUlwYZiy7gZA3+QxRtFBV22mjilHF/ETt4DCgtsqeMNWiQsPGwIU77smbtXWEM
DGrj68mOfVqZFSKXg7bFPBTGyKcYqFczcnffNGlEGQE7PJHOfAvaICST47+Byipg
OZ4LFCbNHsx9aZ1I1S5kXYcQ0Orj8zEwOE+tSfRqRBb3MNGxXF5JqOvY1Vdu9UF0
8n2CvZdTg1HNFs7U+CqczYkgNTxKCaYSn17apFfMw2HZ31EfPrwT8HsyW4WLkC7z
BNE5lGSVcbnUXZ+cjdkhlzZMDHJcn0BPdGvfVhFZhLXfZ8upmBynNv+TLUOhHeYx
eIUZ+iS4y5h0NyMGClHAcp427lVlNLentO2Laz4/f2VCypZJEF1He6IJ4ePqjeAr
ASMmCkyVNo3L91Qa8zhW0gscqanpo+ylL36mFOErgvhSy6QeSwJxxe1jSHUgixuB
2qWBRpqK7BeIPp4puoHWMERtQJLTBBYLHmEhxawlGB0sXtP4sAkKk170jY5hNySA
9F7+JKnXRTWAp9JZiY34RnzhNFP9LktXd98QNUXW44W0/GyJLqX762SUiSwcJoB5
dp4NGSbsmz65GqB4P7nhEDvYMwFQ3rRjRHBYt22bqyKRkcPCmMV8u7onjq9hmbLx
YG1FLrR8LSOHJXHZ4xMgTdre/nEV0ia3SZhsRt/9W+edhHtrgob+U3Vue2fJqFrg
4dVxfEzu1pg/6Hy+c2/nYD1Etylpni+yUEnUGh3vDDuZ4Sp1Tlq6s5xv1R9dACNe
yXb/uXFz3d4fc7srB2dXfd9YkLg2Gq9D1O7arQQrJXojatuB/Vt6P2MfCwZMWU3Y
95qpmPyoTSLh4N7anSoTYWpFkuXibOjZj66MJMvD1uw6oCYdirguhTajtmc0e/5d
vIaC3oexFv8vz6OoZIyRc/HTGV3uyJC7nytEmB2XXI6sxlVGiZO7RK9DbEBcybYl
ELodS/48wwKN5SERtA7VxwdTDMpZSY09UbpUMhp2PpoLw7MyHwTGWbj1NqdZAQSD
F++vHB2NbiP91TV20pZaB7kV73EuBekvDY+GgZMizDiVPK27Qwv9ufBGBvaF3VPR
oXNdRQBg4SMJKI3Hm3tPEGOadmiMYymstzaSC01yRzYTfJP9KWq2Q3UTRfy9QLQS
sFxJJzSd2iRk3KsNBcj/bD0EAVbHe31vonIB0ZYlf776Ulz/8EnZmvpriNzm8/lz
Io73e04pRvx1WTpYJT+MJPDO/vFoiYarOdxi7b3DnFTweN0R4U1hSQPL4GHTfjC6
hPEGfELhOCPBWnxAtW+1W4MQ8euS6ATP7zhTLhNoIuvlseWxZ4dwUYjPB7oPEr11
JoDpEVAOBOIjQ/13NN/QXm/HSFw6spjU/rqJ+A1NzYemiHyjPal9rOhfKmASoC1d
o/y+bUBVbOWSDM8IpyM6TcEAoMR7PkNW4CReN1xyN/4eqDomNmeyQxAS4Fb7vXcv
1lEeeJrZt7Z7/T9sLKaSqTh8R/pgrd81dDJ/YuO6QK6GjwXn6fqELtptvTliJRzR
lJI7toCvygfhgYZTEw0uArALZGNYpY2ep+NMaLP5aadTJj5ae5vOs8NMO0ukjbpH
KFaZJvQL350227AMA1RG0TStXOkoYg13Yv6bHpTsgBD37EujecPFf54D9zmDDQ3C
PzBWyuQqcNa12/aV3tDoqOhLW1XY1lsCN/POnFyvKomIarNisefRjDbw/RMQ6EVA
yw9cVuGA8oQ+8nH6dnBrQ33cbjRYrViegMZN9wFN8olgQ9qEH6G/G0GWzbfYq/61
fHPnO8jX/Axjf6aKk4JuLvp7VGWuWPUr8exKA8DqF/jvIwJVj8xold7Ld3e3xmSj
rXxYWTYAuSgVDFgZtBtnkKHgkxEDGBJhyHHD23nzpQNjVyIiZcZ9YSX7P679+zZX
CBpFrX8QmaWRVZFOSDixejzmrRySg21Guf4wjIfeNEEdW3QUEAd2AozSHFH4M5lt
NaREQG+VxZVx7DjI7wgtmz0tnquCiwPUiVAgRZxYEc0ZCdag4WGndYx4Em9XOOlR
2iHnSxq8hCoJyp1NYQ/smj5PvZXpR/W6WnnAe/mZGY2YBj2Md/rVZI0WjgttRP6b
nG2Ce5jxisZykw+efx3nixK1FBxfXhHFIKgQFOfZzsnxmYEt9E+xE65bMxwmYC0W
9zgQwTEKOxPsiwMgQNmsetuti5OcQcwkfpF6VIliOZzdlh8arVwiqm+QHSueFoqd
prBSUvUGJ97GxS01DyATFZ0L5xDd+BsnU7z0jBxPRaYrShpvTGm8FEiuL81v5poo
DU3Ho93kvNccJK3pTuHLgg9b3i42znW6Dqy3avsrjkpBh7H9JO+pRSFmZAsMjH+N
txthJr0P4Sx2pN7d6U8yX68Uc6FQOX1DrQ0/Q5Td5ife20BYXRiKwDc9PQ3QBOCd
sjIGYmjYdDmbuBEfYjXbBxOfc2gmZ5ItD3Va5E3+iMzZX/2wsGfc0oCWBNYJxskK
QzICUnfnpF4fLbCoxJ0uiMocZUqsc1+WfMfqXabxrJRKXjkHJoi2hqoDk9Rx8al6
/7DX/Xt9NAL8AXKOXUShF/nZ7983AriualvF68gZpQj807rBscl0VH5uumG6EJx0
RFGZXsDT9rXDUhQVw+hJpjIlyFbW0mfMCEDDim4RR0706wNYjkw5x1mh7Fumb77+
VTV7nl/VSdJDHsIXshk3ALraVR2ood5av/IIFedRkeWCiIRgbAn54NDARPdIV1EH
RjNfqK4ZgSjMM9J/rFVFR7D/vl0wqF4dT5aiMUKrGkzygkpwliWwKVHJkEh/eb8b
PkGMaOaTPlRjQPwPS3iuELKJwqETg45+CTkDrrJrf0gwHkEjccrdSFVE/eZ2mZTb
MDAT5nN5JD4f8X/dv3jfQDhc8vXoXXueFOLQhJ+wNdRkrjReLGaATnQVXlt1geqn
BCOjifKpEwbO1I1joDBlB0mC0kAZEoOTjHMrGYErsPbmj6pi1REt7xvrm+WpZvtD
D8hpoYhDMGam3OUenQNbL0aZhsGqc8lroBTwQ3f1D4L37WXtXWAkZs6x96wlS3t4
avQzsxLE0sAqcKBxSOiatndTUhTddIOvtPGEkXANYVXwV/9vy8Iexa+s9oHvXTtg
aeOlCvvF7QObGgpqvrZFmzU2NvtFugstbxdNNTpgtyoZbrDN6qpfbFudzLlsuia6
Mlrq+aQoRuNNHCnlM6eb0JwpjqXJ33rUJFUFsW+D7tBMgHrPP0S6xllL5r15Wl3V
RqZVGIq/D4hqtJRHl1ivyYpDI6GgHQElF+ML9ZrTWzP71WgU++w9m87OdFnswWZI
JzXMPMDaJjSoT9JoE6gyw4dvvhOPdFpkVUfrE8zp8kEue4sv7PAW0b67leZzuUbK
dkV5pT8uMqQLpqx5Ov7hcc8aOTcyYYdh2BXaGWGM8U98EPV003VOLejb6IkJGrDe
fdXlFaqU2CGuLXWaPpbj128S5Prkmt+2AV7r9fSWIEJu9CJBPW3lhIvrsJeqpLlE
pN7q912Nz7oCY6gpscbWZ+96uFb38qkeZnZgsLMdCSXVgognCdwSeIOdtXAULhVt
ojbsBDZPmsQCizu4SDzGhUh249ypOPVllJSWDDD9XVBnp8gtBcNR0YS01kp+eOsG
6b1g4WE1Z6qPCBbE+ljXj4jiQP8niF0sqfLxS6hkMlzv0KCT+dGl3NHgcyabsN2H
7Tm3xBvYFuvIOcBOVIoLVHK2tB3idwh5PCDq3VKTgfuzWYHs7t+65h2NWRAdutv1
Phld7iv18dtOn1BNtJqO1/0QesOk/V9lTxL9ud+572yr+UMGNkluXzdJECFeKV3b
7zQ/DKCj/qV+VGiowpTYm8RmZu0jMBXH2eoeD47ddRWUAmXXsGGVA0GhFsQsvKN3
gVdLWdV6XiAK8HaTz9zj6UqyQqyPqYTT6cO0sFDn5IlnVFJSeRjYNrthhcVgixvZ
o++XajFH/R0uLjlOuvfzFgJyJrgCWn7+pRU6qggIOLRXBcLwDeABO6J6XNr1qoWN
5cx2xGU3YGZow+CPn3Pc2oR/voWKhp/2xYm0rxzsydiHW5lcVCx1e21/tab/hWid
l1U9//9JZbSFm5XNKFcop0TfTRXkpuLSzyJxm6ZqnyX1qwznv+NInn9aEKczHSjB
6ntu0bTW1eCAJa7PYyNAC/zg64DXhWMuNHoeI0eIEwwuS1iTWExsKz9N9LJb6lnQ
3yVxrgXkyQ5cCxAVruUrBt6BnrI9XJFGjZ3RH66+Snbzr1FJa9yG4H9hHFKuJ/oG
NctDdyD28Wb23yL56/yhOc+Y1aJYCJqCmvdqBFhP5jXRzri4cacBTfs5W0vo9EKN
Vv+Ac/ZopgXbUNBpZF/+wbbCvZSp/tR892nUyEXmFQ8e4TsOj5yLibnby6WItZP8
wxRzvO8bf9Dgtf5+SkrGkfrNYyWuuOU9KSuOga5/2yFpAu/ebhlbTOXAV6jmpJV1
lPxKwJbGRbrO/EfIHcDHOOsYUhN9lS8e1UZ/2QLIGFdUZppkTX1BOhpM3uhvlnSn
CcYlvaT/nEppOHrqel8a1jTAg52mDltiARUxwJ4bYn8Vv8xSc0muXtCPKRA7mgX1
a+9blJONwsvgtPI5+YwTHIPaK9JBGdOdL9uMwTrS7txSfuAB0iVplMHPjBAUMZYx
AJafGexhMxIqySUVO8TW6ZPZirSUyDnDpP4pUjYVkeqlPaNZ21wYbt4rrHIm1C3n
wyl4HXhlkNUJ/myEtK1cW7XPYtM7/ggzYh6IIfRjlHpbNxar+4bPOmVKAFhG7SHW
Xf8r/hTizvQhyR61h+89iUo6XtALr8CiIz+Vl+LeagLlniYfrVKRxI5BRAQZSqV+
BTWkR5ijbybjZirk/BPvrF4HIef3OGCIDqeJXvF8ZnTYms2DfYBB6m4aCIuAI/ha
MbS7z8pyVzptf1tj6i6WoKw02Kuep0MigCmx1LVkx26k3rXK7sv0Eao+GBZ3sKQy
A23DfQMzojVBwFYvBOsrJ3jEmgXT8OQAQ/Cqnuxi7sJKfp3ddUemPCooTbTThHp+
jlS3cZcEUdKWr3J/B+fvgdEj1VSpT3sBi1mcQeRedSBbiV4Szw/ojdSg1WtznhC5
0JSiKbSrb7f7SkPyZqzqX2/+ly0ghOitltg1hUqO7rNdrPf4MCPBpQfLkjTvj3zo
Hz1PKaSbs5wRPOcyehAvKpPEYEB0qL8+TVkhmRkSy7NCgChdqrkUCFpWvGFfp/Sr
leSgFpb720W11e55lSJLTXaHywVi12BRyIhBjcCPoajQk7QZGUHU/IU0AyjbXKdM
E66PdrNprOg+T62gbFr1ZJmtxrEwdItTRArWbGTBS/rmiVUk9uoo+LaTTUnyLKG7
RYo+/HrHQyaCbwcxyby3ZDNs5faDvc6JOquGbsjYkg6g1M62t689wXi2S5cvcgln
/Pjs3+1GGhnNvk5oOiyVbc+uEv+YRt3Hg/AslVQL2UxagTddR9efHZ0Wbyiskys4
k5x8B9rmkI+Wktwh7ggiXALT3uIJwwkUZAClMK9ASQb1mVGjPf2DCgZnBSjbK0/t
/dDme9ypcJtF5kFUb4G6n7us+Asq2KriE7LBK9rI+AWCJDVYzmWCRGnJe+zTAYMC
E/9a06MKpeKbvbdQZ6y3vQce84JF5DTltAUvo1/C7kf8T0g6fJhpC/HfoOujmAUH
cADOgIJdBnUZK3zwlCB4APorx91eH/WBSKV4Lbclv4cSNYJryyImUFA2phZ3nMip
GXzGzxtnIMkokpL99SsHM0eMLU/ON5KpNrkd/iJRDcZ00ByAP07IbG69UtD+PDg9
KrwvhXNMUiJjy5nxomgclzaPEdcNCW3vD+9tc7G8UucYMHCYQPVdR9TThiPA2f8P
qeij/UTn5aAdl7KqBxcH95QYTW7v1fq8vWVoVjKSG+rfqhHmcCRxsWuSTNnHrSe3
t7vLiBNjSJD4vt8GV5bWbY9uydM2jL3DsnuhdFSnps6bZrKJafnGEQ/zNFmuExde
LLFkoS5xIe10Z4nu3PgDKvVaE/t6k9iVbptdmCbE/miUiX78jml/p1YLFEI9UZhX
b2GJeCFXfN+u2EKJhtpj3NmWiFg2/3efcTGB+yvQVGh/bCAlufPP5EpK2nDxK7DF
i8E/0B5u+a/CA/cHs7L5NWpMfYP/FJylTndgDHUgUb/WqVqOEE9nDsG4lMQl5lvG
+B9mm7Fkk33eJHB2phrZRC8j+aRf6WbJjfFfKIfVKKhxmuDmKOHrVuamTb412gG9
GZl04TMG8yuru6fl4GVrNLJNBkDL6BALWh6NoR7gPTnroKy3AfYlKoQZaq9k88Bo
eYWTclPSIDJWtBJNNcRrHcDwTrl3TGH/1DYtJ9bGjd59A+2A4/ZECLauoWLjtbrK
X4FspV/PKmUortgCIlp6mys9TSyqxNcrwkNReBjPIVMLfGkGYIz4v1JMqyABvA5N
hDOZVYhUHyPBlf4VpB1kFflsYY/Wz7EgoU10IDOSK3V5P6k5CNVAcCniBwMB4FmR
mimt5oMtr5DIJVd9xphzyPybwnIozXUJQNUKo8Y0Nc418vWTyTuQdg+pGvfUtTeJ
NlIKxNWT6SXpwlQGexZGhlgxQkhRrlVsjPKjAZOyGphHHAvzl1WQYIt60YEyiM0m
NeaXr7fx1tzbQHOVQhzJu00dNrAUwSEDUU6syRN2mPlb1Y4BOeoLOAgKaNIvnVmr
mH5jN65UGp/BiL+dobYp0AEzxY/PFgiFi5eVDne+XFX3ERwoLgqai7fWhEABzJbd
B3EnqT1OBuvxpQ23pE3R5R/TEuu8HMtB4amA5n2NrOKAQL8Rcacmvo7BTqmsxuV2
ved9p1XimzgOR7nPyaXOL8yxqHFKJsagL7XRwRbbKoTW1eDMaaoZ9vEfoC3j5qcV
vuYR3ePeOTjZEnWOX+zsflfJWzxyXSwY/j+eyWSxANzX7hfk7061NkJvTvX7qnzY
3wxywFbgzP3fHimnL97veHkpb+V3+c4s0WBDSOqzg1d1WBb8ZoMhNDC4clnvAUuj
u3H0k+YxVXaazGoU3jq+w8ye4DATM2Nqnz3mbkkaeZbZ4+wbTrkYDDbPU6z7qz7f
lGaJesRuAtXJq9lZYlQ/xHWgraBtfWk1M9HXpsFtph2jc+4YVU+p0ThATlLkffGO
ptvIgJM/et+PAq2jBVwehXxLD9D73Zw+IAYGfhLEK5UCv59QaRnZON6fSLNHuLmS
sskIy8/iiqTdHdHvu62/u3AWgWNuyNBOzLfQjoDqVAwa7IkxQw2LwHIJdW3xvL0O
4ob5MF8AEqSQaoLFANO784q0Mmya8WepLQbzJW5fClQSKMia7twzYSSjr1jLdI3a
zi37VmUX8OYsdB4eUEqwfstIJh5UrFBJCANKk/xr3tCELgf83CkPMnwQ+vCtlxd+
Wn82gil/+EK0B/7loBpp8Sk6QAWGH3FMHJvmMHvBr9fz5SdcAgYiZojF2zQQunXY
6JlSNXl/QGypSvm4ydm66of8MyfjB74xWYAEyV3Anc9x/QXP61IP32EJRtbiM24V
6uIjGRwjUtki3o3afHff4a6hmu30URtcu3Kf46d+ZJyZvBl0csXeyOPWEq7QtbAQ
VwOPk/AMlg6b6g3LE+igyoYiUhBwB4nbQgnUPLjTn+OSm9fueE5NzK3Homknt7yf
L0g/2wNDHJ4KgkgRNSU9o205W5ekoXWtmgxc9/8NBgI0A7IUeRDxx8FLGFDu54O9
RB8GygGMsoHNNfm4WK1phQH2NzexBT3VtIGcVnynIQR2EGySeSQRX2cNKSJlko7k
/rjJSgc6Ezu0GJ82V1MsY5KyN23/KAEy4vIXeH7ZkcxjTLk8iyItqGjDT603GQOc
IDpsO7Cd14ZBt+zll/wWwg5dHG5KGSxuTdmHbuxia1qagmm6gp3UYcYb7aAMDCrU
rJv5WKK1g2TcaAYte6ZY38BBYxAkcuA+t8HMsFNRBtMCjnTtwh+muY/FFOAF16R1
f9H6Rvx+4S1aGBrsw/8dtc0a9TknkL11rcn1GHqsCPGOEf9Cxfk46zqYUcCDJM2C
FdxqiPQez5MII+cO58+L7yuqnvN2tr02Hy6RK4TX4sO4On0jmOJIMDk3WNM2cbbZ
Os5MooFxIaT+m35eV444TQ10YzTgIujMNIvsIPuh2qWUwZlYcdKAaRtr3I7dfRv4
9/FoQguYyum6EXptLc7/D4NyQx5MCjeGZub94b8OZoX8IxgBLvmVxoZs/g2WnJNK
7Y6kJyI2s0mAwxyqhOOgoJahDcLANUGAPBHG2k/9hav9dKw5oIFm6zlGn+g9b5Fs
Ghq80KMT+iPDGgreQonOfyV8eDKn1pGYhOX2QnlUTVqVQgeS/qnEQNIyiocgio7i
KJP7Fc0qXKtEaq30+Z0kshXVtDr2u99EKAcMoCkCq3KvyqF5boQpNgeLJHPkTazd
BkMsrq47DrhoMvG92d35gs3oKIuoKVQf8XPnUFbHpwLoqUfqsd39sVU0LAuXaiaT
/mBOlx7vH6j4lwaQ18Os1uheuWxVPlouLCrSIFD4Nk8yk/t9MG8TOWKMBQyUNEIX
CDz0VpZyNdRypAj200XeDjs9Gayobq+h+avcD3zjW2b1EknWgxIViUvEDw1DqJVh
symkyBu1zF5PpF8Gtlq2XloCLQDDV400YWgltgdug4KDxgc56mfpGnMmcnfwatFA
yxPrUP9ex6JahFMVcWXfDHjNWC9ZPAQq+X6rawX0XS8caPEGY81hrkAoNTC4+8li
z3/9ucGY1VQZfNWcp+RdgifX5k9wPfkN7KaoODInL3kQyv/yeQO5skBIS9nb8Qpf
Np9i1kMqRNKMysSOsKqd/NN7d6VcCHl2wCy8IhpSOkMzjTgbW6dpQYgJbp1VG+lJ
Tw7YmofGoeDWiUKFq3yGA5dl7E2RIqVIwVM4JAe8XDWIUyYVkeEsOMWkBgUN7ZLS
VHmCi5oHYI0GIOJNaVPHtijrajFGQEESpcRu+rnpEWNkv92qkXNusIShCuIJsauB
J1+4POqeGz0xA/PU24O5cB17A+v/NZU+VNALq1JvCKk9UmrITuv7x9PhVxDcLp8B
aVQfe7Jplw2ap67hA05qjbWqlQMYDyyUhmXV28of3o7CJN3bLmou7OgrYk2d115q
+xATHFpW5ec38K2LfRrW1DKQIbsvjFtxBODMMlf3a82S8FMyVwADOb3qtvv2nIeF
WtYOwwMj3GTulQzBum+e1417DG6TewGdhdFH4nNmgJq/KC7XwTbhXF9pl/4b51/0
WSi3GJtJesJkPjzH8TrjRhGVSJetHX1FdK2F0OYRPHzfS+m1FE3fCqcdmpg/jIBr
9Jo+2xfsQDiWHx7slryHaf1Axp/5hb4KZUqAj8jS/p0pixf3Mi04T5MPeCKiIoLy
i4Ly4OQN7kQoRXEfaj8TcUm9xS59ZdwbU9G2Pe4eCdxqga/w/yOY7lSo6+pWwY04
J+2X8bgYcItSzvgzay4IP2HLD2JCtnbVdj7fVZMDrNzhV6FtMCeVysL2QJCqIET/
IDyW2nXPLYtE7E8yUa1bdxxun4cAmAtU460/N6E45ibEuD5ttcQQiPtFOZo2fmJM
IpTA7aJz1b1DUrITrej89kek79xY5qicBgrPkNAY0BFrlTAzZOraSRKzpE+ApryD
Js8aGs/Whzdfs4G0PjkzpLXLVxcej072Kme3pRWMjcp7EhnqVP4vRWd21WrNJu93
AuY/hmxGeKaW1jsqdumc3C+AqW9w2b18C1oH3ZD/g9cnJC7Sd8b6kbDHQJNXIUd3
UPtJJyb/2uT5If4qrwiMX812G4xhCElBmh9okm2ZCpxUrAWWlDpbIpYMc8+fdJWE
SmWCSwEiChdMYzZMOuVwdgWTe7+D+WSXi3rta1bTnryXksI7OuUW9x6fQGW0wJ99
V1xQ42yJ3OYQGNBD7mnu2+3iY3WLl0N18ykgvl2P6XXdtvcsunR4V06fdcy7hg8p
gIgN0XZHmXrdwnIhSnHJVH6wiEaL5RdIOeSbfiNkQQdAdVxsXbDPB0qFq0Iu9u+J
yY3pOd4NoVXxXsU1XgGZS7KNDt1xouf8MkvfC01AodTJ2sUByF6fPefxKfYuZ7Jo
cipPMJ+/bHlFaI0aeTUCvZdc12jLRLlOkeOu0t+ti4BIBkmf7i9BczgUv2EoFnxD
ahUU/o3KdHJXZS7N1AIVuOIy3B7kHI+HzhAVFWvAWFYmARZ3dySkhmKvlRdagvLS
FSEOVeoras546LzJTk8bgDr+MUBe1ZMsdSrZEcxkUI3IKKR5nAUwGhGHUGzQmOwp
GtE25bGYmpSPUaU1Jo+MToZ8BSFr+uscCR6Dez5XzCuiNDH3qzJearo3KPks1oCk
mbPE3jZqWZv4HyiCZVIJBTUibwEKtLPnqDkWJg7QbM1WuH4a4lUq5eFVk985OITy
pd45TpWJiTaLdmwRB8UuVg36/o/QRo2xO5Rz9uAvxMihtlAnFbSlI1xH7j1qVAOz
PAw0CAuLGKDpnwuTatZVp8S68IfNKjxrKITNeUnoEhcbbgbvfCaKV/4YXrKq08wU
cJwyvt5+0y5x3a+Qp3pAIk/1anNxcFbtBDfzl/vwa2v5VOrtMHE+CvAOGP4XXa15
i5riXKIZPVQd8ibJBKIsNe4evpvOAGFegmSCTaGgXYFwZZUPi3KwFqOvKkZE8Ma2
XmsD1M3xBx6GhFsXDP+GtQsYYH/NMioqAUjNTewasPx/7lpifJd3eBoy2cAxc0lU
GmwOvz5WdlHl1QKmN1dAEPWaucqhBBWHvSnDOACaP2/A7R4YKaGt5PhYyZ+gsnSP
r8ouVZiBU6qixOoHKKqGU2UtCfGkuPdl6fYgrcs31xKyDVIvHPg0bJuL8OB8jpC4
zoZNHJmUNCd4LsbzarUa5Z3RxCbmPGijIlngpWPm3GT0pCHBcZoY/KMBUlelQV0D
+kVKtv/1XHgNvgTLd3QwmvKDzt99t4WpQXc/zCvusF6+JapkcBw4nUm45SDPARdi
W1n8XrW0nELVbkN9yPT2fXnjwpSQJPNWkINRo6SIiqS/tFa5XC7RkTLQh0Sgewt2
tICvb0nycHgfTKowzu+aa2hJJ5bXDvKoZ2IipFqX7HZzIeeSqUpqQYIdVDc0tSdx
JXTeieUzsJ0hw3SUbEwU5JwXjoUHQP5p2TP4DwFIWUg40PRsXxYMQQq/eC1zd981
sxJ+h1FKChAm5v86Icq5NdDKFjbgdC1QXaRfl/zZ3JiAYFIvfjD6Pk5DB7i1sdrA
Y8dxeH5pyWlt1jh8g12RlIcQnQIoNRV41lbtI0KJjnWgWeeNur2kumEcZ8bNrvj6
2YRAJguarWPMa1xqG32IXZnj0+ocWjiz5aKwDp9f+eTOHNRT8djvwqv/FMljylhR
ldht7B8bfAA08Gc8N1qbKVQMZFYjHEW3/GAQGfFoV0VQNVX5VqeTDdKE5ZnEpIUO
kVnU7y5sDETEVqrqaMgxPTyW3rgeE0QKvLxGL8JTAMYMzTgTeNBnYFjmY8vGSgkg
hEphHwGTCQQKiouTfDt3tIM+Q8XUNOve6ZaD5Qm8QZ6oWiJ3SffppIUba/ciajiA
dbqaaRmdI7aWE9vJ5nlgI/LUm+ujuy+9Ktn54BN0f+VxA6zgX3s/DpCKcDDtKcaj
ZWXR9GmTJ2mXvNsJe6S8RIZgHrA5C13f/onxWREN7mWRS4Qw6x3449A56ThAUZZ0
RV8Ahg7YUn7d+7tHK5DsvjZwa0oq7BAO/N7Js6U579JLWaAiXI/KsOJMlgd3rxaj
bWrCKC8kFcdMqtIWwlVCW64/RltALTmq8C6JDCcPf2jWMBAFjn0JVxub0G5nlop8
WZ6Y9qE+Xl/kmGLbpdY5Dha6JUZF2VgH6tTAkSs7ac+LOVCdGHECTg7RIGy0w72I
XO5geF593eAl9xMMc281FAWt69QFCkONx2Ouc2mRJwp6mxl8cgEkM+MRs5d0em4U
oyTJm1hZKhuPx1qoJGdITUq1ZcBnWOXUn4b2x1FpxUGWIL+i7HlW7Gbm8W+0iW9W
flBJz6hh091zolVU6RVvZzke9ahlj31eOEGN+BlRLyRnGcLZJODFYbXLwZnHk0cn
vaiobkboisFbO87RQ/bKjAk+mOoIUuHq9KixaBovsEPjutI1P1e5jmi9GnYeGaPr
iP74CIFPFRok3nronpucguw5QWOCK6M79OFmLdd+DJxS354l2lL+JBOuC0sD+Wf6
2BFdCoyj8VC0bJsSbYzQqBv7CsBKyvIzO318q93YUkLpzo/7zCof9TnRetQNsmVc
vqUCDpw1BrxhdFJ8ACihSdDIwUEonaSD/fa6weBhHkRqP+BYeM3Oa23HpR8ME59H
V126Z+oIPTgYct38JREQXiyFW+wwLzqAZlv7fMWNcoY3qpvaL6BYh1ZvsSN2Rzqy
Ya485NJxqpeT3ztbWFI/BzR6LPQ9ZML8BjU9C/IzorE=
`protect end_protected