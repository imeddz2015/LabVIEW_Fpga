`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 25264 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/9huKRhRMtvnNqb3Z+UU7TahEoHV+T8U3P3ufru7l1O
3DlgtZzb9QxCbOjthp9+wDkjygH0eUfDrEl1ovhZG61uSuV6xynAqpK54/DuUkIa
uF+2VhOMk6smVg2/sqE7QwCJludD/8bU1ei05T1AVKOP5oNcqGkbGQktlXhPIOLN
VhMLZ38KEurFjWxCjWJLpeGsT5n8aS6OscYuFMF41dvtAAJ1+eGPLZJmftTAedI/
mtHS6/O6JpuAUpnEt+AH4k7SeQNZVfYsDNvRkcNjOAm4oRK2LmWNcd0A4CLgorx3
9WLAL7v0QvbHIkeD5UfoHatxQLyDq9Jdm+/b5NXNCiEVU9RrrvOdbMtJQcg3PNmk
2DTSU4CwUzNy7WEWj56pdfVMLWdPcP7pjKcNQ3uFCgmSuimHljvknazZ047GjDX7
cE0spJaguyCtPkUcSrCdHJk1IGv6kD087Vwi5w3mMl1sLUCd3G1xLCJihyKisEmw
hAB0ad76ZwAdQ1b1LRF7pKW/JAIdsP4p4eB/L7/A6ncHVzEFbA3dW/UmGN6GmzKF
p2IyL30mEzfQeJCLjYFivkfHniqigVQr3tsqkHmrnnYpKNsUPzdBW0MbKJt9NiMb
V1Ob9A9+rveLEQ4c6ZZHbTqKcwB9QFxMLuTTRRD1G2Mf61yQwo/3c4bQ70Iu7FsE
+cios5xxUpISBTwckAGG7wamZy1bbOxV9WZiwyGj6mzpjEen0NIuPn2xzcSCeDHs
RjwYa+u7NqpbGPCQIXkAuzsFihQG25GmY44dBJGX5gfZhtiR2jEXAieUG60gvBSv
6YQZdhmx/+LV4grvq7FANZUC9iJg+5yfzdSJ1wY3lc1MUKuVoa3rAlhdAuZrwoxa
hp0vjcFg8VrDbmXYttMHaZD0Mqz9lHxSjLs9Uo1Gl235bdDQsKf/w0a6iFxms9dE
L0RBtlcgBoKhbMTDnwy3q+hJRY6Byplp7d4A8tRzEgyngMDsnTVHv/cWvaJrc4yg
pPXupAQkKDy4aCFw/vNLa4pLBUsDVEaf9XWxSw27EIgR/SU0+gPfKStVxqeGc1CN
fbft6S8TDBlr5Tr73v9qf8P59Tr/n2es2lYJYhP5NH1FeOS9zLzQgp0Fakx95RP8
62c+IvW7tsPJmw+XCCPZQYUlsH/eVgDidgL5sXvPTdO8/l4tXPakyo0uuc0wbebF
DtdmTmeI049Dai26cA2Q4KY8UEjTpqXYtHrgvxTXxr4Ow3ItrvW0UaUMrXnzKqwP
TAThRCMYAjzANck4zVR7sJLB/xPJuzca5AOKwEGqGDM9VMhnKKHmjA8XPpfboI/B
DbmJwYX68An8vwaK8sv/URwHIln9V7z3xD6r9xzlLhrlWNYMQjnUUvBxzpU/KWQB
lvCRnWCkiPonLOGSJdoYfFiSQ7afXui9jgmxQdAHlpAoPeUvdI/m2Gq9PvRfeROn
K9H50DaIn4zpX4vaZE+wtbeoetq3IMe4ZQSTqwdPtPhfqkpdzyyKNawXOqs0Cn1p
zFg8T6l55AxEL8MrUGOvEg0rfmPO68mw1/6sjzJEW6UdTM+RvK+dqxfHgB6JyMv8
XdF3c7ffMeHv4escZ8Z646IhWFxHEGrhQAzxrbhxWklRMucRMfvTfS9Y5PbH5WGS
qMbHzUwLm2/UvH7k0tq9lEW9db9TGqmuWA0fXkk7Kk7ybMTi3ljLlcg9wIGl0oOa
F3So4txM4zXIp8cmQo7AwNuK3XEPDhF2/J2s0vO/OIowvearftBLh+Q7AweobgBf
Y/a+ITDTHp0dYz95r09h7Nz2nlio3dDfqYONm8Gzhrtf16G+kJIMxaOODpEhKyPd
16BHc1+lMewYhjivbiqMZ3geFkycND97wl4OdoVDLlkNSjxfeA60vkLmGHhE23u+
rWF8fYhd2WCKRQSAKz1kh8F61axcFPui7lTfaWKEyVxafP9P18zA9Lg9OqJyDJei
fZd3jzhgLV7WDoU1KyqxL0pUq9BVYIgo5y5uy84M0BV8942QvzkxppMyCtHSrtil
1XS2ArLGkrbEaHqxe9c6G+avEdICjHDd49gTfUZt6S4fERyUyRTDG/XNSRtPRRt5
Z++YpD41fH3dLfaYg3LUw633OThvor2RJLV30Nuu4fPaxCpm7ttVpDTKb0AUuFyB
gSIdzudwxz0ooB/u2mqKPRMfTe6z948jupHfml4SuxYu6D7VP1FRp1zdb9mel4m7
4XjvMMsXuVxwdzy8nJgylYxa29dWN/Yz5khcbuPZ+vGXxFRMtWYWr9lZblH6WvCP
g4tFZniA48dv+Nq3R6e8LAUPfRmWwm8Y5Mukw+BDiN/qJ+c3rPcKkxJ4CrDQNdsF
7ed3C+skvxiYEXWUdeXrG1qMrfVXNzsnpIKxZEBWqZRYkwT6Sr0tRyA+0E8EJZAY
7yZa2T4RJ1/+RlY4kAUFoVqqLt05ZjyuEshdxn7l0gPgwM70DiNIicUIEnyiumjx
8cPAIMDG7UrwniLu9mjBHXmmMLEsPonry8MzhmIAy0nfRw6a3xjI2bAM6L+Omc42
A9Pa3wnJeS4B/V8ZXpzVJ7Ze05xX6vBdF16uNHaQIzfusJisDEDvzvqxAVF9a3zg
Q6v0u6ROKuEXAIoRQWbK819sBU+JDBparggCp3yy7rp10X4PfwvAfVENLo1QDndN
dl5sgNjYRBovLLTNswQY4DEWDhQ4WsNw7gV3rVMJEUUXREDtrJyxC2eS1+xyBdIS
rS3EDaABcW/JVQv7zmeoUB6JDvRN9quV2Ckb3RtHUy67/TZxhP+Gh31GnVJJcnv6
75ptUBgrAk1N0dId9IeOKD/bvuy21arzT+QnBKkWKeXvypAQxc4MchROl/378Ni2
Ztibk2AuH8jKKNYPgJGVqmaku3LlydkcQCPP79+s7q7Gb1nbl0yNllZhCdnDFw1u
1cIeJ6oAQoknRxM6Ke9Wuwimj4IinwabkD/h2mSLfNZhDnQopef6WKGZKwaxe0zx
neN1QDK5/JuVmdTRLWKzzys0k80mH8JRhw7t/kV0pbALePx2C3Fn7X+RtHC5Uk07
0RO3R4CQZh7YPsfbbSujGRb7CaSc2SFE0wfehtbN6RTS0q3QN0WzRBhNYt5Oh3dT
s16Z3C+Nw+w1wKB0a3fmEy6Pz833uKb6GHiRD2TARazttnnSz0rhM61ftcQSlZDb
/hAC/L15xcx9q8LGP74IPVOFQB2b86KjWMT7Uny9TbB7qPtPtQFj+ybx0zgBhTI/
RYrsNdL1pagZessf1mQIWv8RsZ10L1S7+YfQpyxhyMxGowJXOM9g/ScR/YZBy/rM
WlQxIOXXBpUHGC8JUK8YffCB7OqqQTZsviOA0cz543JFQ9+qkx7jd7RP3E926G11
FrZ/t8ehaN0xS7xs9ATSxHAWQ1+ucpfpj6CpQw8Cw/Fn5o0J/VfmPEwuqn8BNYa2
4lDQV9nhW7RBzcBO5mBzsph9vxSiah3VtHlxGkaZSSnIIz7X+gk2LWiZ1on1zWT5
Ds2VqzkDAlLFYSgA3C9sybHPzvBoD1rVFntC9BIxe2zGG7TKiUx7Jo5ZDB+PnLWG
9DN6CEQCn5vaxcJ9/nmvJhnp/sFInvBl2nAtflDKrkFqRyfMATgV7drT6BkRGpX9
0IsuP8XuPtTGLwsqmjCocFFDj6sWMzj1/S8uTxc8zSlKUvUN+zd0T381XzByO70S
jG/vCzdo6wN+2uNeOMsBMfTg6fZyi3dVkf80IhlmaK433O/UzT1QMKeNDkkrKRgm
Ak6Spz98DimGaydkB0BJqG6EGd0Kqnhcx4oN9KkVVbSQGxBt0Eqh+GuWuZdLY4CJ
+U7uEDZt2weJpEPTft2jZywxkYjFNWbcmeUt3At7zip4Szl0WSUOM4ryQueyqMv0
j10rZfoAtViBM3DDW0Iu9RMYbCf5M23WHuPbNaO4rVa2wbGeW7jatkL8jbZWm4/M
y9jmxqnL6CqJln+0kmQcbnCQM1JXz3WITlywsoz/dZp/4pT60EXjYG+Y6QHksnTu
NsDd/dQN8EGO3OHq7X8xo3erzzAiADP9X8qIoNEVc6+sSTYDoY4blAr3EWdmYinQ
gnVEeIFirE3VNU9+oaVWdZA2Mru3pu801gvpGWDs9q9ki6UWaze5Gplar4+3Lvi8
N0lxJLQzXvvzBMaFqkJlxSR1iF1HDwbyrXS+crte3OeTblAXs5L7jZGT9jglp7zy
C61k+7T9yCmib8uKiZN7Wf+L6iAf9RelvHLvnBspD+dWba0r6Uh5YEhfF0bLfGQz
T/FK+x/C5uWkz/h7CwE7glV8DSBiABgrpdtZ8ugrFscr6/WKfWE7ttF2eYs+jqh0
paO9bGdgygSspLzLJRlJQqjZDdGAMFVW4SqUlPlT0RqR/R+UKJDl9CMqQt0lH6tj
hg1M62WkGKdWl7czt2oLQt+WwG2dI/A8jXpCjLzrXkW+RP0NHnep+umPDTIDLhR8
bFZcviHo5HhF1MEdFEDNbUCR3CE+d1+pCaA2lBM7aL5kx79I4CGMtij303MHL9XU
VE2l54lbb31EFQzYjSPLJStWGxIVFn4V6a59lDtULoFnEL6Kh7sPwWy0ZVBMBwCB
YXfgCtPxm+aMXJjpDvl4agp0jTOLUAckaH/yqCkDugkY3aZftWNRH+5o2thy4trq
9RFRqMtosX2EpCNUAWVJkeScK7c8fx88GuRU8UeZ5wOKaAcYvYG1A0ikq9HNj1wE
MUSaQkgxjkPfWxeVClFaQLDXd+ko0bK5m+dBGgLV1Foi4hOJHbRfL5p6HO80xmBj
lxAZgV7sWC+OAjmiqMrdkMNGQ3cJDTtZgKrD/IFAtKOH1wmceZAEKThYbI8dXpk/
tJznFQzpCGyRt26VbSc0ckrTpuH4nKRmf54FcdwEFCjmLmlGtMxN/sQSbghwcEu/
CNwT+3wKxqwLZsk/xP2vy60to2yELuujRoP6KGT4BVkJYcRKM8IHeP3zCEnnMee1
Xffj7u5088V/TrSDpf4B3m8sa0aFID9RyGpcG5W5XUj3IPhlogK4wgrCvAVsNPw0
LKR2Ji4f0z8Mc/ijYNz47PbxFvUELu9GDhOtt7B5+jrZH++vfA/4qfnJWLn5lj0D
vzBcfFsNW0RALrmxMCjvwizaa4gIbJrLT3DvRhwYqHZfPM46AOzgG6GQx2rItQNJ
LIEU2xtAem5HgnsPLo58Tr+f2VVsekZNXEbceyrQuuY13pviFB3eOaq7ugINNQ3U
gMS85PV/nbFbofcbnIeKwESWDFo43bJwA7n0AOIPGjlV9+BxAC9E+4Al/j8ZQBvJ
q1oBs+Oo0o0D+BQ1sYY+i/AbGFJFGoE61hmtO/5oTaCB/OO5dVI1PoMDzZjh7q/C
tnE4IJRRCJqSagR7444Cn8v/kKpq9n4f1Xwrv3ARGeZhK6bICfszkGz0AtYzg4dl
+GC3fXWRlK6NnohWwaeBahD7CIm7lcWaJPCLIKwe//CNGMXvPeiu9JKopwYXXtyl
OAW1cQF3M85HS13Tjil96lYg/Zx+yHQZAcbBL+FNzmm6xeMsp6rqlVQuHhICMFjA
WBxLljnAV53N2NMGTp8ioh0bCMctscVbCjS0fXJlYUQy7akep/bQ0LvpM8joi8VP
h+xMrNvHoGCSF4Gpq2Roj7iotTcO4ioqWNse7TOQ2FK7VQx5yefjsDF3+72KQD9C
86+1b4JF6W7XiEgAhr/XJ0LUQMULkOetAw3UTPQ/aiNocsdZGKqzNkHuxVdK3PJ6
GVTYTWJUorDmfS0MS7a8WZn4Le3NUVPKKqlKkBFHO76A0mGrwjisAJscfXz1Oud+
fkzBbcTOGLUcEL+wMvaq7FWxRvr/xB/Z3O7NZYXMXeGf2qJJaAtI1atbtGA1+Jmx
vRgXmvbjpwhqQkZQjOqX4njd7sm1Jl0Eh+NXtfKxoShUdjTizp02/r8vmL4qivas
gzR/GUVoy1lSGo0+Koke7P2eT7+wiS+TRfk0CCDsvZpSp22cZ0Y61cx8LuMXyvmg
ox4518nvkvRpiUk+Yi5htAGKDePWbMfZ7ezK2SyRcyLq2DRRa9JJPvuJZqefYR2B
JHTBfSjUmGaEOXXNUL76U1/fcYVJc2T9LbqmDFyNRUjBj5rlmOkxQ07wc8FNRqYw
AvGlYNm94iYrKKi2hwI9L3EQJpPWfn6SS5XrogHUlEE5iq/DAShmJr/XqYZ+0Zjq
5lxaNb9cubYsUepgWax2OWxXpQ4IMxzUEkTR1Z6GWtQ9j/cw1cB0NVXi/ERkyRFw
FVCWGtps2k8RGKE3gD+ibxhYxBQcYhkMEVy7NVyQd1CVbjmvU5xLCtMcCEBQZpUr
n/FLq2AlxmyLVsU3GJQjG9K1O2Wk8Vv+RXwUo2bDCFja7ID3c+JQrlaRRHuCkTyW
d4PrdpGMuWmESthX4EhXmz+CT45xYnu4/yoIyqHJ6i/NFuch6+VS2im+3+0IjMU+
uc13NANsslo9T6MVW0P3u4Ry1bmq8wHwwfJk66zZX7sIsxCPm46VGVSY5B2UriOr
bmRTcjNognyZ5KNINAd6o16tHnOItXqvBnKnSJlRvqhCciU+xcOhWX9/Y+hhRZQf
fdS1iXj91XIg7my+jAjiogMzO7mEPLu1dBFay67u4lRHzaMQLNH2aB4pZO6v17HH
MmiPwkVwxMNDeaUyXDLtvs1fUT8t/XqIThMpDvQgib98nmhHQIEWUhAy6rvaxNca
bZN4J9lRWvXyToKvlj5A4x1uzY74BZ/NiCQIwuKcLUsKkCT3E4q6Dcxp5yGwtzgz
G6wjOfDs9Km3kYPhb3DUX3BanVQnRyizo34AOIzbmPb9VbrLSuUw4WOitxKBGzMr
0Rqw8EwOQedRNLtVIHJg7qLVclFoTUjnGUDumODGhHdkFAD8LWuQLs2A0fgWPuAG
8gN7KCeslzYw4Ct2BpAXQ96FHYSZlVzRQx0B4VwmAoXfIfcCpHlj9Fr8fc7rLelg
iXApkAh2qM+JRP9Qv70QGVP6mKGKGY8COiBNVck9/zoJ6v2a4zv08Vl7ZZ2jofyX
XNhoqm2yHjPXNc0lEpEJxpQJuPfUCqWWkxfj25ZagLzi7HhfK1t50AYpVUedwgha
Rg6pffGB+SkTRv259ruIeX+q3xRi9jAivwbZ4G+3JLp8qdbAgbB9qSakHbPAqmZP
dnKNpP2FQt/R/4a7clYGB6Ep6tZqkozDSeWP9q2pkTOuo7vYgDMXPCV2/a1vrOyr
XXCZVZNkqiHLGinmtbK6OXlHJoj/jlVbsrTHfbiTHWpVGZEyHd08cGSA1FDykLgQ
rUlflxignyH/PLv3x4q3IGuK5e1av21KesneslTM24lInY4OV70Bm418TjzkF/I8
1Gqr0DzmoXWCIQ4C4D5VU3JPQHT7fRf+xwKAvuF/AIpW+wLAes4bycGOGe1wJiu7
vk+PvjK56jIJoWZGB2AGWVV3wuE6R7ze6Hg12pppR1xgHVOpenmnOIujJ3XBiX5t
LZaVEAR/8qsVwD/fd80jEmXB6CZnKnR9vY7g2WiVIZ8GGKiTnBkASiLvFI56k+ge
rwesQP3x7yywK/rFA2p612mTUhycoXICP4d7IpyccdPye/JoUxfcavPcob60mLcs
g+fUd+HMWVpB5lWMWkrAvNdLAIaCzI+wnGRAzHTWcEvfx8Te1seMh0hj1K6kmvYQ
fjGzGA5bsnO9ebAAvowaeJlEEgjgtsZWtp/5mbNCIXF2KEjizi/1Y7NBdI2HGiGb
JfflqrkPMFsMdawwTO1jufRXfupXcEjNStvjyZVgJGB4oMQA9XygiIHIBQjCqSbP
t58cWcMQWJwlays47I83BJSv0RGMGvWIMD1xTYOMHK9gCAaPjS8CGhHzKWOPDO+F
yE39HKUnzlweRZ+Nc5FCpUiTufv4+hNsvIHnWgmDb2IV09fcKW+d7jaetr9w4Eu7
lPQTY/AllsGqucDx31OjYq4DD/2S3o0BmsmjGX0BYonngaHJCTIYMhLqBROtzciO
4+IhFDOBvdL9mtPQg2wzfV7wr1oGccINeCS0cnx373o5IwPOtzFpe0fJLwt0Msv7
PA5HSUagQlZHBqnW9sKmfKH82fPhlAzVrUyhYcY2UVq9bRhuE1hnjgtgO1je4rtH
3UZ3xkKxIcOiqvxwZDuZtViG+XHFxnqUtSg5LzGN80S0+TQr+gTeiRiJrpOOPOeQ
HYUAWUcFDAlDv+6Qi+CB1p6CGEQv3ZgbQiBr0nSs7BA1qzRdfuHUXcxAXeVnCULw
tz00El9ng/GKPzs9fynmCRhPl8xVnX69TT+XNoXPymD1cgWEajzZM6M52ePozmD1
3zzEvpCeX4xx3lywFFoZXi6jUjsTTq3B82ZhER8e9bsYU5fgYG2tAK5lAG0CMYib
8V8s5c6bwLwush4VFAJIQa7ZRaEP2JUz9Nv89uZtFpi6hoQ1hdBd/N87YYS6y8Xz
Cq08iKS2k/dsJEABu3dpkq7Iy8t3GrLoA/tnmGo0nn4KnzNc99Rv39riD9HwbUnR
HlmFK9+ZXrRXpWa8xAVLaruMdv0UxmUNoW86Mg/d5nXf+rbRNds5qkVFq/Gig1L1
+7TqWrbIqU6+6tYlqcCu/0fDF0+1MqJxj7wC+10FLrGdHaKyjC1woiip350hNhXQ
+Zs/CK8JDEc9Oz8Ed0xLrlR/UN+0zBwxU9svCicKUyiyv+f4If8/zQ8vaTmwZunO
L1wGZUoKpoI7RSAS8mfkjQEIXXZ+P8Q+gx7cFj0lFoy2zCNvaoQeusGwjUGgfVO6
WtVKyB62xDwf2s898y41E/nN0LrJCnXXLUqqjFpUzzLcMPzK+uA7YCSKKck9r3NV
8Ek+FkZm+QJOh0LUe66ZjnSGjTRjGRn9P7AQZYMu1cf2r2rVFrvXKreVGsHY0tDu
/TbE4U/L7Dlay07m/MJT6erTWKPna4aXlr9yLm3zoRgjcSUQ6+Y2xiG0lan7fFuf
qjPkxKyO5nqYV8OA8bEaTlSLPUthaXhB9ft9lQu/VoXkBM5UIfGXuvBYjcdVyKM5
EFBFWcaTdguiJJ92bTx2puXHL9sXzW0kj/UuyFREkvZ+wR4uwD1OlzZSG5MBaxBT
wGh9vEB5LyoiUf5/wQzaoHJ9poEM3u9PTLDIf3L435UJQR1P0VNlq4nXcXEFJY/t
Yce9QPobq1ZJ6CGIyHp2EPsi3ORpGAeXaW83QHPfN6igKtmHgRdvfmBpMc0w8cz6
0H6QYesJhss5YhHUQ5fei8jB8AyQa2NLJ9G5A2Ndq0t1nizz/GdsTVKVD+1frHc5
rTgw3OWY2FnTb4ZmSE+/FbCbE/2/eki1QK2h90PBy+Pmt+7Ewdb0Atq6uKyEuDnK
cHUKr6bkEkL/XCuYADZVT8UpmHFWjl08dqR94CuxFCBfOkmsQd+6nKhLr9HlGuJv
Cm42tN5D7ZSp5oFABqvlxzM+ePxbTtWWCZUNQeTjREsdX5Kc1shuZ5NKpn36cHVn
9EQ2xNuKEA6WC/2HANFc3fpgcEdD39lTG/JvK/GrpIDnhxV9khF6Zd9lddtIsJYN
wJFG+6XxlO7JGu7VC3mPY70tkubrvGG5r6qrH87fAWRU8+IMBJtzma06nzLoIita
EmwAvHaXKkOOjE5v66nFJpCzyjUqnQ1xuUldfnfB/EmmSmnAz+rNpDI77pdnNwt3
HSE0qo7XycJMmQ7wwMvDb9HPtSMfXQDYL1IVXi3LJGZZEGr2ptTeDVk9dEZ7lzrC
L+f7SM+93zOE6omTZ5dfatE3QbPySWYBzileM4S31/J9PVQqBKOKnvC9RQxejVz2
VGsBvQViJ5aBocl7jljGrfswqunzNsu5Hd9AxOt0YwpCtJFYpV8fdGbvkTiMZp1b
L4DxhuAnZpCL17tPLhvHgHElLiunqFIyZ6NU3hyIhGQOxMHSUL3m2BisE33WcasS
XgepdjWug2afFxoHznyPiFnS4mdAsHyVwR1fTNQ3TFMeUHy70dTE2HVoYwor1l8/
FXT3FGe6qrOC6y7VsOsrmTTMrNPNoTwteixhdcuMPHfGZ1ig29JoavAHrfMxFxup
ULuY5LyehTqYhYmatoD+FlMZzcw+BRc0uEYU3jzIjseQ4atDvQZFOD46/+FgyCgK
n3KfnTxFziCieAYS7oPEw3h1xpoqPCpvms3ouZkapPD0U+olNZTgy2tnc28zlPZb
P/27WPqGqKPaq6JniKyY5kIL84FgX4r+KqyruPWm3Ih8lqacuh/7eaw6j1AhFAGg
M7zi9mGFN4NQ0usOPlfEIuXigDNZgYNmF5IL2hX8umS9LvxzE5iDA64mEtYn73xy
22qa3Gm55WxTPUpKqXvvgRoQuNFpm7bDQ/A3H7+psLOHBa7lBAszWpbJ7zAwScZn
uAaDuY9ljYaNBgAS+bmQ0IWABYPDj4pgr7gq/EddOBhY6iyDekgbnfac0TEyCwRP
xL9W3Y1jS6GoJP8pkV4Ie2S4CQcnpAu8z2dBWBNyVQ4V8EiuzZYds9BLl0+kA5zm
cp3F4UkW3P2ZthS0Y/D9GTLBM/1Ivu6ZvyR2acHYWov1VpJU6IQMi5KvFOuGOWSz
41TKdW0hT6xa4IS7Vz9yiG9QNmOpMkQHDojRE+CZqVVGVo49pjXDij6GCUd/20+b
7QVyR7rmaHToYvWsvgCnW1ogJc8sMR2crdh9Og8dKi7D2AHSKhRosEWNBFYpRXhW
DCYRkhVdyEbcOIU8AKIZNuk6U4suofH3BgakbtynM5CGG6O3IQrGtuRvQSOSPIaX
gZ6p4NVvclXE/xxgyXGaVWkdObNEtdwHcqW836laExBK8ya1Ykk5sl1OL7TSo5LI
2ckXyeVp8lIN+N8grqtp6KiBJJ+NGkPcSAOSVo5L3ulWBZudaILKL5p1YqkyLMDr
6tEmL8Io0xg70Imo7ZRhpZ9BgdoZ3hjw0gZsbsf4abCAhXMuOojptmrN9kmasLA4
FC7NZA7qbccbAuPkNkv4//Hgq/s7oSBkMHG3TWjovyZrwIkuLHyC7AvXeoge/4ic
Uh9ZpvZ3PSD+jZ9iNKn52Rdi9sDt0+WlnRBGVujaXNyL+jVfyWb8NOtTr0PDz9UT
X9qXG+oFCRbSquVIavxJMTBFsAek6WJuHU65WzmYPxwIl9jugMH4RhAud77JO8/m
lENjdTpPKNUP0EC7lsiWV8MsBw3R/4yvRct9DvUO4PRQPu3SESVC5Cl0pdbhg9U/
aBLaSFKD0ppEKi8Yi1/5N7xBv/FhwL5tjfMc/z3VNR5RmMREfy52kG82f/5SbHfl
NI0MDJPiqFXH53oQ5t7qcrTEOvdLwjgjrlkMpAwWwjAGsVYJLJzfCi3uB2IoZz9N
el/MH0zRQVbs6kPe9wjGHei145sAEKkceCk1MFQ6CaSZeiYWC+D1dgVtSR8iMzbg
Qt61ZH9PO+90JP72m5raacYebWG9LvuR2VOai9fF5Z1Bkk4CQnzRp0i+0b3i71sg
SM3RShDVWZIhBTed5dZm0MpU1QsjoMPzpYqPnbY0Z8CzUAV0fVbIbdgNGDd63F3h
PCyHtv/SOZAtQ5qKvJ5xLieyrgcDVHe9LZZHUDfqxVx+95F3MQRfoov+zi2cjdQc
9rfFzWnoxB2EzSU39JJA1FtmU52i8xlbgH7i3+KLj7s0p3JM+FrvIQiNIa/CGnvj
W+OVp8E1PAUGPsaJfWjvi/VrekC5WWxaKJXkBUrC0HVHtaboQbLN0s8/g2WVI9WQ
mPnUdrofd18Q46r3I/GPcUmUA5EFBU2aJwDhvtB2tfebMrvDOGdDQJTnEpvM2DXe
JCt+iZNaW+ABrw9/u/JMzqT7lY+Mn6l4OrfTGFwehWsgMUmvahoBg7f0EUmnhabr
PCl6iS4hGvNmHuYp15xQlhmwi9ggSArK46L4Z9IwiEYXtNFFwEdpHjNeU8Vp+eWU
0+nTIDom+B1sKpH66o+U45kqHWCeTDAMh9Uyee0qEE4rWtqhEQTmgC4ZbbIZz9Ta
VhksqVOMT35rrfkO1IE1Yv0oGZPvwpRgH0gLnq1fSBkCgfSYHlNt7Y9+b9xYHaxT
rUrFZvj7b/haP2DoupAoR2smVq4vzY6KtOXZvtcjEHNFSOEpAZW8onDxfeaPs3RE
IHnM9aD7tAuRszmA4XLDC7OoBd2mCcuHt7DSnK6HiRhBSIztmoxrq8VV1tDwxnSh
Ps2qaZh+c0B6wU+/nc0mgvs1NOrvbpeO3s+4HxefEv+MulMgtk2xzvLCWxtV/GXf
IddZbR94y8SL7L4rPL5omJNP5gyhhHaCuEXczpzf+/Ly/l00tDRrqHAX64HR+yJo
pCu4pXthqn9opZ2yJXAmcz0G9rQdtW3livyCnS0XGxBZCgXqFqaUQMuqVdv5UPf1
T3f4NOYCPKOwGKTGYObXBGULsYMgzOhB0qR6zyy9XHNYmOt7ijXJ0OxXcy0efUkU
0QHfy2g9XnTsMVdqXY1O1v4i6Dqh1iwQvbY0uM3cFfhVie+nGe1hlXPlKVeaqF/9
3UcWbLBR0/Ys9jHl6HhLLC/CsjYhcCqJTlMzAArgj9uFyjRiXNycNGqlFa6wlvaq
RL7GZoKCVcghnK9xXs5ZO1/fX0fRjyDqQNpgKFlMmYbauW9+R4A076c6ywVyxT37
du6nCnehOkexUBLsh/P18U4FGgccJvI08FHmlXqNXtJxSIljjL+n/iBfBaE3Tp/G
gduznAUIw2sO5qVhe9q0TeBVEgqE76xsx62L+Dfbxjdg19ou/h8jTwAp9jX+Ncj2
H1kgByxpvLB/7E6RhsLTZ6qJHw2f1LUPFlMyb1G32eiI5/OL4xLfjbI9NiYBQz/9
18e/gKDp8dCMwceqFdoyxUPy+hyC9LXJZi6400Z+qYgT/MZIYO8qWtwJ3XHE3psL
c0dRg361te1kQgGRSfajyOpVT/yLg/ZibOXyemVnPLs5KTDd5RX069SxNt0a4wFb
yu4j0Ck24MsFWLBjXxOdqm939nBufhvuf3XLv/z7AH5Az+W7F3VUWBC+MFGtp2SM
4Z3dfJjZ07ptKpXAs2ryXlE84Mg46t8zVSvXot/NUCSTY2dBOaOUa8fPx2LSLnaI
2AZH90TvDUMpZLnPL1MDELl8c8ZovsecSYMbsNPvl10y+Ox/MDTw0l+aSltWFu0O
Hi01QoxSK3toPK773kNtUMpulDAcGpNSzr+RAzW6igfr7+OiJ58rOkZbJiSBls7b
gS3xVuRch5IUJlpUN7NH+p3X3bloMj9gYw9UXERPpMNxTTiUbPQwME+SrLSeDEpy
NeHRAJ3gnnTtG43lwTYUj31LZuiTtx3ienxT41uOFQigXQsCJce/oN1nitXrh5kz
VIanivrf8IyiYisXFsovCCRiXW84NApAsD2ls6k9W4JtbRnDU354bUKYskBFmIAJ
HX1UrCW9IZJ0GuYvmmEUa0ouDItNXCoWy71gPxk+Hefn0/O19uXkDAsr16TOcNkV
qE0Y4EAxvIKzLL0YOwI/Yv2jmcJoz34oI487gbbWZKiV4n83vYvhAGVwM/RyUGlY
RCIcDalaAQFRKE4UVjCO8Cq9UXZjc6luOcakAl1CPSdul2AaTaEZV9sXU9woXPcv
kHW87lDXAF5Z7Sdn7NcJMSimhSVg6SU9Z33zaWtPguV+2nGma1nyKEsVfOtKRhT3
uakOJ0GT6sqJGGn6TSeinFgETiO7HPwLXhW23RkRceLO6YXAGy08k8MZHtzEgeUY
pg4lLi1YzSie5tP3ys7BpNQtsP+0kFRZ3BdDhsdzhHQvX+Snad8qVpmo2GDyI2i5
T0ZV5Vs9cziC3npcniJ78xgnTIhmsDIMbjCAlTgqzD6i+wQdBlEGEgCL4CXaBjOn
Ve4y9KNDhUs5ZiaJyMA5H1+71VfIJHl9EFozfsVyCI7V++0Mr0d3/MDct4F6dSEP
RqL3p78qqHbUL5YzAk/S8QdZ6Jm2kWrj0Ap4D0YXdCV0DitAetlyy0xsRjdhVR5+
L3eMh9bj8wk7QCpjy1EAtJiSV0RrDSsWGBJttFfGKgwfPoe6utaZ320dq0z/3yZV
wrVxphsMrMRzrm2ERLI7Fq/Oq6eg28gCX4Q6mZh54eGDMLDaxndGzGf9ZsfNJQNk
yHs9pSZ/BeEIQVJXqB9ISSS/WCCPlukTu+jh7dsZXbf9ljaTc6nxvy2+0rOckMAc
pHsXJ559rq+rb2YUy/Sno4Oe2RDHgDQ09RJJdlLi8hMoCSNnh7RgvM8yS5gpVMNk
HH+S1vsyXC7svWro19BHk8SOw21RcvlSzMJghLmfBWn0U8dbo6c/L8i2vOyqF7Ot
2aor0p2UcX9qwTYm3h83o1anCMoEX5Hz0He0lyCaE7hhoLsD4ZVuXfI9aHn0gFCj
mpjeM8zEubF4pcDn+GeN1GAJEcaALPKdP4OCakhX93Z5mUsKBnr/7LoFnrG0mCAx
7o6FazI4rsswn0wMnzgt76dhrRvmgsY+MmLnH9dxAVt1SToQpLEKiM8JwaneArxG
FpBGWhmMYLlODc+a9cdOWZyLQVTelvZomx+0KV6TIDPoE0KhJ3e1B4YEPjvdzrmS
TeBtZQse7eq3HmwKyZPg3n6qW7mN1LFm4+AckF4hLEpcoH1/+LXpnIR2fW3jkocB
j8UuqFNH2GryV73AdkmZWy3cpo3Ytv7fl3HDi/dzm2XYFXR6pyqswlTvJeE5iJDB
gmjMkWFqkk4BY16dJB9KFT3b4lFwKMLIL0/k/MGtiKjJY6PPQQ2Ytw9NX5yUAAy1
5BMfjeHFBxnpdWiVYktF85mQxboE1RYrGTefgHtIJ6nCitQLNR2xVicuGYWdCQ39
0LDO8QWXRaXUM9rMmCZNjy0RDNVBagjCInlAi2itVt8uIH/Dj3akiMSwkhNn6hSQ
D9pdZ86Ut945XGXAtK1+oPjvU1nQ8H2rgoOGN5qqZHuHns6NJe++cLyfWA/xuZKf
1/Dt+f/u+pkfBLFzyoBshZMKaxLy2uLjnc3kXVIWDxS6qvB7BQ4U1bYP/fIXbDmM
GEKaLWsQZCCcnKOuD8xv8Wvu9tbRx64O32A4YSg3UpkyJO4jBaRxsLXkRhdoqA2g
5uUx7XjnFIN1NDC7DWNPrB72U+RHggaYlpw1BByTffOVVCJWGr/fRluPzRN4g6CH
R09OEeR8RdRG118OVidO9yB3vTIhwrljPeyZ/1/DHTc3EHKv2lQD5crTxzB80HmX
IfK4Y4dJFKm2nFH1ExSulNx1WmYDzQc22e6kCEEAZXMeOV+pq8JwnCkhZbCt3kTW
/Kdc0zBciHzvghh3HpJyfCAzd2bARBTkkTeZ7U0rMKhBBXyYh6EWmbFBHyoDcgqd
3q9CABzVJt12TpdMRorKsIADYPS6101SUnPWgnh1UKFXPIO4v0T4yV8W/R5rZWhU
hHX3mMq0xMK2y5DPrsvBtkp7zXAweQnC+I+QJBRBV45VEHCmdO3+epzGxCRKXGaK
YJS/7s5+9u8jaw6p8knPI0ToLtbCUKlTeJQAnmP2giY1d6mne393G7ebmFAgeanc
I6BKIybzlL0rlmJaImhnJWIo8Vzbu1fhrN8vluSXhNMgqpV02O1d/4mT/YjebYKN
4KBVHJppXMHdhuem/O0jKwNUOqCf8mc/vOP6zagZSgKM7zfK5tzjS9kOXN1Jj2CY
wRjtcewmZgseVipl7fcsBz08LbqOp+yQHkgENCa3C+7+AjRoQlKb/fJKxXDNo+5i
Kx3pcb7b7JcBT5trxr9CaiNTxM6eL2n+bJv0HM3i8NZge41b8hgfLWT0sSSp1a1E
x4fNDbgSdW2uYDKwEmKKHyLVYr3545yd+xkoMAqIhCD83GJfFYQ9NA0eedlpF2my
1b/XoeFml8nrEAVhx0tq+iXofFp0cgh2QUEfrVl6kfzM7rbxo1fgBSZtt/YNWRgk
sEjEDk0h78IKKtMsp0GXeqRcst7ZjE15j2drgo35HCFx95DCPa/9jSot5Y/ijvbO
IoUdLGGZWDbywWKv6CNDxGJDGsxIdopknkrQ++X14vicZInWb1to+riyf4PnWlqP
EqCMTcyIMgn+ZTvzVeR7XQb2L/0bX8FJjQB9TBQsezktUJhq2FqB5DR8zDxNH4tI
CQd6eVBnuLXP7jl0D3iGaYb+Wj6pI88ZmU6VNRpB6FvlhFA/ATCj5j2s09wBRXct
hGKkEMX25VWP//HOIKSFbEB7+t5+1EE2Whe7rCfNB+BOf10gDmB0rx8xTtHqeBc1
eWsBmHLZDrevzU19C7WDCfJGwP3JzQ15xQkPmYaRzhciMQCo8/09d9oWBS8irzYB
ANHZM21H4ghwj7qV3Um78qFFwqcLTw8C1s37Sx9JUsHkbAbzrwcmL+qy7VEp19Yl
EIqDZxhTOEi9lPE246pS2THBwzFaX4BlAggiEmgwnqBX62vCKepM5lgHFftkxqSH
HedzzKHq61krjFOjbAcvvb7QHHhSFEXhjm9j4jaaTom0pKCRm3CAa10ILzICGHmH
sgfYFCLbLUf2NCQP9wS+PuPwEQIA/H+B+4KLhiFh78Yvs5jGQ9ErLzbbdJJYRPtq
mZ0zlr4AQ5jCh/rqjqKnyF6jvIZl5Vl6bekk+A/MwCqj0oMaIjQ7pRsdw1I7YarO
bWm2B/4xbOW/RCgbJDDrRkYHC4mgjlQwDYkil1EiRXhQO+odOvbBiGMd9SObSRp1
B23gTrN3qSt8RtI0x2fBKy0fXScWGDTYAvTq8G5QexFZYE7r1exvO92O4uowXYm0
AGDK/oFWOEHwyflrfnXpn0cU8V0TDvtJ+0nLHPSHqNyL/gq5Gs93pTHSMgirR+ow
cyMv2IW/5BV+a481SDU1OeK9ChcGl4ff6bUVmGHSqIELk7KD4ZIox5HtneDw63ls
kApBKrJz6WdbassxrE5L/G355eS21ypkn7/L48nGPFmu+HAz3c9FgdpGf/LpklYP
Fdc/F+zqXCRwxZHMlCAI/yRmlkh8TfjYODlyR871Vwuc6x4GQbRIxFJKr/RPo0vQ
iXN1U4FjiSCvrKooOJ7u9ZsgjedW9gh3obIpIXd8SefJixNV5hEeoJStxOxsAAoK
dxPOvwiJAHo2+bjgJcHP+x3aoZPOmrV1kyjQN+Kye9js4/f/IZHBnXK2EjnFojxY
9dfbVWkcxnKHpNlOoG6FEjVdAtSaHdJW/SrEHyO8m/Lp1XYButgxH6mO2gYksSJJ
fc8coOBJJWgDowv6/tMBcxIrAgwnW9DNhiS2bo1Ng/KsWhhqtLq2e5Ud6ivZoKpW
GzvENQo3ZvsNQ/q5huLxMb99TIEs0WisndcJvCIZGUUMPQu5TEpAZsl1cu6eKHVO
JvNjm8JPOW/dx6SkMb6TI6MpAkUa4zlpaXtSpJG+WsQDUXloAsFL5Eb6xMoi7OLO
iqYFJWu5GSTndsjAqd0w7fgYtk5wO+UyUw/x4DFY+FEF1ekvR/m9xiozWnAj6XWL
wY7AnU22usZf9PNcboGtiRFTtCDBeve6F9M9Ks4x/Yx0IhQ5HjRSddVYrmgBiv5B
yWbDn4bs1aEaEXEp3aVK1zH0bMEcDheXbPp3quZvESjvVJUYZARxhMENjIi2g3bR
ffoet0RlAGzf536kHOD4jnMKnntSM9BIRfFS/pdOOnYMDE7JNoaUgyQ4/SIdHdRk
CUEmTTWQzjY4jhlvUQ5oGlYBohEAEQnqlu+uwhAoD2JVCC7EHd7lrlxQx376lhAs
MBd6IpWuH2FN6O9GLfL5kTZYKOM3aXW7RtwGly5y+aWy3lOUxJDiYHgIH2YZSQPu
d9JgAdt5wlHI4Sd03h7HUqll64gu0sW2UFmB2H0wNo1JL94ooBrw9ghXdWEnoK93
5NpSHQZv7Mlx4zuOqgCU2HvuocC935C5x7cGIZTt9zS3vOTVcU3smrk7rcNi4muf
0E3b/OkKrrM8TjpowxVJQwqxgJ0ltEHFkqoQwKCn2WocDgJOapA3SRx7do/wJQFP
y9N5W2w9JBoNtDby3uZoYMD9rB1ja9ZxPZGRm0tXHFggDaZ/pkoYNWNAxU7/Mh9q
CFULsmgnStVO3CWiqe8MCyPuFrvETCVDB+2+D1YR/U3zKFEhTayKahyZ2zBDREua
FRAZzN+gtd6LtQbljn2T8d47BisjWjCYz4RWhbIjpilt0uH9GfZ9E0GMfPrSL21D
ss+9WCPSTLOJiVvLjkz3f1/mHSwddRhh3DAhR2u6V7Xhzbg/tv/1FzKvP2jRVn93
YBCaVUrvgstClktcZg/2siRio8P5gO+SS3/QgYfkBI2WSpGqMeTDOl9vjuH4Xzps
GJCfCHlnp9Jpr0rL0b8P0DKslRk6EdiH8PSLZdNfl1kgN5lgUzinwRTWyzZmFhEQ
js6CeBkYkJpLtAjv5pJldLeuoBBCYelb20BBDJZfOCWq146k35dkLVDRrHSaclgN
d5CraML/xK0VK91Uuig3V32Oj/lNb5twpq9YfWZahW04pN24RasQ4bXKVJJpwQPY
AbVmduhF5FmOgCi1tkuebzLLEb0HyBZxCT9rlbuxkXp9taRxsi1qtlEqA8ut3C+a
11pgBvG3cpt9pVil290rxi49+Q1IzDRUYwBBLP/qPvE2spMOlbFKNtODh5Kwu6R+
kWBE6C2vHD1nlGAae3w6L87B4ikIIYKq5ahjlgkgmEG+Eocj713L7ErybxGXKfpa
+TB3bgwjKccqSaT1MhTrz7os5cOR2JOH0wi/mfSCg3UQuFjrO81r6UMQPVxGUOLL
y613H0OV/XBJs5WIAF5hpatigP5xVpxi7GjVTc2rOOT24uTYqvj6iUWzVpzIWiMw
hwe3hHltoWyTjVoGUgzMtlITv9I40TbmeO0e6YSHfXk3xIg/f98UUl9qZrFzAGNW
aju7nPvIaWg7ez3EOdODJMNlatSZGMRdeN/BpTQIyCE7zFKVl0fT9ycCd7owzabK
SgyoQcXJGHI83VyVzvJ6tZCDJFMiaaV1Eceq31tDJGSLt/aS70nfjssTNRN0IBeI
lUcTTGL69/TDZafNgmKEMmgj1f9cmMSjhtgiZqCoyk901SiTJHEG3Vj+Hv5IN+1a
4KOvAkaGwIFek4ekZoAcdDntNFafCHJx29Xg3qqWIjGHDml07RYae6ZNFNxT9XpV
rRCXZef2HuXejHVJLaUaaWzOOQFl25llEoMyfRH+ObJexZb+36kRL0V1xuTSzdtS
M087IEpmST0tESOArGmr83tUQ+OoJZRkmpbJBlX5motjoviy/Z3X2PHfLUJVDcRp
5yuv/P1TlrqbvDxmbV1a4q96/ZBJC5r2YiJfzVPRRWD5toDSNbHWM5IUH24HOzeJ
QTveH9NH/INvFWYj535boallzIQ9QZm26Rkl/AL4w6VsKuWaWEccZWMjlan9hnqV
lZYHeYL5plIqLiQtAC1VLkLZSvtDHp1F96iZlTT9IV80yESY2g3LGVaFCcZVn2y2
7cVv8r9EVCoUcmQA+Lgiap6QKDx+ZUiyDgl/gJgl27X9+Uu9jVuwNC/VI7iBeCiE
0H+a69Aijtt9mZEsrSFhGKaNC+YFd67DuZL3E2z4vMxFZTl9OcK6GfTxx5TkrAHr
tpS+6R4x6LN7DY6rdmLQXsJ9gtWNJ7v0Qjy/e2beoADOgvHv6lrMMhz3UdNjgxqF
HxmloiV4KS/mbUDR411/EXsfOwlyeie8xuWvoys3Ur5VTRUA0fkll5oIhrUTv7/Z
4Aa8saZgRzeEjbsfGc52cYwgMs6odjl3HU0KSlSWvdzJtBZ2OLet3oHB+dfMbeAE
3ams9WTy0uSGi3iJXuNHiU5Ko4sjaA7YNh+HAN9DM3G+UqGYi44NPVVxjf2cbY2u
K2/JaJtt4yLIb84vBgaKE1E+uzWsC+FG3W5Xkl97oqLmVTLNWbtIyJBuvj0cNwGd
TnmOzQ6NoGrzRder/mvZXlDWeIIME91WrMNLAPEH4J03QGGJIJ59nwCedXSLH5O5
yP1FUG/7wEIfx8kMIBM/cnK878oHG/MzrlkmyBn4keK7VIVpmkHquFhPwwnjGKYI
VGxntAP88ZNfRtSlhpJLo/0haQgsuuMtmZZsIEYcGV0Z5K8Y/CTsXcJ9OjniZIME
WPvzRC/w2WT6bHN6yJIvc8w0oHEDEs4fwBusnvjBvYZHL81lGD8tGu6PCubwdfJD
1NAOqdNsKjJs6yfG6FkYa5AsK35dDLMYpLwNb6iZXPz/R09ytGVYRsHzjvTR5sXH
vT8nGPrcZ7SZMcAvOTFW38O4uIVpW6RAhCtIUm5WY+AfptCuZs6fgMEb7dFc8U6q
+zI9XrJk2hBNueYunJCIDdmYYgLQk2QTbFWwVMrRyjGttTnGPGqpYzRfxLAzUNd9
Za3PxWbrR8NDh4uJhsh4HuyOZfl3yarjk403o7XFId6s/JyvFoc/Tp4im/+AWYgo
CFrJn+XaglYS87kZA5OyT3AEITlAmfXzOEhAiOq+dz8FBre3tYn6xgkGBqXxe2n1
GUvTkz44L0KvftHpkwrw6kGs0tWwp+cCsiPL3bOTP1Ha/PH99FWHDyAG8weTO6gE
7HJXs6MflJFcPsMQWGouHnasncmiW7vZQbJXnx6TaMDxeN8CkPUNztzbrzkfFvvY
v9aC/EADpBVaLBR1Fhp7jTwA9b1xVc6JQaR2SUcAbxRpOjhCfVPSvgSP06juxPlL
jEwLgmeOLMEAyZpHU2p9ECRpKozgW+OWPrReO3Xaa90xoDxUUOzVsTtCnZpZ9BTT
XJSLhJ9yVyFeSSUufn6JD37EVRGd0ktx7zTyNKKYMGQyF5L2Tw7YwfNbOFPFQp09
hahsYRuVOVoPtN+2MS35t+0kB2P48kKxf8XfuZYXP5ZiQpTlDXzzPAiEOEfoO7dd
ihgn9JUroKtrsbAV995xuKFvEwRg1qD9/opUWck2rdPAPc7F4dW9KTiM0nd+XDvH
izPdtiSI3NjqM4aIY1sOlYQR44llcSVP4wytetj0A4WeGj8wKTmmxsckHFjZhrAN
7XiHtCBSo8IU27mbxJGm4kpyO/1QXXOdzCP/9LuB1RgTPm+vGwxM1s93Y05smbwv
jlBXtwK6AouA0q6TDYwoIRijbYoRSvbO47aqYO6gGTHLTu4uS9FllVndDxLsn2ry
ulmwg1yU2P4SO5R/yXK07cD9jP1QYedqbjwPa0Ek2gnyHgGuEcNThZi2qUIefwld
A2i2fEv8OQ3rML6liCvBUdqt+Lorj/scNJEgQgj9TVDPg/aFGArg/cgW33tC6cst
mZtLVFl+Uy74/OM/IKqZ/WD5id6PdJ0ek/Xm2g9PJBtcX+NoemzxW1E5Cd10cahV
3Mfrt1gcOVdENvs4F/pawDaqwqGwUKnbGNqfIzckdhsAU+MwzGC26ARrmXp92OVL
CQA/xWdnXRfHtAAyEzABhw73zEPRiY43bfi/zpToO1hzMyAxjL/J3H9MBHobIRR6
hZTfOO7U1jAdviOxaC0JFS516m5iGuXS1jClhrrWZth1pxu6nWPF3H5zGb2nV3oh
rBiQOi2YK75jGQdJOH1P9C4Iul13HVtdCHgK6pWrybetlKUL0J4fXeiTaXKThvDE
Rl0g00pU/sKitZw2z1SUsU9GKIw4F0sbsTsMrPIsG42ue3BqgJ9IVBOZ4lhSyIsc
AiCfJIl3L/HD2Fi7rb1CCVgGaQEctOa5IR68+c+CpP31yEYaUe9CtrINoAywHLVq
yrs34Z03FJgUn7EWpMmdrVDbDTbYoVa2jHxhHGzbFyCB7TD5Lmi8h+hjVE8kzDoP
DRjmkCjiVszEtOmx/i3T1Wc6xEGei9wni4e6pszEXegh2fFI7SeJRjgwqdo79b9d
A4JKGAN0BeIvvpK21MFNyg55/r9olX9pRhyB0+KWva6DUouX81US1tSVUG56hB5u
i0yhUMEpj8DzWNd+h1OgaHjPOOVqtC4vClwcmxXMKSR1n8JayM7aE6kbY/LsHmn1
AD/gWZW1vT8wnSFOMNefjmRoFGGm76bhrAcjCQR0EfLLvckQwA/trZF6A7d1Fosi
XcDQxOfwPqEKuYo7kWgHdCUQSqDgqcdkLKRLQ7OYAuF236zMIvftzPHDL+Wabe85
5b+W0IRRT92++4j+c3D+2zdRVikENC/RQZltZ5KiKnv5V68GtR0uWDFJjg1Hwrgk
MlA77Im6JflGmjNSLA2XdJ/LLaOaXuM5KBTfVbxc2o5hDIWah6qbv1AW4dHkoy0q
QGRnYrjTJyxI/oq0a6xzEObHP96ED3XRQRFJCwdckOcyfrQqW3DfTMT7z87C4E6C
CpbwWRWthE9ZzUqbkkjakGmZSa3ZZzrxyUwbzne/qEYuZgt6NoicbTY6sANlQOjZ
q8N+EbKOAbuYGHh1elbh+/DJTJkAIauRM/+wGHHzj83AjLPWUYII0kagp6ono4mc
4w9mJXy9TrognIFFkW36x4n4xm1Dge8aoWl1TKfuEEze55wfAVt35b1eRdiI0/H2
RvTewLhWRvqEaDeF153yp3eHs3gLbO0zKcwBq2/IRCoOPvKnjrV5LetjsvZ64t6J
rZ2vooEnOPk4LPQv+9JXyA+oHKuJUS/LQrTXBbOyBCxg+tBuEAUZiyaTbXdnrWVe
Ds06jcU/299YKHAxTB3FNohTWM81YepNp4CSJEKjZjeHjGejlGO48gHZTpwvVL9o
rgFk230RPKYJY8TeWskidWCVq0d6aV9hx1UGqsa6ULqMAMGNqNP/D+45kvv7jU+m
ADNeWRlWbyMkMcE7DZr6zYD2QS98HN2Ml35PRUR1vEImuBesAtrHH/yqlYMnAtEB
ACFswMYXQqBlbGcNW44jijNvqZEoP/q+v3yI2TFIQSq5hWrAgX376Ov5UXv4rqM4
VCdu3dhfC8EHz9yjKXaHV4TRq0ayOTXjD32qy2ByiVEa9fTqGDe8yp+rgK/K1udD
0zP4qnSuPEvsGBL81W3jAOq4JtaCwNnRCoJIiRfncjV8MDcncdHkbJb0gEreNCLE
2k0/uZeQHCJlHid6UjIJFOuvPNnpVjaIRJw1+XnP/oXq75nn2/4jvyVAx186W3Tp
2FUNEsxj3ZjKIvoRUvNwnm4Dzq0j6DrBQwPvCUb0Viajk6CXynosXGmX6bhZLn/Y
dDrUDIpsXUYMCyR1twi2Gj3Y/Cb6qMMG+aMkCZILH2jUxAQEV5T9Kx9RaLTJ5Snh
yhfun6a3ysH5xuoRnI8UDAFU0hu6VhZAP5Z6YYS+0OFSDXosVKtuDR/eupBHhySP
A/99AioFbP/BTI4kFqmH8lY6KWHyKDrpRdmqttqhLM5nCLsO8llt/CVrdJkdLR1A
vM/bR6yyLhizS7Hqk9wjOd7av0QT7fNH9E1BPGP2SqMUe2nRrjWtiO8dVf9627Bi
6kQhoXEOq5I23JGZY9axkhMMvbJkO0JtGySAPk3fxsj1dG8U2sjRpXs8qJaeyAoT
gTZziquLPPl3Ttsd6w8+kPTg/APcbzwsNcjv2X+PKBeaBvuvSTfxd4MrG/xQdkSU
4/9cu1tJiu2tUswA5cO/ydIx/sacNE0sFYsAPn2zbs9HHF4Ycq2253Cr3FcvSusy
Xus03ML3vpv6IJpUK5IHTz2Z57Fd9cukCa9BwSNxo9i1l+XzFqg06UD7jFWNj3Dj
k1sHyQVm6xMavdNhD3G1Mk7jluM5kJiwGu7E1PAv7iIhSJOgLoQ1UtS5f+rFmalj
BLROobOw0r04J7QR6S4aCe/wQi+o1woK6CGJWW08DGxel21klHpVi0xQpWTh36T3
/01Bjj1ms4n+sj/NM8+NN8/tLNfDWjacESImoPmGfTuZ70IUBTB6zWBnZVgrw91o
3MadQW3bHLA6/BCuFwdQClj4S3seV1HE5MBWn3RYibha5JxP32A3BTz/NtDTR2yM
Uhn7AyGi9NpNzGXXzfVDSZ/+NuG3d2Ab5qsZSNPxpRE85l30HymQziFTwEdo1HyO
xR9ywpRFSCkJAp0MHZIBTUjNDyPojh6FeDlqU1aYjY9GupWZfyNsezgypaW/wyYt
+oB/4J3kkQu5dTBIu4vmcRXy9MKmgXwcKHFaADVyflPe7UR52B225ZJmmmdP+J76
X6kK0xM2twBM5V+Nsy09/gF+ROgSCy105CAm/vpgdHRir0VkRflqVYn6USpf5O4O
zWxhyZraVkAijcqrbvrn2Sa7MyNemFClLAYrYSV+zY4dymM+TkCgEi9r4oTWUDSU
RqE+wbhO/c9HQdjWFRZCZwDcdswb8Tw2Tem6e2VzSw3SSQuifeECwOWtaJ27Df69
rOHmmYucd31wvzx63ri5TMZk25hocakYN7VoKFq27CxU58sVwbCCNQB/IimRZPL6
jEbDVHabQCDqwt1oA8f2FwrpqZxnVprBYl95BsxoCsBUfDVsytP6NO887Plx+3Wq
2E8leeaLROqnDX8w0YEbCvFH0HdEYWw5QWOAEm6vTDflacpYlU2iY7dz7bK0hFkO
4C52IZrZ8Lcdgdta49Jga0z4jK0F8EYbURq3rhUAZoYJqBj+eQpFVwpFcc7Vyzd/
psGMGtQDCBCc9/jau0zntebX3qRPuPZzW4TIial1GXDvXL5sd+s+iXL6qPUgNDgd
BNM66nfrIVyf3KCHBTYP+MLlDZz0d/rGwIriQEiyDhtIoeelhjiWIBox38YWI4tM
cy1dWBH5Szi4f03Ee5gqGKRD+yfcanLWNJmPJ6VxngMv91YkY2NOO8P3yjZWP6Nc
Yb/CSQ5EwqV4YIupXqPs0vp1yD6ITYpH0mIxjEUhy1ALnvAMRlZXBw+VWGjH1X2M
7L4zlSuoflzXCHGO2SbVv7JoDGgYxm3OGzZCPlJqmERspWzGmq62Pzh7ySBIdCEx
q0Rq3PEy0Wtttw2/kO5OZ54/o5u46qHBqWljm9TUg4R/ur4wHtV5OH5cC60nEvnZ
TD3Dep7NubkObat06q3A7nwWBznxBg1HN5M6DkHG+A6rHo4hdQtqzyK8tmpj+Q6t
8P50B036Ub1GV0Oe4PJaTZHUA62/U6NbVNa6KmtJs6viZe9l+hmdObPvUsECLH6e
V+LSftGsgpcpzBI7pn56c/qd2P0M6WoKPxlA3NJBRL6QkJwKT2cZqLFa2+gfFn61
uC1le+8feuxD6uysxxi1kmiNXhT87bH9i90/96dXW4sVDPwMZBmkoJV7T2bJMj8s
JoUyligsvGoKf/9qa5Rd53w/9NwWl1rVBv9bYhbJBKYhp/872VQlJZbNIi0loSzv
h+21iovjWhwP1ErueSx4YiPBEe43XasoqWjhhOAk0klxpFfj9kYkvdKclJx3P9/K
l3+lRXvWr7fs3M/7tfdjj6ZlwxFbKW2seP1hi5LdKgRIsQ+dzmGwPdBWpS+Gltr5
rvlOd1ANCYBje+QyqwlkF6WeLohs3KVsqMPjCiUgaLUL8uSd1nl1/ajSl2WefhcP
qUP14XfLzhyghFLF46iBHfPKWmtGG75PFGjC2HMBRydD8URVTXrqgU0Tf/q4g0qq
EYzAv4R70/+d7SlNyju098vrNFdPjhTqvu0Any8a7a9O/joyBbBflhuCQKQP5hoO
0kUTE430USfm9Kf5jj1tbnl/0FuDFKASIfUK19Yz8g4mDij4vzsSxbYyHd+Dd4wk
v2pC/uA6tK1hke0nd54q1bbaSk1FhI0NlmXwZl1QFCs6cmVUUoEMqabUzCIyYEKX
M71o1NRsvBE1YL9I8hUtsx3ihc7tXd6QdEJ+xddQkB6pBcAqG8AVspwIybKoIDNU
3J5GHOBl+oGsL+vvXUlH72kLorCmxAiVugrqsWoF5/VXhtqOtRbgda5dx1cYSi5m
diFQQ2i8m9/gUvzomfPrQ5C8W38ol/KRKZvZfX+I+mnTc+VTR8bY8eWBYypH8SL5
sUE3OOceY7hahtUfzYT3mmjA4diYsl1Gu8TPo2y4+R29jVFPAbgZ/iOJONevSYRs
AlCYpIg9K7b+Ue6qhmhPypBXo/1ewbB259yOYPX7a78ONTTx1iBLt/KJx1AvWXm4
nzSlqiirbdb6eDePQ+snTIr5K5tLQVUK2URndaWKZYZeOrcSvgUJpUwB0J8elHkj
iev6nIGHQyazms0DLf9kurbBj2DGAqQqMbHbvekHyVCG4W4Bb86HcFMvYLxc3kQX
W70Ms0/cM0ffJZiTq+RnZl4BpGFmwNlXOQehQboV09IcxlANqtvVIeTTS0syjExz
9KzLFLFNd1Wnv76VbPjvOREqVeJ2m0H+7VfcsNqcaONVKz3QX7ACG56pDqvj05gs
BGJI3mu0nsVY9OVHFGyZVD9B4N486pVwPXOwoZK0R1InNIvIG3PLiH8JBtxgTIZc
IaN1EFj32W+EijGQkWDhpO+fsNkPCCJ42uK7Pu9WOmbsNjEvNMCcE5OScUvF/3Th
Snhy6/ClReedX6NIp3OWdomtbBr+5mCCssaiAdcqdsy8c/mwrwx8rf+1hZVJcoHO
EPHSdVXuxbSXFvX1tRE6xMP8Wk2V6CAdT/Tu92fWyDMHgJT2jHnC+ZsEuqbm1pFz
5WVHorVngNM/4XMo5Im7t7fF36YvGznxZ1TGMi0fTgHhF0gqmd9P33v3aeMnvZWz
8YsPASbbz3GZoD7Urs3gbpZD1WNIyNv06xEC3m1VpxMj5iNvI5CnOv6eCKWygf3J
ZeckdL8iqiUJzhqtK2NnQMwWZHVW83imMdKdPmkzYF2TThqg01wDdcJbWI25ngng
Zpyu2ecVCSRmoKzWIuKMBHTSn7xMRV6DLubWThUnptBUE1eJgtw/mLVqNGxlSDnY
4cZ69zULNia0LGtVeCFYQKAp2mE2sPM2klW0XzupF4Cgdjf6aO4hG3WodYCo0E1P
v2C5XxIvkueu6e5zO0XjN4kewnJupwtEVWdyKZzbOzglKxJPPgFACcgezdTaCD7y
5xsHdwb/5TBdqURCq335ZWEbbMcQOlZ4AY6MWUAsgWMpCYEI8pcDxk+pRsry/Rkt
MiEC7lxr7A0YOZ0CQ2Pr8kCwh8CLGxUyY+Zf0tiZCXd7YN6pOLz9S+dVFdpCXFoF
6ks28rhRyyGxd8wdpeBer/3/EdgT+RiBo5P5kCCK78ratGsXjsTbDWCre2E9m3d0
H07fKC6gOzd/X6HK6cFGSyCIzwkT6KzDImhN967SVPg0KDViQafC+7xPZ2nTw4A9
2PtFGLAFYUVI9/g4RADwgamAPRVtwhyzDyJrzbS7jtZatKFGLffy7baEBx2qgpSp
3/48PYgEDR3XShDxnJ/6ScrLrFJf5HkZK835lS907adzID6BG4rFgVwOKulGQfY5
cFKuVcqk6Tqx3/VSK4phEJcjf+wbLyCfrm/JXR7yXPbiNhldnWaOkE8yWfeJ/xbc
14F2N2QF2XUC4g0l5mop4xgntzxzMkJlxlIIB2Q6qdLf4Sp3Yy+zmjtHX2pAlAqm
qWFopPsnD5fHtvILk6cfnFcj/PZo9JUip2XtnMDCtg8iggP7M2qVhThk7Urraba8
m4XlgggwUUxEXq1NZHrzFFMlhUmQPOp+F3O668jdJFYxQDjgIN2zE8X8E2/lyRoQ
XxXlHNscuHygeUIBAaf42y9iOvW2ORlKsrNzoEl/JCn0A9KuppqaFI+WLd63rotX
ot1kpHvSFT1Y3be+Y4zHPqIb/YyOaM2ml45Iln/qRQ3cUDP8keUaIk3Sjf5HeedH
EwEAWbdoqaOLXmsKd0VxfNZ/KZW6XdFgsQmFdADQalcQ28dR+HCISWSKJzFYf9nA
2kSysfvhjeOnplcTAyBCfEMpDO8yutTjfkGHxqPi0mD/aWBvFINmh5pJgzwLzEyZ
/rFtW1mBRGr1MPoijhi/zcKWeAGCBtfgn6spPEkeRCUB/k9dywGS+5iM5gUft8Pa
8CDXuG5MKu9MNH+QLvEXQ6rbo/Diz3L44SMPtAG1SbIDAX/E/CWGxGYqx5FoYjyU
GLuqivFRnss738Jz3vGsZYxo9eMz+TuGhLTL983+yvnSqjzjbBsM1RyIZ0smjBcE
hkfgR/shDPe1uqJbPatRqm59+P6UXQgF9YJgapb8TjjJdBCoBfZmSnnKfAjkzdTh
C83LT9/9AG8zIi0DriNyaUbcqL/TVCcu+kulR74VLPGtRTL+HLFG+aK/5KppWOBh
mHp00QWVu7oRYJhRN+K3XlVQMkH6qTkFb8sIpPLU1Wfoh2Ut7eU/3VB62dOyXCWs
gzF8/q6IQ7bdhb5W7VUFx8jihYCjvIP5W6l0uGs05Rb2gKZMjB97hv8Ax/dAbx+m
FQfpJkMXkH3jeOhzBrKtWGI5yU1BaDPuLCafSAfPU95LrqCtvl5ufVuUiTcUQ5de
kXmy+rW20S0aNxAM4Qvtx6GA+DmdLzY8iy5meFyy0lHCdItIY+GHHzaB4OoZADt+
RZ0Nx3USZUj0WSR/ml7fmL46FZhl8FYJD62NgCQJcfr9fga6vaFTPwVW6xyfuWt8
JLiQZOplEj6BWNnEbj1ewbFyaXk4VXFUK2T9eFyv7tzGX2eX24KFdcWq+0e5IR8T
FtGk0bQEQqlxyPbU7SBAXfbx0l8P1gI7DeR5DfmA56u742uZp9j1qsNp6AbI3yXi
cBzgWemng4b5LqgWc67obDyFKK88nxD4Le3iaunYfSMu2xWhT/L0esiMBQNDYnbP
plB2J8BhyWgjj/4jFNly8OoB/0+GdoEs2zcZqusD8KVkQKD8phYJbQKJIgB4GJm8
E8YZuZ5JxkE/xU0tUwWz4RCH6ixMPRpOOP1mvwfSSkHNBDMPCrQEc/bLxu3AsAKz
z1VT19PCU8r4YK79yvRHsieTKE0hfMHvI1gYLRYQbk43iuMdEChhHmOGPXZQJCUP
nbITLCaGH1RNE4ndb70SL+fjNGS6lbqOc1u6uMWH0Q6OoEPXIgOdKb00KnPPKDGP
B+A+4PADBePiu9PUKHHQJy9UENnojzQajm494QCfj9Ol1O8fPFqeakJM+Ijddzf4
dSRG7BTAzWQ9cLHLYOhc86aElccGtMMi0PgtAkToIg+jDORRy6ahpAHq74o3g2pT
md4/S1GBDt4lql6M/nrjnaFwIY5566hzEGZxXpRwNZhpRdmcBkqmi+azYkPuC7L+
0tDkiKmXzfSoQStguHQ9L0aSihcX3sIWAvifWYUtOMduks+V2Rb7UrarVK3YnnAJ
/5XTcrFvngxifSglUcDpXLREzm86yUs99bhXSZabBbNoSJwS0yfO347xhBYdCP9/
L9GgAE25QKqs1J9vBw1S53xbmKGXUG/EUKnRMoJ24j/RS2MFeADu4y2t487E441z
GL9ws7XQ39NXq1TZmaY9GwWKhfu1ad3kaFtrdtw1GIUcJ4p8pZYWnegaofkyT45g
znDhm8s22JisPJfezIIQvMPIesaZBlyye3UIDOdmN62mJg0Uo02vJ6joNST+g8zp
XFk98xQtywsqXRw8IjiYlYUfIgqhd6a+kDarqU6WDFkZPO0KYXoqPjoAMOGMvinb
RuD5Kt6qbqhIvZGeGuQ/lah2PZr73OL2hSh3QJoF9mcx9jMalI52y0XeD+vSZRqJ
1c87nbUvqFoEaDhbcDhVy2j2CLvAavQNICFjN90QEHc728/w0fV4UG0cvjp5IxHu
qWJhIxccIxAmZqbM8s4ySY6sE/nA4fskcHnKDNS5YE92CMJwI1mJ53z62zl/9G3h
idVqmM2KI60bYlAH0oz07NRZGCfBsj3i0hxac7JhGspMo7+2GGfFeFvr2BeVNPwX
3JVBpFQZwdNYVTcj7cCgU2fOt2SYupGxU8P+tt6dxtXYR7fyVfdlcRqpgsOZZXH5
8akVRSJABw27UOdl3PG6J50igFgbi6Xf6sCM+w7AN5CWBoq1lIoNi85TO+oWSFwi
eWhd2FIlq/iwxBpqeAe2D+QLVoBb4MUrF8LI2YWGPlIXKhIjvLGzFSbGfm7G1XQs
1f1Y0eajyQhNa9IkJmgAF+nmG6GrSVTrSwMaYewlsmeoRE/FVXaI5binI59Km+9d
+Jp1XGB9EmxJo72a+FnVGo2xUp7NdjfGIXvtu8BiMTyRLyK8FINHOsExfGHanQdO
BVXtB+fLgvE5WeOA+LSTLOWJkMQuUVWo8iqHeGmKE7BBg8xhGhlTE4EK2h0JSKlX
/v77YpCbWnBTa0WzYMyoWaVGQfGZaXFdgC2RtifwKY67ljzWprLyLlmH7+Yd0WPR
a4P/JRvMx5njAdrl9ZAXOpgN2ToQ1qmRWCIJWcUXmsr9uY8OJoUDy7SBidk1prow
9alK6gXr9dRAlo+sAwFp5FTmeEcaS/QzG4o8AO7qiqTHB2lrETpihMTgTnIhsiZ7
n/PySNiIf6V3+0Hpq4Ie0dhQ03SPYevAyc+BkUcg06g+jpIBUntm4EsOkXZc73An
+UXcb0JiL6e6TKTUjWbsyyBl3lVokubmvc6PusLRNkvKMTKll6DrUHDFJb6/+B9t
N++ZNz5nmPgX/DJ8r4BbTLyOsWN6hEAlCrXWfmzuxWsRKW5DN9KofR2svBfqJtDh
Bfglno5AnA5CsuOi3E6i00HS2RjEedix8dDD1mYakH6LKiQK0hRUp1YPrb1aI+qA
gWvcba17h3Dxuno6rbTdMvuHdw5UTXcHvDpIMXuPY+cbDGDDJTk/Q5pQutzIGb8z
Hk7fv3oeo9qtb0f9EpVRye6qTynmjTGGWvgzyN/HilH6BaAXIxBCxmbcogH3Erzw
tKX/KQKkmYNeSNMmzVCRwOeLDw4pzzqn8t5DJY4UHt1GXF5vYerJURrXQZ16kOPk
J5tbEWsHmnxOT2azpj52A6d2ME78UOMrkTyuGr3eLK8qsjObw4mXHe/0Dalx6oxh
UDtNpeC0viYkKie9vWPTzCupdQ3JvKhNDsZY4LuMiX6Zq7PIdOVSfK4PB5onRG4c
h5FvL+G7EHQaHupmBAbav2ywIicrJ4d9+O89xG5Y3+/5XiY6WoqHXYLui9/5YWDc
9nOqIYuBIwDNqZ6E0ZRnj6qrAIRHB3j/RqEO8b6usf1QdHdadh9U5s5WVUqcFP76
xXGf3CvKftHa6JaipMQ//eTkYhkjh911wqTSB6hLmPCjrwBvqVlxl+Td+dFaEBYZ
22DRtcf3fLYmrVZK6T241XLKDWnzIgp1T2lASe7JRt9+KE2TkOVM7Qm/TzxWwHwl
MCmltQagxcyg4FBMqKzIfHCjwl1tG9aaCVcmKsMT3EckSgwAQH/xUEu8AtLba2r2
vxhr0uqorkXiLLFXTPHs/1jB3gdAG/7nJif8szKisAAs6e8Kp/pDEYhNNigpGVpP
632mfXZa0BJlfE6Ur0sdHxlrqoHtMJSV9Rn4AlIn5XEW/2lZCzlyS4O8CBnBoegK
+UW0tt2lwZJP2xiDUuaBFEpQornqeoLkdgLIyTWBXETDkBy7Vs0wCOq17sBJf5Sp
GzgnSmEzE2yatGJNbbWhI73Wc8Wq/pUM2ZkdTtdgS2JvFUi3eJDVCaFzLd74kEqS
CT2/9GeB51pdDPxnlUINFed/xZkfSug4KSmlExvZSC8G+bxAMVH2aLT3xDtl25WH
RhEXR81nX51auQexXFcOzln6LnbSEgD4yTik1k6c55JpxivD68bVJ57dlTaflDeI
pIJAZAoxECDa/yGN5VHzykDVhSfOS5EpiE4byCOJ8JkASaPn1fHXUCYVY6bv2ejK
VT6Y1GHPwEY5TVn/jmd9PlUZFYozNjKqzLlmXNnq1UAJNtb8HEyQolcqHafKNsMZ
CI/y7riuxQmUCWGalmdis7ONUtJ3E/X/AIviM8Vq2T0+98zH62bMW5oUm7e7Vt62
zL/Xw8iSSTftaO6w7b3TeDta8RMaudi4bXVZC0ZsHKtv5Pel1/gA39URm35uvko3
ZCdTPfYu+KmeS/gL9l+fpxrem7pbAI0O8Nv5zOg4mYRsSw+9a0l8DUalN/58MalX
mBfFg8Tw/NrFeje0WJAVj8KM2ttRbRweUXg7+DrzMagqbejaYyE6cvx3gwIQ+LrY
G03oQiU6HTF9jasUegr4jHte3zZU0frXwKdxTdQWMfMZo9sS6Pc3XZ4DjnkuYj9D
629/ajJh4BDPYNrJjrrc3ttpkZGPIKRBBV++PLUC9S6UTXHYHSWldKcdKBeoH+J5
Dv8XnfhpGdLcGalpYut+s7Q3N2SdAKsZJA0Jki2T8+bgEX7UDojPJp0HeaQXb7yP
/RMd5uxHi/334QZ7PMgS95oNOjhTF2tkjCwMTZyuraL7ahimIyZyxduadlMOqR79
70Du2YDXxA0qzyZZZfb6khXBt+wPPDqL0TmKyNGrkF264hN2RTIf6qIFfbmBwfH4
7guRFwnmxI/kRI0xdv25rEkn2EQuVfjqh6zQqbrTkWimdKhD12Mc7dcPNzzORyuf
BWVQy+ljChBgeQFiGCEB6GPB0N+TD24ksA/mcHsTnRD5eLZE5/UYMfgRXPlYGxYE
V4Ht73+MwRgX2xABQlZ04x3ZQ1q30yhIFQD9NhBpp1jbHwFew1qFq1f1yoWQwgd/
I04phL9VaVwy6TPeTc765NlZXepLc5RjNEZm3IkniZUzaV+pUtuBqDBGfptC41TS
OEfG5vQ1TSaouCdIQzyY0/QUagypODBrg+OrX804Es+IjDrihriha4icgTh/9yGx
eRoAU9JQKXO+T/3sp0WrYlNtduvGWgEyGIuc87s34YEcTmsFwkhthRqr4K6vp2fm
gYEscHOFa2/woKaH0W7GxQUEhZCJg5nGB2dpdIgdiwoeYHAvwGbtT3m1WjgSDNKH
/w0mw2rD7OpVcFrNs699vDYC1ihX6orUo6hLsEczVbxJEj6HUnZpcRYtmBlzXPKj
GTlVD780thQsWHJHU7wP8YB5okCm7uhkn3hKl26FPH8FlHEl6tniXEAinFUGVuC9
LNJ4a2t+XH/vkU/gGCVeBitbJFVC/xjOoNF3HwJgTjpr5ckG5BeAugVA4mvCWGnc
8M6YrgSfgsMlwSDI4LLm5bQDphcm3NQVTRI6l5FJxBzcSdb4Tu/GxYFShtSfIGKb
aH0K5EC19qPUcIyaL0IYVZe/pHvwHZckJK1wcZJ9ZPfp6A+ys2vtyzJfuB+euyqE
iVuVgaUaR5oW713dHQ+ZV64E4B0mLoRQAkRiOc66ts0dmvT8RqJdgsLndEg0btoI
X6Lf/4k7+mIQ7NxyoXcHj2lCcjPEtLoOkX9/oQeMhA+HlKX7TdYugJcVcrbiZ3DV
3IqtZ2ek+Xg/v12uacdrPghZZc/rstwZ9smJlg+TJbJS7z2bJxU1ycJg8PR3n1tI
OOTtu0azz4dkV5AS15ia5sfgL0NxhXnYqK2KkzsbQQShswS5D1ex//RtbKr0QNPt
vjc+w6G5rpFKBMOaEu5fg/t4+x9ZEApIxCyAcK18LtvIXsUOOF6uPkR4gsP5g2Eo
9z2zsRbgzrjMJSY9SS/+dGpGTowliqp3ORVxM6GKcRJFH2/Q+BAorm5YGF5CYhlp
XPPyRFLVJeD4lSpvQUvL+ys5Qs93xIk3N0V3yXsXmin3jXtN0IBA4g0ShflPqcFQ
ISKcNJgCuzHSs8LpSBI97gsG9u/+FsDnvCSHHRbcdxJp6gMWP+kHLa0HgVLcnOZZ
ZMbJ/47COE4Egt3qda3AFVbmS5EIlCdQq+khxWq5vwcRMdvrRc9yuuz6iOSt3CRq
r32KSC4Ke8iq7Utoj6wVlSjPl8QCzQ/UQWJU6fPu/0nE18YJvf2PIAEjSuRUxfek
JB+DqIOqP5eGpN2meQQLBtENayGq65GN0bLFPTaBJwTDnegSX43rWjUOY0+C+sAu
28oo2FrLPeU2bX02y7ZJKQ==
`protect end_protected