`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 1664 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/9huKRhRMtvnNqb3Z+UU7TahEoHV+T8U3P3ufru7l1O
3DlgtZzb9QxCbOjthp9+wDkjygH0eUfDrEl1ovhZG632XOeaXNBs9G2k1gnP1bWy
YGPCLxe7B+3ANlnwq8p812WVHkQvH+v1u1u/ozNvNiEPmssGWxIw1wuszhatuxwI
Ya7e6y27rTWRPWwc6AiSlwMQl7TmgLMRISys4ocNFdYfm8OxCUg39ja3lWFgQes4
r4ULvqDSYNfuJJcXY37Ul7qAnIOGA8yBLs5pg+cfXbQlUYmBPNhdz2Mn4JA8Z5iT
AAt8y/6sZrt9YCU2C4kSKXblz70XSW2Py5EFMSnuzOW2JL0MgDfF7nLmUO3fM66q
jU1IBzQgypjtYXYdWBSq3N0JgzkSSEYcbJ5Re/OwrRiBQ50HT4uSbtA/l82Tg6Gi
FULQoCXSFXmNKwLpFoZXY93lKnoCW9Km1X6hLwEENbtSn7jfJmFS1CRCfOpAthUE
z/PMH3eAw8WD+/spGh6XEQWFPKFCNkI0dBLXKGIa6FE/JvG1QCQ8DOi3HUcDz5rO
gWTn1HrYkUVlN3OPbtvTOaATN2wyfjMbEHrq66lfwKaEMRTSu4NhY/1aNjywxcxa
FP44tyJurmKKRIEwMWQvinH3HAjzjo8fDU4bnKWQaTBdcGg8PKdbb53fj8Xp/MJJ
UMWhnqbaRVYDZEycXqBU+5qXfIrpPzJpIfQiv/IBeC5g9N7Vb/7En37SXpEOizij
hYcgtrxBiomk592o1L+AJHLXnn2BoV3u12p2v3ZAOLotbPPaHAxa9GVy4fQEhm7z
JOPPZw+eo+z+MyCvAzZZ/DFbtub3tzKGj+kZSuOJ0o7FX7k8fx7rfdPuotelFfwl
+5zR8U4GAHSCCOXHbneCTdHT2c95IrhbhAtrPBvYqs2QQnGrZp7ACMgIJVuarCkt
aSHh9q+O7pmyScwbJeJ/WYmrVBCuLuPtWoQwiFzySq5ZSAPXBpy/LlfofKJJ2cS9
hCIMjAvmligRRK+8nfmmz7pLrfXd9odvlYCryX9v93bXP3Kb9i24I6YOil6fqzOM
YnGIcHd/m4A0YmOYyXoLg4rjwLpnnB00D1yTM8W4Hlou4UzoDgL5ikTnbsvgtQmP
U2vZBjLxqcAbWlEGpLfgoDx+TXfWkk78TadKvnrKlGkiu6eG8/PmGVNkq5jK8dbB
YbPcvQxMtIiNhwOoGSpXyCgJXPos+Vu21PqUcFCHoFFM7i/rXUIy7Hn7+hUdmWbf
ESl65pBVwuBL7HfpaHdQfhmCyI8RZMLHtqUO7C4yP6s2teXKDSySQ+l1hueJTWPP
LnbYFmPYLC3ix8UU5y3dub8RK3EKKUtqIf+bBTKQiL4LUCe9kWmo26GkF3Rp+ji9
6zKSJXE+JGQ8tEW3dbP7kXtQCop3Th3IEi8d1dN7JcQEdA4knzCFrxpdtoPN4cqa
uX6PiLXLEFi9DLsQ93g7FUiFJAnUQj9xIGoH7AznFfuODXfB//yoFI2UINIx2or5
dFiTJvuNlkIg+cJw9TURx+eLMcJHxobYEgVNpL76bGFHjeM3V4G9LU8Q+7mjZM+v
spZW2XIXjeyak1ZmnxVRfrJ52ntGrzuJIwkR8EPbpquYq3aB0k0E4qUczq1oI6B6
5gwzBlg1S7ph/V1JCPi6YOppAqKJUH1kRH4SeahSCI2Vsj9KWzAbZs0ILd0xnOPg
K3nfxOxFY6PrmIdatph7Xw9X6GV/yQ9lN0kRbON9n+nnkKRvEYqRvIAPZG9Pbwsl
52o4JTeXc3qD996EvwmbrVC7UCKvVHH6xQVBMNlaMPB5H2H2uLmyIjYQysCQjUHb
Buh0OjzYXE9+fnUNEBxV88ZFJfwBOe3e51EOzkFf69pkrcjKC6+8SGBjmE1cbWFW
Fyh0aN/xFyrQy0RQ92cuAGBQAA1KfbLxCQNSdYY/wE9FChlZLaIeMOTMKmKTbhRx
Itt7HRxcUz/G+hwy8l/JaFs89VAFriAHsUddyImbo29ZQeYnEO6zg5SP2tVUm5cn
gLYUFcvUGuk27w5q91Zrcs5IFXwqsfUVNHTOHkV1Fw9+Kym+mvjpcAGMoVUTFyve
syDWQHrHIZ0SoD1D35rd26896X6r74DMEZXoPKzFWAeLZ+PVuxYMzemG9wtCY1Vg
KIvGqpk23lvACAfliygsCbn+onv+z+HexkhEK1HQoJc=
`protect end_protected