`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 10656 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/9huKRhRMtvnNqb3Z+UU7TahEoHV+T8U3P3ufru7l1O
3DlgtZzb9QxCbOjthp9+wDkjygH0eUfDrEl1ovhZG61VSER8bz4z9vRoSvozvYaC
5vgpVtE/KEnPBf7cHX2czsmgc1ydvhgzZEMTF/RQXnzFV0kFJEyBQKhAHle3mE5z
YOo00cidzpxnBOo96w33UreOFgkPgBMGqklWL0YVHKgouwMF7MXKrMz9JFBzKeJ0
LsEZgpQosze3s7jxqDWSfezY0JIMM7hV1fmzVLS/jidbv1jf0JBIXRu6U6yPvjoL
eMU0CHF7ftTw3XwCe6m+kAcxnhSrChS5cKG8o3dc763vlg5Wqz/q6pF2BehpHe2B
zl2NAwB+L8e2jPlFIUDfVxu2Iv3QGSBU37F7n2r0vISP2fFO1Cn8kBTMZ/tL8nDO
IPx7b3Gb3auJ0Tgl3eun2PubWk7z8f5FuSvSrn/sTtvBdO7UVupeuQ3aiz1tg+mG
IDSEDs9vBEECFh/C06j3+JzjWUiIEkxkhUJkD0ZTTs36mv7b4KXZhie1aTTe4jon
8QEcduUVGBFN6DWg7EPHnx/+43zU1NVs+OH67wYakw2ViugfJuKVIIc39y2Q9fJ/
LlEnExe+SJnJsQe9iN9azLZOhGtj2cdy1KnVJrKwVba6McdgpELreLuUxqsfqk4y
d9Kcmlk0jxs4JXwmHWHMq7GjPrx06HyQGhi7HKp4TXdMMdyMWUtbyxr80rJuraHB
1BUOLSHyG/OqSnOjhF7rwEzCgszIr8Uhf4+K+7YqAMV7ygA8ct9Kx8rDyRcg3Kxl
047B5vZELs1iB+W1BGIjPbBS0JT6Ap2w1gA9opdEee8hhkaNmQz7szcCDxPhHIjZ
2kPTSpwT+D9qpfr1RftjZQxeiidONXnzfgb8FcMgPto8UcYwkn/hJ0DPaHweLszY
a7TJImMJ8w+SEjjRcPSvAA4KgZMRUJgkryvFPltQkqdvynMD+yEZkhB4J2I21vT9
WtnIVRL400hTnnIz+fywsgevZ1iLxuqZ49DCOWuhyfy51piOxvEOg+Wx1k1hu+2M
lwhjcAram9R92mDSAIjyJvpPgRR2/Ettz+ORBv2jj87r6wbLpzidvNnZJpiMtBeK
SNrgpJGMGWp43nhTymQvqlGmSoxOCeUpM1APJvA8xVUnaQVzYpjPVsuO4SLs9Khf
6ietMzUrAmg4rcSBVjGPEk3QehUOs5oIfjiRn1IVPRj372KP+g9MB6wv7aW2tCLC
McoUVaShajxYV/3JmSyW3MLHtnjoNDmSEug4BKrMZzl166V+wPM71hrdQZeq0kab
jCydrAS1BAAH7z/FXOu0gPrOR5KFxT2PWdBIb4TI0tWG2qZU3Ex7zYHC5sP2bmqH
9Lvyci0rSD8SmaQahLjBGo3s3zMB7ZPfRG9IlrlY5ruROp+VKt4zXlRXW/QJTvmG
CKmP+4PJkPsV5UbzmxaWKlPBlSd5R9czofh4ckccl8K2FHOZDHBLaAckKL7GPdKc
cJRjiU+0gwsEOv7ZMU5gM/x0osI6WutOZ1G2+1BdiB7jZ+ZSUWkYrtTK1BUGeFhd
UdCQoJ9vVD8kjENQ7RGcraCG8SSzRktl3GdMq3SCf6/+8j41YJnGGC4okzy15YKw
1EoxOKY+NC/Kcdyxw26ZpQX+cofX1zNH1SP1NV/O5ysOLv09p/r2tM1WVDH6cwP7
03nqEQ2qdLHtzs+3gpDkG/y3Qe4lOMbWky0f4s2U7CINEaqWPG899VlbT4zM6tAt
ZC7LYKHgEAbgfSbv7RzBZ/cWA4ZUZPVJR4tkuf6vI50UwvhzXHxC3XhLJVv3BTea
I+nTr4lzfesXCW42+7m0ue2zylQeGJ3lVCvBQmCrLd0L7pOwdWdNZ6Ve1jjUpjDg
ZHkrke0Yc8FcqCJxXp9jIiMcDFwe5fARqvVu/d4aUES3/WJqAzZPtpCdaF5CkErK
2ZJ3xZLZkGHIE6rouUYF2iokAyAZnfy1/8bK5o24mO0vEn5o0MKHBYrFvtQYMQn/
8I90PXeVf+QaTJGKbcyEsNyBiMnaJsI4WLrunEXCSAmnpkFHFtQn4lB0ZEG8nHVI
oFHcPc5nCMLDRN44wIk/KnkmJ3Oo9elRSdrpIWVz/xBGdGM69TTPOj4yPwGo8oZJ
anZ+qD8XBVRFyo2O7Qs5NcPpq1tNIHG/lk61jTNg+FOD79wUQA+6vFueTV+t+ALj
K5ksg77IsYdDXtkaT2JdIyBKV0wbhwhInZayqGCb38Kny82M0v9ly/bIkxYCor6H
q7YDTpW1FpXqOgcw82ZAahZ5konLG1YxekdcVQs8njyB8qipJMu5QCnJ+/Zzj2t/
EcHpBCgLschY/e/l78+S04arM/kEnGCMi/qmK9LV4gA1Xyi/cHQ5OGtayC28vzlC
c1g+eWMDI3CcilFNa6p1AidxTdjX4lp7IDoduC/IO6PZAgKPK2ULAYUeUVpkjhJo
yjiVgWHnBF26v0hX/YI4jRr8WizyULc6ufNtNYNwnS/UPfk40Y40+CR0vbGejrKn
DybwFKlvIMuOxbsMjXjAXMfbNt+SW+pOh+9LUpmL1x1JWUvOL22zQn8kFyrC9nLd
uDhDnRXiMv6TS+uhTRSigO+VZ+3gzxdgHAds821J6vsaH8v7MV4qIrGoXkYwodst
qF0sttrJaRIFOjDPFXGDDw2Gm8O/oO4mnS5nNjVAe/hkNVqOn2fJnr6HbTyQoeus
9kQTpqwuRs4e7DyeDkHOKQE7F7dIhnNWqTm7nYMe82EWYGlgSgcMkVV9NYxLFBhW
36/51Q5orfWQfCE3WGzlU5NIl0AM2+AZcYQzOoyKHT4Wjiqi2REjBRlVK7wPMV90
kxAUVDImCzCLaQ15T+Puw4TU4F66Jnun+tIKXy2BHhzxcT0e+B26ldZ9UVNl/xaC
QatZN9SSHjjPz20vlKIxhZeb4OWQVZGsuTcxcaiXB6F1oYexFEHn/ehmcnX36ZXx
ofkdzrP7cMqiHcGGYqTruATfDGyrxCpHNDZooJDbOOh+o9UEZa8H6eujrp7B4gRR
5wqO9lK6OenPAMSp3t5GU10RW1fpBWPcRO+ur2HSK0GswQnEkN3FQj2J/k5JpwiN
Uh4X/ABsSClK0/sokDW9vGI/q96sB9ODUOJ3UAZx5grrxSlKCrMzssnHH46ZnSKh
EhBqLVz99OXCi2ozXMhhOfnqFpuzplaVjIuyOzJRw39t6LnbyhV16iE53At2OlAu
niWVjj4o7ji6x4eL83vzRY78iTAZxQswoLhfNcpMyYA73XDc2XW08HYv32BdCv/c
9CkewLrUVAFNWI++7Do+6kSnQ0gceNylfufuGxgV9KRrD1N6Gwti0QbJFu+8FFic
8fBjCigUfXT9OC8IOllRioAZb/0oDHIQYHnOuSiqNB67cL1clTAP2b+m/UUidWAl
d3O1nQm7sd1KZHUld3aPupfO7/qe3Odp/ttcD9xTK5XlgQAUJSPOxOiaE1wsFVpC
oiHDHyo9Ajb+unL9kfqqKUNDnKevYWHNG+SpPOuJJL1irSNWnRYHPrlHFy0VCaP3
v7EbHgC0xXXiGwitp1SmxGX5rNyj4EK2S/IbJ6jkzWSQVqRiywzpmqvkc2aN8Fq7
3HkRuZlgoh46lNkkNVPt9lPBregVWihE+8257096dfW0WANEtyLcklvVVNqqauFA
zDpO+A6j2D6BObGNArJDWJJ5e7oQFEzk1uBUo4ODmzZTLnCHn8wprwNV3jp5tFnb
97sqD+L61MaB5xjXZPVQhuao2MjWNjUkN793814J8umGqm9w5hUlZ28oO2TyhEDZ
NqsYpYHxuE2UlNyMUcLxSYMilfISHCM291q0F/CgYmK9MgMRp78kQzkpwHr9kcCj
2znpqQbDlLy3aT5f+v9/X6MwGDMWRzyzHS0qf9ggkQuVs8gosSR2BrCOXkPM9yy6
Tcds+QRxHaYAYiDNVwWSWsgwiMbB9WiIF6Mle/EvjLBwuMQmLKRW/nQqde3smBfP
0L4KmMs2ggnmSYkIZM8Y69XStdKzTQ7S442q1nEac3nqQUsyr+RZqT6bLMa/E6hz
n4M1qON9W7t3GxPaMp2pYEg65Nr2ICIRusSqRdjlbRIzbRVYMHK3AQqoPf5rKSOr
vmYy17ACR1S0D1OpYmWvgE1sAuy1ynkwkQMBkbZ6yUxZW/0wy6duwu/RgfZzMJup
JYCdd+5Ua/fCQGx+dQg+NznjbwRWggfCGkk23sVzGX1I1oDABmSJameVN1wBFef2
d+NvL43LV6MyLZxxoEcriSOPBl+FV065/3/onXTUvzS+6OVjXq9pvzl5RbdOkqH5
WREOx84eiNORVS9jAq+BfZ48GeGZ7BUpKA6ets4tqdXknuew6CjauXuGO9LXSsbD
DI+z0pMGGzaO80ca/9J6S15kWenHTYtxZJceQ0aqcg6j2MIvNTSrSHQrdh0J7zGu
/2R1flVNn3Km1qriiC9FNJWErmn9t7irgf1xGAqfjw/obo9sDUiG5l+Mwu+/QR/4
jFCFgLkFq9Vz9gqdG6heHOdil1h4LoP00N4H3i5DLzMvl5n7yVWqzhno4pxuDlbY
zClGHb0SwvPzLrEuuDt+af/WHj7kGeIxuCYg58aQ82fm5iyggiBqGtnaV85swukH
2pP7z/gKZT68Rb/0ske6JQ1kcftEGulH3yMPxeTJ+BCKs/1Gj4XdQ+kPdRdfzTya
d2ubOAfK7yFE44/qrEKj5ux0JT49bbjyfSzGOBi2wB1if81fjI/CYFxPJg0e6M+R
rSCQWLlsgMpBUhMgpz8q2e2e/QcuvYtUboOllN/wfnsyg5K0yraGLZ0ovFXWcGSc
r33Bp+GdkYoxD5tev5tNb824qW+7g0zZCorwmVoaNyf8+fMP2JKZgke4DDGhqazh
66TXWT3LCyfFeydj40i/4aS4Jt2J+FZj2GpSvg09UD5D8gtaukF1NcuaR141y595
4POLblbU7DozyVHH8SXwlXUJsVyZni56ku+8GbrVaqz45Ii16cDIX5ghHc47GL8U
8PfKRRvxmGolwbPlFqlJpqRh534waDtES67Zx2tOE9GbPybSvnvgnxpKFpTPvE9w
fkSd39O8zJ9mZGimaB8L/3wgT3ib7gNSAj8gQNT1Ck9rRpzHoGaIglQcMOGbICo5
vjuPdaEUysovHWIiIh1m1SL1dZP9rUbYJxJ3OulLicfiodMOqywRziogxNQiXoUa
aqNmkKAgJ6cG2OO4Vnn0dCi7sK/+Zw56qBpZt77HwdmH9UvmFF6bvH5EqupExr3z
IDt+8eE+9WqpqXMhbIO6E6O0ZodB2gAjZ3+hPK9YFCjoZrdYBhRlLUOueuEa5gPh
0YTKOE/k1oOi3J5ch3umYkKW448cX4JNWKQOm11EpPGd5t07QuK3lr4iPpudNYwP
4QeXsYqM5iApHc6D3tQukNVzm1cpxf4H0A//m8Aaa25N1tNGtv53byTip+5w+hlU
wAIb7vVk8oMXgin4yfH3uCGTFg4X1SYKqpYR/PUKgd9O0pKji6k1ZgkHHt5asU2I
qCUpZlqURSyqaTE8qUlCX6hWmZ9pJj3EaWo16GZzSt4WYnma93OSjXS3pMUbzn2P
q8EXzCIuaFY9c6KC5WCoFv77dsn2xXcWCM95EPxfVDstFc00BL3+sV8/X/rr0ZhM
J0FJYgvXIRHbJI3kO02XGHYn4oG3YmM9HCRGMFSgJ8zTc4NCCxhrCDU+vi+iMJse
S+AM7harB4GmbeP0wom5s6Br+6c9IO/8d3P+boIApxapoRAuTA9n1fOLLAZolGj4
6c7yuuFJoWTNGsmOIZkaoBSxsiHJ0m8cr9KsJMuZIIBcfy/sjvg9Bb1GCsCiF12W
AHSRvKNgvnlGwBG2cP6E0LcB+KGm+gCm2Z6vprjYy7T9owEnkIIC6ODX4jAukF4H
xF2aNcxBivf9yPqQMyALYl0DRWHAzjpE3UEWhL1UOHvy/m3k8tPBdpoKQCZzztxW
wp/tghGydqxAde5jBajPs8WSo9JvfoB9RM4TyEJPllbYP2eryuVdE+c6JpMcuUrJ
S/TTy+0fFokCO16Tb8QeddyqFSZy9shNGRxfYO4siw0cq6sGtjoQsEf1rqDxMy2B
pgN/SuJmzFjcKxRZLTQ+AM3QZrPnVxvLSl+M0eygb54uI4Rx3DVqHVCXyWimxLNP
9bbFMl0YrxLASLKAFx8OAeLlCYNPcNMQ//splwGAz4v9uXdVHWGXIMVzyC92+MiY
qzRXjwh/AGekDrHinm3HOq+6oGmwRLezSXIagIzFZQBCXZIWzqcG97E+j92der4G
NqxGHNiyNG26MWDpUWAmbmct1mkWwKD0QMe7GLq7UWgUouSccMhsXZ1o+ktOrWED
W3GqrwmSUCZ4IMi/0Zf4Df+ecgoCtjAGDFWcvbn2LRv6pMz6tj3aO0XxNrSMTlan
6Gqw/+n/UOgJbpKjr1YvtymRWr2/CKIjCqT4OIeRMM5IZU/9HQhxHiEV2ZXrA1Fs
0rN3f5GNKCSeO0MjnRixUx+TEJgkpn5qatfXytlaLvsEplP+g70N1BIi/9R3YwqF
iJKK+brI3fki62pict+JsRm3rcqNzxZys7LFs7yfi1MPL+2TFwKpqGBwRaopGt7Z
It7dH6EDCmhSONssDb0/NgU9rpL6LnmRw1lVO/NOvKA2VT4gjUY/dLUfUX3nM+5A
WpMtshQxe58WNGP4DXfkRqDB5ZHGJkCgwSnvtAbaJd2vRWlDSx9HgjCQlLXAwchv
CV3XXnjkefizmLgs4YPRmKcRxwurLZVN5bguyp9Iut6xzgIHvAcWx7zHWbLrP2T3
A0fdQ8NoQIjrs3Qslbcs4PG7+4pg1mOnVFJYI43tjmptQ1Py8T+noSq6O76/QqUH
s7JpJQ/xAJT2pq/BTKeaRBjPVioDfVbrIautpv+ztZYdo/NxEDTC/q0ZnGPbj10G
lnmWjgKblQSB/4iz4uzaFtXBnlgN5iIuemV0CliqexmBepV+gil0+FxS+CK7qsJK
HV2FoTrRBOrvbUyA/1wtN8AFuixasLmddZ3qdLkQwhQ0Kgz6a8dzowkQvxl7yIcA
py/qHfW7hw9pDa9NjA8fEjTUfSKBvcrCRfybGDL3szwE6CTAbEI5K1DKmHFkCXC9
aNzgdznreUkunUfDJYt7zVvGvZBuKE2UVRrh3hBtkW7eMsTMjd/6N9eVPlNysjDe
TkyIVvTsazYYK1fsQf31tfRdQpfi7KgjapYMnFo/vouWsJ+eWALlDjVblkdGq8bL
02pKRfP11VgH47AuViEiuzXtrp4L09rbieke5xPyj2+0UOEaXogVVnQlFzpNHIZk
eQcCaLwWJZ284qVkVLglHPy7Qb7IQhaYqF4RgY+FeXBQWZt6Ww030git/5CWB8XT
hgdzcDto/6wW3vcMqBZ5X/D61J1dnGPMsBTXuKnBBFjae5ZqUBTKL3vdm7CJMkYl
906vOTLL5A0zogIj4YDhUrv1PF/OKpFW9/7tct37CYnVsb/gfx7ec3hFV4n7D3c6
0cs9/hrXpS97jR0gNS5JtgClQ3QQICn0c8yI3u1TaHOURo+9CtgQqvq68ZBTPT1i
SIZs5DIitj3QXUsEYPOJFN2PO2f48/fpCsUjX6LveTHAIFirkJ85L9DrItQnEji9
EHGqJjGSpkknnrxq5Kg9Xn2bVoySHqtMdNyNh307pl4er7qdnqBdhB8h+ny1B1NY
B+Re9q5b9ppScWW73H7yNKghywUy3oP+morIIYxRQalq4DmIyoDSjfMoEnzZcet7
ieg8UFzv4nFk5p46kipu/bVkvNB8yzQwAYxSzx9cYRkkPAd1b4eHBnamhISzGadC
iDcF3hB4yWWkjXFkteKtGfsGGLyZQVOkHavr/8MOGwzu3/w4osaPQHIzMnQy2Aku
EH1StXOgXbcmXFy5gVYWg1vqdGZ9/md91iISDuLMGBGgAHYoMWK8B2FaIiL4V/2e
KwqshtENUwHlVL99bekbIaLL4RTxGpyEw5kFNUyHssDoe6v83FTzXLI3EXC1tKls
IirDg8gGzAJbsy8URbaqYXxQGu2gDmRYz2mSUE/Wx1MEpmMKOs5OQ74/GRtCOMH+
Z9vDCjnicFtCodGs9AIhmk8JyeTfbscfj+aSnnWnGllY4aeu36xLOGwGpYZoAkEx
fW3L88HC2JpMJFNYj2foja1Czesbbxs/x5hTTRinmX7mMZm8/ulcHGyTt6I9uuDu
iitO5WsKzkzHlqqtnyamSsMZVu8oYU8TCzAHrar9QdE65NtsT/rU2TqquSkvC0/g
w/3Oj51eIF8TfHmEFbkFwge/Cf6ljs6mDti11Sv3+VYf43v7L/hb14MamUSAPPQK
4DHAWt7rJ1hi19Tx39ATKcmbL8XFFE9xaNaSBLbEY+pjG2BLmA1oAUBh79tFw3i4
PB1KZgI3H42e2B6DR7R0iwNbc0tql0aTkhGAHwXggfIbDeTlVhLRAajm+WE5PvhI
qflNCqjWJitr3Q2jtEozOB4oSlzlBK22CdhUGNujb4Gw9g8PMQHatlEOIniG6Tf8
qevKbuSXK6iIvScxaK6KbHnsq0KEWjCdspifrAH+5v4ANKCJ4gWbPe7Iq7xfK/6r
KfFqHjRH3xiXjs1naQq5I8gSTkUs1A22SOi+FRZJ2XlG7gse2UAWbSj2ZyhNMCfO
lk7BfEtx3+uhE6mftrhvk6bWrUU/nhZZCXynhqQE3G6nIermHPrZtLW8JRMr48Ym
Kge0Cf7F4BDlZjPKX4tuFyHxk7Vwg410N+xA9CNu0uQpa9a0B0v4Y4kJGw/FTBwd
V+4yu9IoJ0rHh9gKa/9gG1cCvTXuu7u46U6COPgM+mFMhn2nMautxOSnG9czYcWz
6GgbCTQL1HhKBro2gQDdSDlVTPcL1d5RiCnWTzCQkzZO8JjtmtWT9qiL9EFdy2/b
NFE/a0MIqxbKDBAia57RQLN59CRLnHjeAd7BtBJKovFlKnFQCXhqmc49DhZtgA1P
zTjCyx11lYCTadyRZpbExp43L7AIh4l9jrlg9fspnCM6oUFl06oxhWlNHC95fq95
1xX2v2U39UHyTil1SY2IagjS+JQrw4qjrkXZUyt5Y7Ekg6aiwCoyt9cOheeG9S3w
7Bv7GrmDtZ6tlptPdZJApVizJeisADWZyUo3RAMhxmDVDxvhU/LJKM36N4Sv33Wr
lG4O9kzksUUfbRzEYC3+TKCIlCgPWyTNinQRnvNLz9z5fUrKGYM/dWoLuROil2Wl
IqWkIvPJ8ysTwB6jceinWNVaCq18gUDAKBBM5G111v83MLo4OPoHjT6aVN0v3Xcl
6IFVIGk6ga0mgkvomtMlkxUcZl6RaUgtm3esY7ZZvReSgzaI+qG8nv+ecPgXvLvq
HY2VuMqt8kAB/ReyR2+avFIn7F06uk3UF2scuj7E7Ubv59xc9xVW1ldhYLF4MXSF
sNc9My1i7Fmg/ZSgdOB8l3RIzJnlU+GeFxoSNjySZtGh+KHVty+n7FPlegtCafee
cNJj6wnx2A8waWB9SxCXPF75SxZWv/kEFRa04/xgQC96PUfuhVQ0clEH2Ws7AUAK
5gJevzupnnIrLL3LtspM67PKaM5LOyMpvzRlzRo3lWNXsH+hePjFVKxcin8XDnut
OXbAfahMR8Ny+dz9PY3RLy2mzC0xASsIO/PQQotuVcS+f+GTTLdzo3AZxcyxLGWw
OwgijUO1MMMb3xg3w/7QTwhXZ405XARfKdbnQY6SMKsCqzzK2zH+KS7a+16DvhwV
GHBY+23IL48X3z0cRoMi6nKtv5Yv/Wrc64JTxj/kWbUogzeK6j0HLnSZQ3ZkbldK
Ykh/VWPPOchVK7Jhm4kvKAf4Ci4W/OPo7a/aWBUbnf7q2C1Qy/mhFEmXcau8A7Uh
dnMVnj03Uf4NnDrRCokwsjju6mkYpXKjI1W9Gze2m9R90yOFs2g1n1v6jI+pyFRA
U4kafY/o6f0jkiXy8z47vIwAwinTJeeryPGVa3FxCymzuLgvLgEKmDLWkFWKcOkH
tmuOuX9MAvSsaOAlV0bzq7WSMm8FFlvgoKu3VsD4TSYYbjpluqlbiVdgps6RHENA
xIkqfs00BTZiZPK8PfVyYA2Dv3rCmybj06mDlFYv0sTtCndeEhShBHR0uXXaWMSr
Tw1EOOQo6SvGYoiiYVVLG20GPTqOXs4DUNu36pgk1xOnMnWxE7Jt824ubnAE/Pgc
B1puBig/4VlftGcKSPGGNTrHRWCKqbDlQRbgWIrtY7r3KUiYEAfLiuAbZJf+w0nz
qmo9IoPchQgBtJQ6X50G0+UWpO8PxaLx98hL5KK1P5ZtDV+p+70feAncJyB5mRCb
X/W22Bo1YuLLfdiUYAmnn6ZLuONjWiynvRa1ILqT7b45n8ulDdFl3MtjAy35AIvK
yP5zrcyftCspkzAjOW2HwL0CevLT9GAP1EVuX2Aq6bj/Pjo77DpgIR36v0ETiZBU
BVCI/fxYb6ShV3v2bdpDqc9wV121AjaddMc8bMf9gLgi+EG0QDdUzjE91cE05A1U
Oz01TcZUlNDb8Sn8tz3hCrMHHuRar80eH9fz3Thmg1tgpDveuacIF6B8wTa3NFxu
2hE6Owlur2IrmDzLS2Xv2BZ9/yP8hUZaXtwHOhAkiH5fFRqmXOYXjn/NAPx4Zs06
U1JUSGKtxCeeimNktib2Q3+iZrnsHgqxpx5FtYLRagX0HE6jcRuhaXpJbJdBDaoE
urUAEuKkR2lwOXHRcLZwOX+OWLFrate8/idgXwGJWsGOpUXEExMkiE2wtUhTWecF
18AenPjDPDFunaCVpYId2Adbw6RtttHc2WB0yI2CkTjXwxe3/hZJ2utFRGyKys+K
0c8eGov91su1d+9OS6rvXucCL9ApLDDFfyvTKnlh6kzwpXkJZIFuCmC8aGJn6LAM
dRvBW+DtRHZXayKMYUzaNrlZVCkn0YuacrEEWLhgOpPBclNLLK4K23SKIllH60r7
ewz4ZShhAiWfldmly5y6yZfMzG8Se6xcr1xVoR96JdcL5cXlUOQdMj0n8j3Yx8GT
JfL/Bx4y7qfkAlNFdlDowT0O6jpIrrVs1m6vrTPruH10sOW6C7Q/2EsrVJF6t09M
Rky9G3IzGFw2+fiGv0f+hC/WDv6wVyiIBjr4P9Q9RQWsh/cs/MTLe3BNBRJeey7C
ZQdgIu1Bd3+EVRF2y15h7lOcFxn4UdA6RR2RJ5CmifsLa8Dn0sjf3caFp6uyJX5N
tPBM8WIm/XRQ3Wt5ptsR5gixKslb5b00BPtKpCwYlwRPoLB6rXi5IbLCtxxXblNs
8lKkNeEd3k17f1NUX7sMUh3CW5p92q6cp6F0ROHhf3wC/r3drVM/RZzbhDkRNDte
nyGgd4Xk+QhlmsSPcvrZaaaRXUbEFJ0YESSzEVxJk/zU0UoJDPIdKjQQdMcSXxor
sAYBFbQxEyNwlo/ptkQdA2n8LnXYkEHH+Ym1kKkvcCCUglGQxHxhDEI4NkODzo+N
BPbDiRmbtIAmUAdcDfdkeEUNIj7/KsbZzw7OjrttFpzW1VLPCqu06vvolItlF4L5
0FdPZsrUkWzSdTpKUCmtQxH1n8pu94PWOoQYA0fmPNGjvwAeqCNSFxbVOCF4Ipvx
+XLiJ4PdOZhuLNARtWu5jWyYjr+QBPGTjFj1Fv4jYLbLVvM5xLLENCCZFiaQZPLw
iP7uG84ho+5B9dbOQKJYvfPnrnvCk558U61A2hen14NQh/YI559yhHMirdcaDTQh
aQfbeHHCn8z6VqYDb49j49Yhbym+ncidL1trCIlkfYJEsQ7n3lVffcF9Y/1m1Qwh
hDkF9e2+fNXFkO5lNzrLvt4r89oCZ3MHOZamXkkCF4TgthqK7Hyff11Nmzbj3u68
vMCYRw8rBeWWrK+LTbn8c+TcGHPqCj4oFJIen1oBlXU0qNeFFdjVY9oRcelqljhs
84HdEBrqZEUIZaUG20fjC2hnN1NGwafxDdtvtjOO+AAKXQkuTJCrdptmNQtFfVyr
AfrRvsq2w/N2HV3GvjmBbqyPpqmM8iH9JIp7ekaHrCmNrPMIhqoVP1nGQ11LAyOx
sHddo0nPfgXchtSZtJpB69xcXQnzsqrs0w3jxKysclLBwDriSq/eSszt5jggFX9q
MaYCmqQxb/bcfS04PXomLR23ry+gqFOKMk4nnjax2bUdt1hcOHhTNU85je7hcQlo
1CMnbtQ4lZCkkxz6jvwdnKyZo8fINDa/ndHcyyzbmpDe41enEA2t/aq3cNjxzMRX
Pb+RBK4k3wbAr+GM1X+u5R8+ZMxBXXCJ2Xwu7kJP3yRk+0DtdhmM3EMXoQ+r0qOC
yodjZpqkBjIjL8iYkkz+suB5Os7Qt1vi7PSGSFkyBn6rwm5wnT595W2yUJKjp4tK
ogyc5pmzd7OBxOCokuAVIyEkubt2iHg739le8fja4XgKK04dDtNwbAYAEM4JU0Sg
ClvMRIse+QOBrUwVUu5+CKkdpul07AHWdCwpOJ9SuElL1laZFq2ZjalDTTRb7LSm
OFDKD+e8z9HR0//3vd1sO8lOXC/26J/keMKnJJfe6e3NQfuJpFxNgXvzsUHK8BKx
i0NhGd+CyjeZbskqULYMmQqLq3c5igOx9IZsfXh/fL1QFEC/0VWniXDLpcaiMye0
ZC9ofivymKkX6VlMbOHCr6gWbjxqN+lfSdOYvRdS9e5aomVsgsbgoxQQwlhP161f
JG9ebSDIQywcr7B1lAnnSfVCwJJI34S+/Wmecil9Mou4gJBEwZ7DnRGj1HmccqZ5
kNtTEtWvSNV059P1VNpbjyZVXL8Ais52CTbHzMY0KAM1Ezk3kEk3BQp0DlMLwwX4
IRIfssDF9+hiZ5BCoKNaROWvJu5iviGk/bD1ahTcNByS/ymtKzRFtzgYGU/h5ofE
2L3F/Ow7rD6YCk7wO49RnyOEH1bxqua8cOBr0ReW/GIZQmc0fZNdqb52jOOjwU18
5xbOAbQJW9lPaHGKETUwyFok04kdHOBm1/cyHmdHlJnG2Yz89CbJIatq4DqGHM5c
ihhITTKSKjYmx4oqWoJGA/WUPidZsda7PaFpK3n1KR7ga5hqvMrte2iEU0OQfzZu
IRo2N/LYilU+dje7WyLStcczlpH8lhMMU9S9HMEJmjiPhU0IqoNwUGDNmd/dLdgN
b2By1Q+eDoqkpDHX+jEraNYl0twPD8GXBVjIEqRH8urlBrHbgyUqdK6wp6mVpe3Y
pvyyMvj+Nx9SALR49HH1QRrRX4sJ49EqutEf5ALNRegedSSGCIricAHnOweXyiMj
Wci5sYlT+VNIe3W/5aZldE7TDjN3liCiomNQlxGl4cR2jysA8uxewwzzO4ZtdE4A
ryulzkF3uPKYf2USeiJJhkX9XYNL3FzjPkp3ijh6yZck/oiq6Z+iHy7tQdBRWVoT
ycQwCxZ215ycWys8vBL7zska7lHuA0+AxzYDAZzc8XvGCztiOIbDb1MlFDSILfm/
SMqybtm0zhX/wIahm2t8iMTLJjm7T/fzKPzWlXR33yRaCDXVtzIiPWrCJcWrP1zg
mLdNZfJ145SciFoVS+rS6T5iSNps36gmR8waCsqhKp0zEG3poMjUQp0iM3XV7npG
932GM2a7QBXOmu8iISjdk+oLQILuKcnJ3fN5RUGiJGuHlqZh5l2Lt/FKztUOkKuh
fBybxRHqhjsoieQF6urDpfUbR7VFP0xvWhDQv4DSndg7gydGhvV8VZVNTFswCoZu
RLrfCkzkbKeVFxJOa1PCZiWLhaErH6u+rpcOW/8NL+olENf10yloVo2ZdKSgPAiB
mYyxBIkb4BDApFdvOckPiZRskzhF/MgIUjs4xATNPUjXJCDAa3KWubMmT98Q/kRJ
IW8nwX3YfvtIR3/WE/mxVe2NBxG82YkkSbzJrMtpobcYhTLZkoCdujhaUWmCtEZ5
etnXNDPszItq0ndJD2ruxvUx1XMg9rXipJF8sb1Ng3SM943G5W9AI+VAq8E9mt5l
hOadS05ZIxX5/Aw565e5uyqiV1OvVcT4WSo28WGxJ/ew4nqxQKKbY099grCSLdEW
nLj3ypobE0WPBZkybNF6ZceB3Bz6D6aPwOrOTUMosAaqGF8mV3IE0/evMgnpZYIM
2PxqDHBPXSr/eCa+86hp633anwekw0tsPP8x9zJt68vd1JtL+l1O/jxzXy6hJYeh
`protect end_protected