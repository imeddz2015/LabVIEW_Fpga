`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 9632 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/9huKRhRMtvnNqb3Z+UU7TahEoHV+T8U3P3ufru7l1O
3DlgtZzb9QxCbOjthp9+wDkjygH0eUfDrEl1ovhZG634qmAsksck45UkVlLnexN9
9uvpa/F3sqmrvn2O9I0e4X8BwEQkmcS3ThRMKClTJWJ3MRH8oyYvHCuUcIIjea7L
kT6DjN35LyWINhTmwxNwFDXFXJ1Ilulesr5u+2yApYZAAYXx4RK8NBQLjyeedE7s
VCttdWsVQHTCjpAVMiv0+X5ffsD0b7uf8AnnGEh6mXWmaju6mEE9OHUaxN71AjQm
HuN01fNyPmfaSBwaY9FY2HSr30haP0VBYz+m9WHMUt9CBo9sarv8WvW8GPi1m2oL
g8ikegz0Dh0zYp885v1i6W6T66GgI9Z0nYP/bSrnp+E7urw/MojLwdiOpG57Ojzh
k0OdoBgQyR6a52aNot4zB9J9+0lHfC/5BOm9+uf1vbRdw3NcnesXhPTlovA07mlp
41rF6q+DU/XLVCLRxHAL3ttOBHEcP8KRV9xiPDKeZIPlNdfyXFJlkANq5vXlH3Sa
Ax07+txM82zl95OnD1nDx9zwHgJJ1RoUuqnbz2iMCcBl8pVkwWdt2fwiUvbjR5mO
eAJKF0j+JvALF7xeBq8qgIw9JC+n9JCzVEhDomqotTFU8vT6jJ1JLuNdb1poBwrd
Z7Wmpd5N6iWSUVNy4EeBufcsohFfEyw29raJVNjbD4UMq0gQHlRT9p3mOMUOpvcH
U1y/ujX7b0BGmtiCWWDU9V/1+Ab86vOiTDib1R3f5eKwELAHRva8nldgNbHqtSgg
+ji3GqZe7CDFUlnkRBCsW1y9S3gFnHon/66Qs7Ov4DRWS9iJsdX00CW4emPKT/iz
87umyWiTPUupkEjyq0nBQMzRAq6xzA8AZ9gODhJoBA33UYjHMn5TLbkFGhzO4uAa
0ZbMOxJEV+qu5taQF5ifFsdI1ufCVy0ibv3KB28BZVVB1J24c27eWMc7aUBasVBP
Q3scmfO07iBYftCoeHEjK0937Kq3Y7FmkfAwPWMQN4sLcOysvPvdt0HNkvuDqusB
KksmwnwBZgFuNCaU97CH0+vCD7ucEejX7srlyoK0goFQ7m9ydeZMOxO3jC0kVUCh
7FX1Jaq9pc7Xu4QpC9uu0WMeybIiUqJwbQxL9sg45KPnQd55QVnkzNELd6Su9vZw
fr+uco67Qb3MEUIrvMVusOYqPuqRWi0bwq64bxzfj0+MGR20kwdSwHRsKhmZaHsw
4fJzhibHpNN1STMP3aFBkB8FdQkmKp502GdIidj3km1hgdJ0qkXsmouopVnUUpMB
xzdH/KYdcIN89tS7sE7hZRnv7Hw9UubFD2jcxrx1HFIaAP9ckTxYFM2OnsEJ7H8u
He0ZrBm1PXapOnQu/BiUcbV9DB83bc2PNp3/IEhmb+GjFj86P81uFi/QFxC4Ic5Z
BuTSg11ZWIscOsbePcgunB0DYwqm4d6E/daJsq87oA6nr/RqrkLBq0XJ3DBbXzcO
ZAbu4qwxgTy74qCwhir9TAr3bvUmnheof+IJOI0ks5g1MtPY10LhpoHeqGN6FdFh
Zlkn2Qg8Yk2oXSU0wxvARcaOW1HsqKhIjYwymgObi23ZoReXJI0SQZXOUlOB4UDu
sEJmCBnaHKnjcqmFddAvaKAYXcKY6N/IIe56ln/bEgMU4L3MHE9yCVApxKWjkGBS
RAydfkN/TG4uRACINVCLo8j7qk32YyG9VngbLrVwLLYLYpQe3OzNgQjUxwKKv+l+
QIPUg3zu3oIXOWViyx3L//9DpRrlE1TRCvz+0NnjtviQ9+UeGbRDEcBPZrWO+F/m
L9btMFnmZdsVVD1A4VcxQxvm5+YHJjolU+938nfyeb13mjU+I0jkgofcNPTkbr+w
mqbPegQvs5Q/JKqOjqKPo9rGOTig7VuQ+tK40TB9G89m8+699vGTqLXV7Q9LJU4B
h1Ocwko1wa+6On46PuxFnvBBd/FH+aqP71y2II4BSRwzzxxict5lvych4P+NIWq+
QqXU5OEl1oPbp9kNj1QiUWpYzBG7ULxd3aZOWHwV/owFM70dU6Mo7OSSyw/Rfa3/
DEpyac7FMn4WkL3ywCHKeYglsLSHfJKie6LBOH4dYmiSKzQ/r1bmIsNHqZn1G1mO
h/JARxJWY1wVy7wJJdC1pL1idSVkMtJM1EDugqGQvgZOx7lzycAbJeAU/tbdxkUw
+yCyp4L/IegO/79VtvtlHzucvCR/PMZrdvLgjDzL6KJWZ4TenW3P1tuDneg4yP5z
h/WgHmPlWir+4CM3KuB0tSk8PPBQtBNMTJ4tusn8P+plwwkN5kJVb0TG6zERzABb
x+2o4YSgIyY8qy/HP+J81vkgGVTSpKW1t/rxGE9RL0efsAXfFwAZhoDD72JwUxWR
kth9E3KWYh3vHb+lM/b32I7u4uWBxRv6JD/bDUyX4cJd5DoLE0mLmE9m6aDd649Y
u2kqgm7iBqcVPNvLF+cjBS6s/FfTQx8DwEwhJOXTZStevY/xiiUPLWQ4pK3OYCQi
hZH/GjYqKBfMg6s5EQCRkbP/vM0qnwzqIZWo0VKE7cJDYWWd2SelFMwjm+T8nTof
5jpqkk7NLafXrVIWrayAycxcFboNdLJdCXYDs1QHtbrGNyTMbchLp+/t1pgeq00w
bxXPdy4JrsIExg8SP9uMddnvzfq/DWEzaGUaTxoxgEUEfUa0zEH+gevuoT+zqUrq
Bv4zy4aLfQZN8kuETS/+ft4UMGYJVsqNXK3LA8/NErqITipURthYOh3cWXq7DLrc
6GMo2q6n7Zzx4F7WMVhNtGJ3O3spjrFYBXjYS5DwuWE9PrsTddkAME1qzt0oXboa
tAIGSHc1rgmaOClca51lSUDEG3Q1Z+lWRJ1lRxHZFIqV4F/9XwCmowmDu5adgpw5
+Qf0Zc3lPNIBjwrvLRGcVeSiW4X1XefS0Pk0Dcuhg4zySrP0kYR90coThA+lQq1P
6o/clz1sCU3MramESR1fiAxNT/S/S7dlxmf0iosaCDjpVw8TdJRtEdersyGxGeRz
/rOQWQILmW2IdEPhcM3MZEQXv8HQKss3wVFr+/qCLtvYKrDeO1hl0jScBJ7ZFCCb
FKe9ea7eXluRyf2TVc4pBDB9PLU6/8nXTbsg/IiK7BLapuZWsobisRSvS/uU/RZh
ewEtpisV0zIBqPzibq0P0sitjw4eYebY9JCPHgY9wtMKCzs+gusrEu3jwVkOOewa
6qmq0qCferZ7saHzx/Hj2O1I7so0HZqejfuYuUsvMIiASNqntVeB1Y/kOEldEZnT
2WzPalWjIt8dccT3dBWboGmKnQjoUaHHqLzR/jIlK7dztZWpbeA7NOR70dlq48ha
80PG4Dlf2AvDMf7kF9KivhPqma8pJLYnHUXrXsUixyKwaYXTmW8x6ijc1tdqhhBU
8I7z0tEjjQt3y+SSG4wHHY/gu3ib2GU3B4KAJjqOEdrQooGNdtPwOol+jyLUwv/0
ZhAnyw1xoJYxrVJGvWmZJfophfC9Be0Y6NHyF1ntr09U4ZCFUruxF3tsi4A69phs
MHRNPR1UuAeXrJbR9UzqggPKaXgfnGKPgQUAyvuFear6q/xXigcIwpJUdzJ3UP+l
xDmkL/vnh1aZ3/hfEz/LhVrZkFS/epibOHmCnAgH/hNeqOxQr+i1tASAlNiX/qsL
IzIZgkg98b+ID2EkMQITwMPx78tellgaCpKq4cudLwTw5a9uugGMDw1tMGEF/EAT
ruyxBsdTz+3RLX4cPZ+jpPnGZR7otp6B6y9mOk/yxYei0OyYtTWtUQZE6ptNa7Vz
DnVCX63H/To1mnmBuEBLSNAJgLCal3EBoVtUclxQFavoJpXoztvmnHNkXq+qeKQw
Urd7GNBMae6bBbaVTeJZd01WD/axu4876e7JsV1Ot+54nUbCa5cKhYrVkz+PNXbk
v7e+Ub2aEfmsjqGi90B3yiy0CaS1bEDICmuB3+wlWFyrVtaBTrETICdtZ/gcDRMV
3ZE30XgsJSR1j60sEjBIxZHZpcrejzN+DapJgHg5j7puw8nc2Pvboyw/IvEbK8HN
ub4zaehk+mE48NjIYXoDmbRDIwM2Nt1fqoqamUgBaeBvwt8VTsQmzgKCOuCkfsMK
YbMSHA/XFzyhU/HbU5eWA8WWWXo/wPblRXGES05cfjqYIzIxD1ZhOXb5Se0wi6V+
KXBtHQbPLSn/x8TXxwtJpdLvJvK0PxaADMvy/yqEg+Sv2Fnf9EuAivOcD9BLcUhJ
j2BJ+9ca67eCUOQ+GE8x8aLUr5OL8g2nedTVSY5TGTGBwbw6FHJkq3JcvQfQzJWo
7vyqG6rl7uxPn8nz3pE3SffAkqUwteOlAvN4xOhj7R5mT/9ZF3xMfsqqbIBYxf7+
dLpZu/UZ2RaFSPSGKYmfQm2N1nlQfxWSvtvvLQsuviCXsGtYO9hZbgV42lauZuyp
1LKBN9tGpyGtzk0iUThp9PwmpBYuGIPNotFU3uHVaB2FoacWN5LeSjLoCTHeUgRj
qLq+Mvur6Uhu/VLJbMXq6pvl1Ec1eQDwg9A0hxnhV2bkDP1UaJowMXqZFDn4Fm4h
7Vi5TCVs32doLBTBI70PJoBYvHRvdEXIW5+GNISDP5V6IVhUmEVBBif+aIIVAZv7
HZWdRN6Qx/VTkGbvsStGH6K335YA/a11dSOnWoGZhdLSrkYXN9rkOKe2/CcM0YtP
NPIfLwR4wIqwW5p3FliM5NwMn0P6k07dvQIVqyCLATeMbY+1+BNo6t+qf7mej/Nz
rv8gBTNVo7rty+ju3sZSTvZKzOMusYp4/lsiYEMNc1CG2QLx/O4C58h5t2olhVfX
XE6VGkyYRT0DXCSo7TiZxqXHCuXUiZrNduhBj9JMqU/UQuPYA5WNNxH+klpr3eIi
uNVECiDn51pE8LRv4a4sNX3+H5Lk23Hq+9A/opc8MhXwGJ//uu0gM/gKHR3eICck
5638vWlQe6xFy8llM/L+4BAFpg3PNNVGQtk6yCZy88zt+oDATEcYNn78H+ZZ8f3m
D+mNQCVBJxaNJkwogX//afv4wwSrVvZaDM0I4xYhSF3oUMSuqmYS7oCbluZPRkPD
m+zlvzEv9u3XZgx/uDB0hA4yEhZF6rE3HO77edJhzY7B7ge9qZyvegxG/7aFFbAF
VhkVqWTH5z8nt1S+OtLXgYqhfurQWXIC74DO9VbAJl4QG94eAToJYyjNl3FhsSik
HdRqjdkUq0r3KXfY6ah70onDsH+PChvj6QISCBWbc+Y4LE7AONldHMEGIXT4mymW
PDLUxj0TOuYzpUi2X/s5iogOB0ll8IHWYqMJSSZ/744vuTncNOLNtJfKh7VxfzQt
jOemiAcbZiUpShB4Voa+mf4bX/c9lm7C7dpzT96eAiywAqvCiMxd3ioGpRGVu7Os
32Uib7rWGbjUDAIsltvaoCwMWL9n80BJQQJUPYyJNvKfC7tTWVxUc5sfcfz5Jnru
vl/mKs3qqMK2dsVQecDanN6TS8ms7Hg9WvaTZSJwcPiixEWY4kT8Yj3lMB49rYYX
i32KbvvvpQaw4Jppis6R+Hr9P8xhqugEJJTzaJx/de1zgyqDfU+QyEo77YLzv4xe
HoYp8dxvkFFsM2VbPoqo0XNgHE7pVCGXG2b/shxDMA2KaoRYZXI8IzoPdIpmymsR
zHvbP3pmfyZc7bFZwyxUGNlPmeP52rIO+QkmDampRnIWji/odLKLWmq84jQrN7BQ
EcjrsG/21vJXun42RLrjAJQBR8KxhPHeAZN3Q97AFli+Hg28O8o26YtnvVp8mveu
VU47wzuOvFJAKosOypfWrXYp7QVt3BlVqBb9BXyFQ/QQe5K81VX9lcf0rmxasyF1
htmF19Yrnxq0W2UCCeA9paoozgIUPyi3cadkSZJbDFfBqssuDKui+T/gLV7gyI7V
6OwE2PzDlc2sJy5ptSQBPqWRjgNkLFLr7y6Z/KLeu69mTTreZH950vTFYuLZoUtX
i4hQw2paJW3OeU22YM6NDc0/M2zlvkyiVXIHgvECBf/ZEOg28bsnu1VdJ0EYG9b6
1LPhZOfMi8itEQjT12gV67lYoti6HWnlw5+89Kr+njyfglmi839/iaiocfs3TFEd
GBDTuemnTS4cVrEeX2yLdVWRdtcufnysvcxSd7LZAEAgdUAHIUJZXm162j+OFqtA
gCkp12fTBQFq8P3jtenJTwrcKO3rlHlu3zUJE2tQCJA9Nh4Ykir3Tl2kr69DD08U
s1I/WgnWE685hRYrRwcJkdHPXbV+IHH7LKqJgdlhdpzlTWOhmfGXkiLLspgtXSet
eAqRbJxipa3zNLQ7EcWHyISXBrkMrcx5Pe7ASl6n+Wxe4+1KRR4+QrzMxiz3NWRJ
RdtXICkRIyw3UNK0LhNC7ah+DcstxzbyWcKj5AfqkXYtLbhrzN/YBoWGIVIksnTN
C98DHfkPAuAuVbOuMpQ0YsPH091MMwFUSjpioI5JvroDHcRXSLXWsxV/tVUcj+go
C1kcAZ4WX4pR4ZMVjsltM92iV4qQs5Yfm/I4dlKkCigAww29DFbO0hRKvas5fnqC
Q+GpXkpopTyx0Gatk5nw3H5kTtXjGza9vAvoAB7lRLQ8F4a0wU5W3/+tI0zOJj/7
DX060Xvvc/zNTuV0+wNxxc79MLrnXLvSYwEEviMaTS2Od7h2fuDoKo7p8kLabEBB
9ecOA6y8dAqFLz5IQkgMEyCDHuHqi0aRdsekpD+zMpF0tDtibKeh//dJOorpx/+d
1XqYOjCygZytnxPhi06oIAOGtYTNezm4KBQ5G+6PuqPJUq666uY+5Xbndi+FJkL7
tJlHFrebOHf9eGu5GQWfDm52Vg5tqkj7aPUTzmUfG8+xrbOCn7qUk0RaDSOatIBJ
q/d6fjkJgFTkmFIXokAKyn0pcBn2yqPbSo4AeP9534kaFkAxcs/fg6z7k2acy5rr
NId2gw5Ow9PbkBt0RYlI43MA1UaiztoBcAKtfbkU2O9YOQLKmM1fhRHIRkC0TS9p
eQk9WnMRa7hNkkjcjDkDPBy2ZajwXxI8o44x/j5NXZX4AbymCICJ1aigXagqadW4
dEyecpRlAS0hYj+rjtg+LND5/R31tQd8wNl9i6qIaqBpGh7/xazVzVKtq1NIXfqN
mLdNKSgh2wCfEWCX0IgFK1tWGkMMFO9LXWcU9bEkbjKi1h+hMqVdxvsSWvQKwN09
+Z/BdLsGCgxAZQ6br622JHKdQdt1WJQIolGWJOF6O0y+WsWJkPF5O8AtsFq74gOx
eKLAbq3z1PGDiyXFBaSEuhIjHfMUC/RJm4FJSKk31Fq5WLIeTEwlMYNZcmpbhKlW
8kHtEgi2vC8UPG0x6w7sxbqOpTiM2uEk7+mvhWZAEi0wXSIaxdFF3iYR9MXDt9gY
/wHdpUTiODw7Z3gOpjcAWusLtvYTMqro4rFh9mZwV8CCUkZKt37MtSjtsZtAwLrN
HsUgsZxAFcfUkMxQrARafL+X2ZD2pBb5+Fky+ROFGlyBpu3vIQTe1n7Jmsxla1VF
mwp5Ke2ze5RpKmk2N1Zbl9tANoIZbZfURPflFiFFP4aXesod2fpzhjTWCDAKv8Lq
qj2Gt5kPeDmp5vkgWoxmlhAU3CvZB4G5qOIGcBMbXvjVUt7KaIumZIqNpHglmTvB
EjgnEBZfrYU5siv7d0H0H7i/emwij/Wx0IQR1ffTibjjwLU2Kx/FaDsVaxRqsPi7
nQ6S38vNO6ZRtcmU26dJWMUgg7Ro9c8RrPt+8izxpxBlZxxl4J7QLei2XKPNSbZQ
MsNLcDF04rrZatcADNvHOmeMH4gwZBtEfcTz98Dvc4a2p0ukUvv50sM9fDwWaZb2
3+c45nyGBUdMiq2n2d9wfj2ii3p8MnGfUssCKafxECBJA2Mss3S5G6Wf8GCkbFRg
aJ0+mu9h+elhopDSRU7l/xD3xtE1yRF/ectRnvwBFvSADg6oZLR2kS4C98j4GfK1
6EsqoXgs6XcFB06wA3x7jIi9QLf06snfFm1/LQMioa7mcPhqmrUCYfI5v8abrhzH
gtmgzndVUksXgi34wJPVmNFfdlvd4RqM0brlx9qLfsEK7nTdpX5YhAoYff2CHlNr
radeHObQelO15pPB4VXBXEH030L9VLfQwLH9UUURxM1Ms832VQiJneQjL/HpDuPB
edO8R23ymRFahCKg4pS2XgY6MdenNiuC6FtjBuwPSr04h2e3qw2rLIJYifUzEb+y
+brghUfRzoCv7NfCO8yt5/RlM5ETVyUF5Qfi994E+RYEp6l2TPb/D0afhmGEgSBb
b6J7BXj+Pid0bJkMgOlViYqQOQUl5ZRD/IjhSvfagr1Um3eELUHoV/OIeApP83cr
tU+3zz0Gad2+ZkBoX/q7726tjzP+LefIzNwUiyZxzjv1qWflq+/PdoSZfPi2ZR0g
B3zujnjZ2WgOjG6hYEBzlaXtRPlAQhF7CCrCLJ/CZoGBNi4EDPIMHY2A0ydaXoMW
9qvD+KShBIfj3NkygzwxNvcIs6f8Gu2XB3KG+NjdaJiFyt8Nz4jeh6Pnmq4xItMX
50m8Jn6kXMNvkZB7VVZig/NOYmbFeiXo2mQGAzJ8XjdmagXjldfjiIeyAfyLarNv
OPwhvU1Vm3iB21YUbJPqOz14epXXSygusVtzC62SIvRDPoTN62Uu2zskInUwRbNP
K6ACzDVm0uvVXNVgsodWzCd/u46Lc82TTX3wc8IOMmn0KLsJdKdYCfm+mGnovr2d
PVLrWuyJxBKpRc13lbX/kVtZFkgAuzOEFuXeS1WoT7YnzqFyUSTlF7GcR8UgA9CM
o+77f7loEtVH72vW3qlNDDgjVVl6xYOFH4jcqTf0Agk98xANvrQqwjzlVbxqKfWe
x4EJ7uxKyYKFoMZdYayxH+0c09DnqqWJfG66/+9wpU3Wy3DVF1IMZVn7BulVFchW
PLPan5sQSOwZ/m+Y66boI1Je7hbVFwguhgpemXvMOo2c07O/lgbhj2a+yMqsc05T
Vu6/njaLH5oQlstl7u2g8gQRsfLEdx/YUHOYhRDIbB7ZJC4LJaYvrKGWIdQ7yivW
aPX/9URtTfzXyxed7D9ayf44xPKdGxhKT+f4H51tPIed528/KfekmXr8F8o3Sifq
ZMRLl4yY1sf15yKxPczmYgGLuqhWgx4TAsp7WWShab7Znc/czqtQIOx24ldVJJw+
Oq4e022W/j+9eBMMWTzfxPDXiyDwxQziFv9oW+Uhj1dFuOYQWweegS8GoP4+HL+s
UVakoQl8uB0qV6PV4GEIs2IxS4d/JBHjvWF/3jD1kKqd5Mvyp4rF5sUFpwrXUZK4
Wft/QqMASpkZVcwF9JmgRFvf0yER8swJzNRRMPVDUr8b26MViBaENQYLTlsPVhH3
5IwENkb8SQK4t+g+UoanVwpUHq260Ab4oH+mu+8n3ucOQICCoFg2qGW86LUkp2HJ
yq/8qNCFeyo49UWhwuBbXIVceqvrY+Qq8IN0+7zkpEAcF4jOyZoE+BLtERGezTkj
GCJrp40I7QFN/aMAbM2aoAsVXMA/pzUuiL9AIsHzR1FkfL/R8bJCnrOLau0B3beD
5pbLzgEK+foTyqnUFf3RpkScMJnHxkVJB3t5VNrFB7V0e02iRKggfMBqgkQ6DgFb
nJTkJhbiSwEFxSJWk5LlVyrsbwtGGXkYV4b4OOulSa7eKdscF5vDJCg44wjTrW4k
ZtM2NDhwz6YlokJUc//l83J4FUhJvia0X7BX82DHXlv8PrD+K+k1l1+sxsMOniCx
4ttDvyIc95+jWQwIvU6MPptRICMWegBB5nauvw+gomj3VD0nvcH/yCzfpVjJElM7
dfwwYAAlfx7AIdVQ82Xg3+an4TIhO1xW/kyln4k5b0aZmM+p8Y3ieGQKAx+1yZjv
L3bdtCrRYDXgTrYLC8msz+1w8Ou77SMlYN5tcDljsyynTCu3lNG7b7xvhQQ496cN
IIVX8yMq/iA3xzzAGY7BAUOl7VXiyuZnD9DfTCT460SmtDKh82vHtys3bFcSvmqx
ncrYUfwgYowQJOlIAJIfqS5R8ONeqGNfXAzjh0z9eUQzrHbV6QUeaP469azaRjOV
LofWPUEKcOXkHVVE8GU56h3djh/JsQRcirQyz81Yy6QUu26OLwOZQqC1Nub6oDwb
V9eOqJCvRl8Gx61RAx+8+5uGcBhYd/QajtlVJH0KQxdsvqJGafoJfAdyIRiIo2Ne
bwVtkTtkrKGzWheYCBZXpa2LrWa6tk7aNJp1hiWSqtawOP4ATOtGD6SU6SniaBsf
5RCAoAb7RUfJTBMinhcbKuoiO7zAz8hU3hd/O83yKk/D5TeOy2Yd7ajOjwLEN79g
PPCiV3dvIDPzvED31yKfRL2zQYD8F/dAaL7+76WEvXs59xLdSeRRAbgEU2JwcxaF
a0xeQXKlV+qxPCGK3NmJg4N0cic35M5LBoeAplmVuhWRtozgeLrf55cx7Wvc6aRr
NM+Oop6uGpXMWOrAr0uKBh/cmV5R6jqiLDnx5Dim34Tztxhfwhsvg+IUS35aaK4Y
qWvmN5HK38Zws7NaOfyuEiRSdTsbs+b4L5wgA5A7jk6GRCza025F79y0aAArVE5o
fJQvBFIgdj3WzWo/Szso0MXng50O+9pgz+ykJ0bkpmwBXq1+hMroeeYTYVYM8/mA
xflkMh1q7xagx6+t8Re/WI85LByvma8fNUlUatwfeXkYepM0FCB3ojtWu4t+twyz
a2yfc/DRM8p3bO2DND2g6fOWnfYW7hwpPkcycqkp1yNhpJQSA32eyVoIX3iqe18n
s6rFnYwbkCaB87q5d23XLxJfF+zj6Y3CRJ8+1pU59waLDpqsiiYGKa8ws4bsovgf
q5QiusAVpE9kyd6yyWl2qJVeMVILQiMtTqNuze2F8JkDFy2bZx6AT7aELBZEMmaY
0QSvenE9v4+cM86LHy56V88Ze+IONdFuco2KcQsgAO5bjaJeLpRUXZS6HcmsqN8A
Y5HBcBNuI2+ryYyhxqiaz83dPB9zzBZbJHnT/GyRFExZpox7ejuNcwjrDjQDC82M
LrRr1l30wBZag8sYZYnVLOMONfhWWek/hd9xqKRT+hMRQtIwlQjc7eg4Z8uxvaxv
NCx5jFR6TlZB/WCz9kA7YyAG56fgyykJCS1jQPiYidelJoINZNet2chXphxPJaqC
Nm8HjyIiHUpbkbVj2T6oWMXRkMEjU+NfHzFsCe5Az6F3hqhUFV0mXLyUGOxOxyb2
6VLnZA6PpJGRkTyKV3lLD7dZT8LwzzusvC4ZB5xN3zI1pRSIBrJvUQhcHz8Xj7ur
7G86nK7NObhQ9p5/uZRv1URQtjjNDyv4cP6rszXjMrbq/QAsmUjBA+PjxNBoj8S0
cPNkhMFXeT6MP8R5bNrfgj3an15bxDNep2jzlev1vbt+kxOJBTJqsJdF8mzG06tE
Jgw1Ve5MxoSoAif1KZy7uAv2fgNbwG/ndh36vtfq9lVyuKdLTDo5Hl9ipmeqB9eB
VvSrEL2iAQafPjAWfzFUD4pXYy6e1Oa0yxsvpXCFufsGDcohPU5k3yLSPyR5ZdPI
nswYjCxD+dJvYtb+3uEV/jcZGnERx/sYUBRkLWpxFd6IL/Gfsd3IdQdJAaSjiAEf
lSnIHcF/gNPHCtWghd9s1jE6O4WbQ9gkTnp2SxvNxS/EMdkxtLnxwqUYmQNaBV/L
Qblwc7s9G08qupDinTFFkoikl9OqkdjwWeuaxEwgURBl7nkAVDZrBFnTLwV5R2Q1
XeA705wiCZB2Xo/fx6IBCW99UkecCwMDtisGP46AufA0EQMn1QawMHGYcJHI7ITp
CzbHeUXzGdUBlZJxaccDHryRKJnREA8hMaRSrs9DVVMGPf7jVCLzyunqFOugMQ+u
FseHBlp+0/etNVX8oXRGt9sKV/32BkELtoAopBjwUR6Y4YHEI9TcwO3rMOceMVCt
U8tQFwvIjNHy48I6AZuKb4dV+BC3fj56nMqF5T5oRHLbdBdtesR11GqHAusYujO6
xOVRhJ6DdzZwvRKClwLGhuJpbj/M8m7GDyF79LxVZBx8D8SFXMi3jr06svj4k4JD
VRoq/LYWTaxP5uiXcfYhS7Skroh4C3RMezPyufVhsBmMGeTt7ux1xe6Ws23ZgaOZ
kswX8mvoy9BGjly5f/rbs8uxjLl/zCucDk1IX/C0FfG+zkUhSykaTYIARs3KOFyu
UQj7GNBEgXW6R7QeSiKamNhD5ltfn/e+Scd9DdGC+exd56zzDQxlP1feflbiB98G
xvYt65XiMX2c69IaGoGHMKwFMjnXpnyVnrXHAj3uP/WCpWy6gZx7QpUsPNUZ2w6S
i0jkhaPegjayZAFSwrKlGJNg+uzcoF2cSMtvdulzl5nrJQlWyVb72ZiTA3+ehrpC
Z+lEJHWWN3FawmpNImHVkadze+OqtjusnmyffUXMIDgNvyszwXZD/jjdfWMM8i0o
PQ1O0ncsGfaqNnvJtKNGb1o/4EkKTirxy3tRfo2zEsLQPX2Sz1ygC7gt9Y78XiTg
xJ8LwU0lSswCsd20xOiT4IrupmoxxrAuca3mryYmr6LPLtPOBcz2z+O2f460gy6R
AZ9hBj2VcyWJHTjGw6XIxAK6tWtBbGVNKxbQGkv7jpYRVQs/7m2GUGf5iNObXJ9N
t3SxPPpeHXX5PedSQmDohmWgahMYzZF0NcfGj4EN1UCtn0YfYCMwyP4ThRiRH/zz
/k+yyxA+bUWx1i55I9ajRXC6NopDLnm6jIDvF1UbSYhi7Md3Onq4XCFC5T4zOGil
ZthxpYw5WGHiWCv/fnNPCEbGOMWtAm443aqj0JIvF20=
`protect end_protected