`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 17840 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/9huKRhRMtvnNqb3Z+UU7TahEoHV+T8U3P3ufru7l1O
3DlgtZzb9QxCbOjthp9+wDkjygH0eUfDrEl1ovhZG60p+KlP1rqrt7ixBkHZjY5r
854TEQ4EnNlIJkCT7saMFrojXkLbTJk2ozDSwbKtbK1nag9D2R1/TbBJRhECYnJk
r//uDdrfP0o9zT9N+prQFl3Ztx7YFVw+NMfqQewfq8wsSLG/rSB9LV8if3urRfMw
FJMk1oq+saOuduUIFY8bQqZVYuAJlzfWrKKvKdCWM6x23X3bYdk4RcN0nlPsk+uK
dxTuVCqN9k7zdidZi5PJjRmEQnFP8oS1DL4raQZvWjL/2cXL4v8IHkaYwY7mf7zr
Gw/y56H5fLIXgcqmyrIvy2nipp6iOKKOfXrC1PV6yNu+GKqxcs8PNF4Y9uVhseD5
s/vtpQnxZKAOKPM+wj7OSoD2fSbaDL/uZs89ceyA80UYej/aH8M3XpQA5z3g2F6a
4ZCH7BD+Bp35W1snPOfpKG20VZUv8Gedv5m2A71ycIMfDWeAexPblvX0YtcHfXgL
QLJ9Me+IW2DNJhOnMS93mzs7QTgDyRpGUl61X1kDwLFnGlamNzidu9AhQs6Wu2BU
6LPqiaAgpqZiHk/B/wB8GdPjtCpMuCblz6gX2CyCcqADdLjIZNaVU/zd2aa+bTRf
t3QzquZA+SQO6OnEftT8ZGQxa0fZVbJjKTDD1ovULofFThBd01MrJdiFUgIwW90o
9gaqPA91bCBPEvCWx/g6a/wd/XJZNicL6TFScJlvUy4epwvH2BR6NK1szZ6vT1Fz
gvMpjUQ04jR/7VPZ/SYg47iiqPPzpRZJWZHZCWR1OgtPtatsWh8AQMMV0v9aYhhK
aNJX0dGtshznASGut4FElRraYR6L0obai5dr1kI00SxL9hxxSltpQdByOkoKUBq5
KnVGZjAiMg0zXcNkZoriJ2s1Az0eGlKa91vNXUxdihtPAmmeugDEmduWk28dzbgx
ECUcrdD5HQvOOvfTM/k6BMykIRzdc8nhOQIz7hg6OsUsdfNCxcOKKO9z0bUIY17Q
cXHB8CqVzHloVqNe+5dZlifL+GE1o9yW57YY/UIAt4bm1g1Z0AlxvPECa48S1G5R
DjIY8O7qzPbYt0hNL1hh0rOI4WOzkIFq/xmnKWcKDIVsiFVk9QabTd29/j0cK0Ll
F561QVOpASEYbO4x2Y+wn3SKhBOUVeYpIKY5WsdIJqGALdI7Ch8pmhjnQRJwyQIz
PDWGMQn3KtezgXNhY7YX+lFI7NmMtfD+r7S72IrtTcQJTOYV0AD+p3PKLl3QQH95
szGEm+PRBtaMrnp9OfBldLJEWstqPM8xk8cHSc1SfNx49AJxyWIRVZgg7VAnpq97
EwqcyWP3pZrmTZvLvAe0tZ7YT/3Xdk9qaHAvaNHX65PFYWYp0wXNw3pL8RER8xJz
6bc5JBLg6QJNJOV7MBuI9wr+kJONdEoeWu/eL8JP+KbgNj8U9fm/iv/EtMxk1NFR
Z+Tg2iDYTrRoUtHGBfTsNjo5aZtPk7Ku/x0WdsuOAjYDqJHwYrdy2lZmevU0jw30
LZ+j7D0CixCY/F3u4KLcwUbg/eu9q1J/iNXEAQZJqeIGAGrfEjfoiCGVzDwDAUmL
4Kiy4pYGOfessUOA4Yz0dmD1tzYYgcur3tiqZa28DEoIQlPoc5WOhZ3sEVI6UHee
7ThklgTmw5cJRa02zjbnf/mJmGYuurABx5+ppVn8TqHB0Y+zwU2d0LMT9I2MDLNO
KQAs3Mz1Butpbw/Hl9JaxB0iKD1RZ8zFsyiVQnllCmc2KQw7FU1bkQfZLbyTuxhM
F5BFOXStLhkgA8VeP4rQVBBptO572D58ocQFM42Sg2gAKtZqpPjzkzBfr5kWpHpI
C/S/8IPLATpazpP6S393srKHz9lEwATEj00qU03ozTHTbdvynmQfebar8s2JvGim
l8HRpCu7HvRCE86eVbvGcmTkQ6n0/ZDMSr3+O3ZjL3uTSPXWHeT7J5UBRhPLkpmg
b3W4CIYFNsNcdD4fD83q2svSk7dGpK8z1sm1dxUl81Bj/zFU2XyfRCHOVQljQ8o1
r55+io+mVUzaii0nPDaN7mSDLo7aLWOShm3zC6AvsRGr9pjJ8jgRf9TYwp9S0lLk
yPfHtMOk4YL9kkCzEno6LkyVyZ0v0W/FAePxkNa2NwwnTiA/NPYDZwEnoHox+t8B
XxiQirDW8yikLV+MabxQZiTa/jOGqHQk/esu0h2/LxaHghkRtHIecnpM1zE7oo9O
qjNBnGrpNP7SpdIo++TPhV+Za+6un/spiyWII4LSjeFKT22pFhQPRFOcaHdVfEx1
vz2SWz2gXjdPiHKssh/ZBADvASvDSdWDFdz2mxhh/KHMtp8eiQqlmAijMzNJgSPy
fz7J56nDL0p1GYNZqpIpCtx/p7RsZIHdFWEzjQ8Q0iwjgOb69s3V3NrCfk5GPEwb
cnd/VTp7yx2OjKV2Hxg8jv+PC3BqYYC8KKTnkCPejcbuvLLhHN4yQ5NrNk7LbYnV
4sTJWB1jiOaA5n8Q6tjNgWm8rlOl9M9htUokYAz4xt7xp0sFIFOLXCIDKR1VoqIv
Q5DtasiM5D6YCS1z01N+a4NFDlJQ0tWh4odReo+FRB6dkQHLT624Vi+3Wprjp4ZZ
SGOeLnYh6EtsKQLJXtVrpyZEf/6Mua6rjAncbj/RklapenF6JYGab5OspW0HMYH9
HWHXaiRjy6SL3/0o348gP0wGV2N7THnpFn2C6F2NxTep2cIUvNv9xL7020gfW42a
qwnrfr5Mq8vgWaWURhZ1J5PUWolxoBADKnIGDpRc10JZglbYspsefJ2IoZNmSn0a
Rs2TXtsRHguHMJf8neU3wd+40TUkhC08aZ+0lmAEP2UnUR9xmsXjnlWVh+FF+87w
Sjd2dX7AixIFo+F621hXIqoM2KgFq82l+tVmqDlaFAAgEAZjofzVRjQR8LwuC5d6
c2WgUn0Nmmj8DfyCZQHvUgTk2pPrWp87hQe7ejNRbX1ZTgLHuY1fTfUHiE89jdgU
4Yu2aeVuH0Ylh7AFjxPHxZ/uEoEMHWv3UuI+Yw7rm7eOI24NEF8hfSsMuCbFeijt
nbmW+2+wNto5CSS2NgDR8TFFoQPT0/98Ld9uhl6fT0Z2pTHt5t+etIELlwTgf6oC
vGr0lTCeRfKVb5F16iTl5Gg67lOCaLq1HvvfXFpWuOl6Yacrc0Nan6e5kHN8mxe9
91LobCYixQD3nIW8d/GBHTfT81ya1rZV8/UVq/MSdDFIRuarrwWUpGpIwRo9wpq+
eRM48vr9++xamOs1kSl3tgvTxpCv4Z3tv89lRVmqo7O9P0dTUiioYhwKUUF3ymcP
inwWZfQbZLn+Ryv9RI4nOCZ7UFRSapSzChiPuProJo2NzY+lMYWYIWwWJl16+x/5
LPujZG6XgOVPZ/WQnzm/3bzsk+dtwg3np7xUET3UzzHL7T5acnUr9lw7LGsIUlYL
yr30SRZkujcSI4LjbEq9W8roC0RNAg6cz0PxolJQm906LPdHd+4fLjAl5rtOgudD
X8ssa0CkBgNHPFUz5edooXROevayTYuq1nC3TqOFLHwSDkwk6fjhQ907D6ZA5Qik
Piv/D+D9YR9bsnTjjKzgqrLjKrZRtaMP6QByrQLK6hK97gnBUyM5VIbSp7HmsBY7
Yn6CurNcaoK3jcuYhIiAvMg+bJObVGG8gnQCY0jRo9fNy38Obk7oLSUVVsr7+fPv
IL6pT78FNkNYKCDA43OLpxOzEve2qaz3WBs4jeY1J4sZuW20laYTTgzReH++20dH
7wcuEbpunA5pSlUzGuLxGjEPmfvIsSv9VYyawj21Re49zXybc9Ud6RTatwy/Yf/e
Dc/Viy3sGBVnlNtwUZnVGmAtB/6n/GzeNtRGSnygJH2XXBsdsMwO4wB6QKubitHz
OCKtEhAt1mKMPyqh+EhG1TjV9GeYywolekRkOBQXB4XHpYD1pQAN1r7XUP462azT
n0XG0ax3mOcjW6kT9ih7m49NQxxgRNqSe9mZXRIrwlSUZ5VAHTYs33zrkVpHCVwM
f2BgNs6BfVsaqQQkbLlJtt71LX5HxUkoFKRPYCnkdHia1W/xFWb6KgL+YzLaNqZA
5BJ0U4/2D8d1FH3TT2q1NMmkQ7Y7/UuvWIg3IHsKwRXJfS8/qhsQLAmE6UsdTxUb
UFTzv0tSu6EYXR9SqTNesOnDt44YqRnl/AwI71u+VpaAMlTEZsACLBce+0AXMRKg
asKbUSHwseLVzbUCLgudqPJOZAJciytWOeKzbiN07ZhHNXsYWu40P3zjosjBhfaS
bJfD+LDn+YJRVDknHmw6rJx7wz20pDH0LPM1XgVGNBoFYVzfhAzMoYd3VYqdgd6V
sL8Zg5B6STNzqOQggYhUqnJfJhlfuhnZW962CV32FyK2GxwupVyp11taPljcPmGT
RDJK0b+seoXDMd/xbH0XGR02ktuoTvdVUU/XUKT6jj+6DvUgbaDSrL02eKhxwMiI
OK99lRub/p6oYy2IYrlmJ7R3U4Ai8X66QqEblFgIEAo5uWCPekThLW6ZdqtDydi3
ONhaWMr3sR3saB/OwMkLhc2Y0LDSjWwxxJ+bVTOabGHKUKsrO5LW+W5F6YxJJ3nf
kZIelZ2ZPciwUBFZmoH06l2VOdDTo3XJEktir2MEu+qMSscfLaZGEOrERLxvgr2C
YUreM14dP3XGxMEMDDVN/vNkDe43zucyFWQTd7VSXFDjr0v+oqKDsnxmAXM192FL
vBhVZbbtoGsWYgQWLlAU37Yj1S19tEoHCjkxoBn5A/XAHHeTggsQ+kWAnlZusmlw
N45Zv5gIk32xBoqFqxR7po5mfrZZE4Kiw+Gt3NLqKMrKloIqQB98ITT0ggJyc4V2
jaaPKjEqe0WM2IDF/xzkJtViC4YrvvHYHQW1Mu7oM2GMn5U3MmNnSVocRPh7b2If
KZQREI8Osj32F7rtOxXYC8Nji73e7ePesw1Y88NqD61ed/AZcBlvsz/kGbbkbOMC
kk9RlC/HxN9Ktj8+oXGw7sZpT33CPoWf7e8T+A7XL2s/02kvzUlaXr6i7Ipa+r0/
SBS0oOb6oGRz0sRI+nBE+EM99YVkmhvke/iUHDJs0d+u800c/hO5RJHu7fbSan1j
XWMeKzUvLeOEIqnTbnSyX9oDBIJFf/KbhvRq8MerzQ3dzvzGbgR0JYIcYA8Mx3zn
UCCx1d5bhig2QZzkW93S7CEiBODrC7gxA/P7PruTakm6CJ/vRoaKscDqAuEct6bS
Q3mvT8bC3pEjfUsqfaBW/GqbYmDoi2qz6QroP6XSXIviRL/RDPmgNAdhBNsLr1Z2
LHaDKljPZW9yHzvYuvrEgQSXA6wqcEytRdxkgrbvcmmbcEJyL8Hc8ceb1Cuy4u7H
cA1kwBzlJWYnv4Ys8NOIEXkwtD3FgKRBVdhdAlVC0kz+QEf8a35Kb+qSEUNTOUuM
WPb59Ds92r7ewOLp2GYXB5tzevEwExdt2N7YnxPhQz7HuiDV3L/dGuc0BURKniRb
9JPs66s3B1MTtG03Ov8LLCNiUwaJlcIvbT1Y7Nm5hpXkDHAsSdXN6/MY7C+EFtN4
3iAep3VVpmD4jbRqsWbouqFBr4+mPfVo6SngmPSFFpQiP2WCVr5ls97f9WxcX8cK
rwYb5mAOKJBQ0tm9OMeIYJAQ4actTNYJ/m2vDaffBg+EepOb7729cQp4bo3pUOH7
PuOA5G5OemCKRrBGIZ7wfMvKLRQ4ejMDFTHE9l/0kRvoy1oMcZT0983Oc3pER0Sw
tUGaSwA3sRfalJOq/r5QycqIrClaJJ06Yf6R3hc+2r1+vTS1LYQuWkJTO8CUXCsr
XLP6dilzojWRksIpfEWzCmGARrcOZh+rbMS8RKJ+dlQ9Ga9g7oxVE3E1ZboPfNKq
HHiaLcnfIT+4Um9ip2vz1AwTU7GpGWjc5Xbp1/c2Qy9X/ITZymrS5T76fVp44O/b
2+1AS4UxJaIStRdnsUyZrm7tYB1dj89zLKLil4U/iGJGBRmJBpQTKJVMTsd0OkE4
oBKZOdsJei35AG/nb7yQ9lDjrxANyuov+CAyrb/c3N+x52weIS5g3bipgMj5ScRx
s5WbNB+QMVt1tpG2B+34DSTvHxEOLi1pJkTgN0IFku/Ee1pbb5dbNlNdR/OJ7/rL
OIUs1doErILmo/nGFLXCnHPSvWou3T7GPJtyIOhi3naV7u7crPArScbd2vv6+oji
jSk7xzCaPcpGggcJNGrS8hPjk3zWvJTCTHJpox032bAX2pEa3bI2y1CzYXXLC6t0
++yThGqPyWvj1E3PvvZBZDExFyp7otIup0VmQA1rHPyHo1GqF0qwJ41TKMrVHpv8
qeDYMeVFhIY01KEqYpszMUtE+ruEh6ovzx+ShbByxZwxIgjy7F7iVymRh/aIQPr4
Bpr/MG6UWFYXMTUwUKIcwmT6TDdKLgcgLQr2eVMaDM2xtPMHRCqleWN9QOauhky4
AgTMCf9/tZ8/LQyvJMKiFMdQNA1737PTzi86C9IqXAOS39gP5dmvVFxzv3hmayjz
eQtFhYjzPPMeNcRFUpDwpaO4kJw0BOob03m7EWRQON0CKMjFRDKShLRsnX08rVUi
7Vk9NJYgO1rtJ93gvL81lWZJ2JWeiUj63fmzigb1+cY7oPmF01Y6wJtbAyNRCx6K
aFe9HjU9gQwR/8+a9kGJUCfch1gW6kipzOEaJkfgcaItFCaVm/pZi8ADIE9GSbPC
yBlvLKkjkQatwT09eJcNPO1Il5NgChPQd7o6RE9O8YQToSBM19fnKkH2XGhh0Nzh
73ZDT8bJsjnpwCC6j6mrhXyxnh/wItq4DRqYFWfrzehoNRnmw8XpmuY8fpfPqD+E
C3fQV1IcRWjYCmSdywjQc06G+SIlwTmuZ2GyIIVAoTDUfPKg6T9rx8EP8LJBJCIR
E49ECpDJureOHNQQPvTMFEm906nQgr+viD7DoFlARvMVabBcaK6o20xUw1TSs4GI
r0vKLU3wlljoXNxXbdqycDByD7qmEmT99QZM3Vd2xt30622fANj9iJxnVKrctNo5
+QFgDAHUnu8wL0k8o+5EwM8YrA7FrV02K0ZUIPS7juIS+m0owiaLZiBEeN0lQow6
g0lyl9NSBet/XfLagW7hy0DByTsxMVzrS0IMbDRlVykgYWU+f+lrShqJIFv6S7e1
iYiOGkclLEiqUgECbs6BmRLO8lZHyAUu12A6af9FGYjbpAlNHpT0DPvcmRrBN0QK
r2BmfEc04+OgqaEzHxnKQIC9dwpM4CX2A6hVuikmmwmIERJ/rGOiA/8bsM9dNKjU
66VfJFQMUg+euTwDKfioAH1CgIMZqflq9HPtKXz6Jiw2y+h3lpQeCYzx5s2opXuG
R6wqwTDl7I1Z1SRHJWnjYgFiyGlpwpk5RCxN2JiHJh3k2yA8EsRa6iNUq9K+8t7n
eszVhpq9KqVmWfaXArSQU4Nf+cvNcpq8/pM4H6qrldbURHuZno8KC3BfLtX8EgY4
7ndJyMbz4+gVBTrq0MNIo/bKZel7xlX27RzJ/mWfz2Gx90bUHGeEQHIHN+DvRJCr
v0OFcOP1lop9QCHJ7Un8BbVKpHacdGEzi+I5DtL840YpllCkg3NFxChL3LG+opZL
BgPg704K8CI9P16znP0TCptM8TOuQJHIQ2Zi+mzGw6euBsGHHTpmQJ638Yh2wZzq
LE9qRhFhJk3+XczyAjvU+PqF2VQSiR+/KhMVUmnDTFkdYlQGbIMeyT+lQrFuaI4q
GCB64cMqNt9w8HcaOGohJ61Py/4wB/pSU5Q1I5j/umfV/j6erbfUvMVisiPD85QO
B5fHmw7q2yp21qMntxVN3nCo55+Ra54Q24yNnEbMrG1Dt+LZ995Up35bg+XAaB4Y
ipYQV/PEl8LwIdcDtQ+XmFZShqF6kXR5zBlo9N3uTYJXVqwK98YQeFhC0ei+sKXz
GAKhjdSGB3bm+OFMHyJ2ikISlw3TfIITkJM3oN5VcPoOJEK42MhmGOwk3Jbo7itd
UFRFYWNX5P/fnP/El+M/De2/QkxpOqJWLVVAP1GjeWwg3p69xF6I7id6mrAJR7vz
Zl5+OW7advdV4+D9zLB8x937q2IbpngdAJHTSX2vEVDhuhESuCfm+KzdEj9mmWQV
M0EFEJpSdYqKqCWQrLEHzETC0d4l1wtfxi6bsTkd6KC4fWchWN28tu90UoJ0howf
zp/L28rrm0kIIQmgTQ3F+EHA2Wxrfnn/pSEaKIbS08FqrZehx9Sz/r88UbJ4TrzJ
m2XO6unyAN78c1n/u4Vv9gm3nhZDPovUFVLbm2c0NfzotlVUUw4gicdCbSBaBsmI
EcbJ8mlaARybbcMyusPzUVHTVjZrEC7QZxx2SUMpe9NsL//3MK1XtnTUiqZntya+
zkN03IhhbJDeOGo5/IaEUV3SfV7R/dovq3FiLog0fz9c1e5NQhcaSIkY/9TD6OIJ
OHzCv6+/IJMmoXOzdVclQmG81dklpCGG1HqDpZ0sAOiVoXZcrP2aHngL+9BSgeFf
2QyGAi6A6vgXQ2Ukg9QFh57D8obv5p5amKAaVoiFcQcoD8csHIqLj36m29dL3LsX
Rf708gtsyHxCdB80hq733AyW6+PT0Qi0tVbDi1crrIRzRiARnXwTbYtnHePPxK7C
lG8dB0ZoCMKpkPlhGDlGd+HusM4YxhwrHLRADltegs3ZDny6dsGw5Q0JkMH+alS2
Z1P8qBCFlZVxGGQUPU7ygP/+jV4bEt5jYVeWNm9PYwVaUX6wW460tPTT/JBkw12r
sv3quF2I5rXJgKcJR/fLiHUg8VxBvrSEG+aors4UnMS4tCpBNvidpJUVoiN+gH6b
iNXf/sg4pBQztwrPv80nLtU8KrALnLs9Lne68ZbKaeI1ZS7k9zGFuSuQwh3hrW1E
V3STrbEfML7hLleV78YGU1gMjwr6ucr3hWNuq3+hjCEDjv/WW2qPY78vCYDcP5Vv
DA9ZddQu7P7L5TQSrVZ/j1U6G1EuwWBTRs2rWsKmAGzYqEF3roltmAW1xAZIXEs+
hVWCNCYB6pbBZlzpFLAoWPoVS5k4wVpI4ZTtrZYNbxkF9IjHdbvRzZZy3YwKPLBD
U4cojYEV9YweiDaLPfhvBsRfTDScUrEfMHnK4+tNZVmjOZLNBs2dP6xsjQrJ55md
AyFO45v76Ji7YBPmIB0PhMu13BcGd+az4LwNrZHkTlmaHDrRFi6sOWaLxaNFk11u
oWxO4j56IvHv0pMbi5byJlFWq28te94P35HR7I8lNWvMWp6Ru2p7T/kOg6kBlh36
nTgt+0WgXP3KYC/zI2HEVbqYeWrNTDtV2oqoikCqdrcUgLh5qZORkubSG3jLbi8i
Ix7jwyZ82DsEpvEKbqchudQdzR/oRuwgWjBGsSi0ZcxnU4OxXMmtIqxk8s9WbjwM
2uA2I4ufAPzoDxstoCZ1n6Km88F6P86mTSKqt7yJ62KUUZPrVGZ1PQkauDRvgytI
Fj7e4hX8cgeeZi8L+xcVYONoIrQeomXUsJb0hEaNe9KsgQySKQDLmk7GruQrW6PJ
u3x3K5pb8Ls8/2CxBYlzTxiLI3L26mxsdf+dneiVGF+3nJRgVYjuM9d/kTx7RBj/
9/c79vNlBDsbVIiTaJ0Hhb8jnGZf5N65TJCcU7+XBLfichBkF/RJyYu4901+upKj
Lbj3rZgCZSXLyPKMGGE/wL5WBzij54Q4JhVMHQzBMM8YwrZMQpYkwI7hEhi17/vx
FT3pXXlWMRE8BmZ89jri5C/CPps0YJnJGd9kT3OwWRhswZIaOFyGpUsgiK0WPqXw
hNygTCUY34oq5zVp4xFa1+l/Fel8JCL7lnrLvZQPPngoKUwqLwJbf68P9cE6bXQv
QdiqjcDGAXxfv0QPmAhzinvvcNmhv/MPua/PcpqimPbDqraJ5hAp/1Jd2VoFC6HR
MWiDxrPGUE+g1KobjwDu2RC8gWQ5UTxJoch3BQQz9AHcHsSSOgSf/Z58yQOHXPAw
gSfIuX8L70DaGu9uadl7NYFD7yqyiiSPYnK/DnLVYnEnc5E4ih3nPHPCOiKhpcPJ
o7hrEAg/CT2OXY/CrrdEkFkZZGxiIAisiG1di97PjtGwvXhr6BpfexrsBYsoAM8h
0hOM1a2EVJZPfIeSoSRnbtqiJvDggrDyYtzEZ/VWCkPDD3yVpYV23z5BVCcLPVYl
FfS4gmKikeOOtlgMiWLrFcK3/ucCu+KMRwZ6APwxxHuL8p7kzlfRwZT4BrBQvIzr
btPZxZurQyOMJshQsrGAXIoJ4U6k8wXARkpxSghM/DS3EvQdAwyNRuO+mY6TA1JA
4n7YLaTkTBrRu58U72pC5s8gHmKb+U2f63IiQ0sMvoMs3uchSymnM83kNgKsuDJj
/hufMjJCkDzYRUMyFYg3ar8YA7rVzNaCu4ldspdA4ctsaiNYIG7BslQPgzieB3da
5mlZoNaNJW95sgIXARG1nvznIm58kNyC5cy0q3q3F4Nf3xAdEyBPdtFPuowsZFp8
oC2Fo/Xc3lbbakg+Iyduj++HKtgOgKSZ79ngpqPB/Wno3l9FQb7rXTxKNIuUVR21
Kldk75md/xZ84vsu7DF/lVL1WgOJW6Eq0XUaKlZ2Nogc84ozAYPqDzzCd3+pIiNr
OTaq+0O02KPHF5Q79IpQ2IIk7vTyqv3Wh0rSeNMilBK0LJFRn7wGza5mqD/WzNOf
HY5Yiil82y5uCu50G3JsQ2b31TKKTuKVop9st6Li82gpTq0wKWPhOU7r+Ye9eSxa
342U1U8IPEMqvhjPAb5jZKB5dX0RitGw18iKnQn1hhhy9ERbpDxxyMyOrty3Dj+j
80C+AcVJ8r+/9eTKar9+hSx/jbfDP4CQmcJhraYVS9XktTJQakjq60+qRLZDOjDJ
ZzwH5pU97yfjP21rpD3Z4Vo1ubAFSY35kqfTb75a3kouUMA3yjY0SsihQ3JUko26
bA8+rtf5zrT0NBA9sB9GIYCDA5Thv5296Py/feG7ZOwTBnC/Ob0+VMchBVB8njEd
QRX2Suygj20HLVkFtU8eUBMEq/SQafaw6yhyQhefIJ/aPUgxeFQBV8eS8jxM1adw
OdGvzBGkDyPwxCThsGSzmE0jKjjkb3VdmV8c92Ms9nWIPIK9Zyrq/LPO0jZBzk1G
MdTcXe/meKdfFnU9mQyz1zCMXAxLUjLyMmTcFccAewcTHLg/cGc2bXxmc6/OKliU
K+XDKBdoXEs9PeXIZdASq8Qj+CPYEU80sKw05sWQBpBf7mFchSaXDA9J3DOcHRQn
EaHCjhHlP9/3Z7K3iC+rHpdKWxX7XN09GDlaO1xFRytvxmSYV47xP/Xh51ljFuMh
u7WPd0OXGIQjblSJTPlTA0piIHc1VuD/MCQxsBWzzMOjY/AVzv1UmygPNZKvmI1h
r1zmHB2NmGydwI1kkvwsY1BGQ0D5bFCe5JbZh87hNhAA9hD2qy9/tMCd8zG24z0e
jhwHmhd0bJrlpdiABFyHx2pYYor2uoOfoXPNOdezY8bDBOufTd8Kr7GT0UlyrANS
Ma3Ty6BHUfTXRCaSjP4VJ9rHlUkUqAMHXxUZH1AexZmsXLy9ooWrlCkFYqHh2iAp
HNXYGEDX3zSBKis4V+BfgF3ApSYfZhOfaUdR5cMNKnFn+R2ruAcUo5JcPqAcKpgh
XCewh6KscO4GnwruxLaHlKOUm7RbnRpCdBvRRLLoW8HOU/b7AlOEDlcyXnaK9/Xy
kmv3r/Woc226FCccrOm1AD6BJ6MwkDYmgfMQPHBQjzl6SZB7hnPTslvzqu0JIFVr
/asRdh+UVJmx+Ku+daSsMUwTPRz2/8hArQQHFXn1A8N7QA1+OHxq14HTYFgPG8n7
9e/KVIz1uQppvbGpMXZqvYrf7AoHSF9bYjkB7xOKmIN/p6H5fwnT7i4p62RHl+qj
Nza61sI4j8Ozl2LZ1J9t58Vcv4/T8eyFD+MabiY9CSFYYT2jub5OKTKkRz+dVxvs
Sep1OVHxU8ExjxT5NrSkqbAvRdBdCDiwCHKzXjsw3si1xzmZSGh6AHcDfx7qYyJU
WTikxfvWB03NzZqc7kpTQ81dLyOUJSFth1W15+MNykdOpGXkec3SHF5rtFhe1hG4
7ZQsKkO6SiK/Gu0d4IV/VK9zUtWWefN+IY3v+XqpSHMllF/s48Nx1+A74JZuZOye
nTuFZgPk/kxq94fBphu4SJliRJSOmrAH/DWD2mkNEnJ0KXodOVislaVWfY/ENayG
UyxQB6Jd+zhpTmk8PCr+i/2XGEhfwdco42mP+XELqqy36gHKVwRmRIhmtD/FixXj
YKo6FRFUVaTceAWyD1S9E09RhmD6n3a0BaxsdTRJPAJpPd302L0KWR41c9+xzIih
DPvG4O0k/SV5A+BTlzCGVeV/DCo3R08U+h0Ph6pGXYzmT2FGHufNatRpwAEqydbt
PLjMrt5Qd0MmI3RLR1WDAO94ULtA9T9XZqL+4nyukFAsxXrj14er2uRrQUp00M+u
shcSxpVWeYm73Ay9JXJ++FqnZWtxoezSlGqvyz2qiafwc0AdmhIqv4ABerScoWrt
8zEyWgbCAl2mkE89Qk9KkQiunYBcdP02JDwbhUQXRI8q4JSqL+On402wywSMH4PX
7T5ceJvIRdZL8jIKzyFl12YxYeb2QLXWeakOxpZVY/MyHPlhr6aq2RpBK3EZliys
kY7EW5ffV5Fzx0OKD7HjXpWLpDp19+TIuh46zPqI1vvEZE/rLTFnG3Rd5ZrBChzh
3XwcEzyVDerul7RNokQRcSzbvf/ECgngW3+NJpuoMdFPkrwIdJv7C42Wu9GV3Xzy
Pf652fxF9wlCwSkuxP7RjOhFWM9JoykohvG0uujWhlNlbkm2lV9V54RL1FpkX9Tr
a539mu2DGzF81yjgef9+QA/I4SFoHp2XMzD+j1VQb2Q9cdCcoaQwDWCRsLTut0aa
4yv8tqNGKIgHnve32qB+IpGzp4BGiQkg6B6EaudUhO5sQtdOWqocxa80hSQEZZxB
/C7Q5ZTIB8UN/vrBksQ9YyYcHwrYndiA11cZMLF8dNxDCoMwR6KLF1QOy95BuG3l
KLvGXCvXmy8kWGzWpdmrBqOOnialRiqsmLxPnEsafO+iq8syvyTK5+aau2l3P9hm
Yljlk2Im+AdxNcfxPSwg8qZj3Nahxu5FUNZzdWyW5fNf5wyAyeF4UCasOuu/htTj
SrbMAVPEDHMYJhEHJJMPoaAmctnkWW1mPvKYR4D9ekt0J1ELRUGFxLga5JV2c97M
wA9nbOr4HaTZQQxolQCg3Al0nl2LuTcS/XDecWKwGOn0/70JOo/mHm17xgOyTkC0
D1C9GGSuPXztZtuDDRQitBnW7Srt0NqOkecXtesk7v5bm0rmdeCvjBH0RX5RjZxL
x2LrbfJBlh1DxkWeYDQh4aRoJSu5ATWNHy7d7nuS3r5CaiEMRC0nYD8+aFpsI7cE
bfzcs82TlVLW9qnf3aLKqq55mqNv44zo8MfpJHiKJUh7LhbAJSQHw9UlBJV4eqjO
2NoK2Teg4qUQYEquIsnq7ZQoTr4+kV/bSXiwlPxMu1oy/GLqSgrlJXyqpf1VmUwZ
qLsoOjZDqXnLfnraVFHGkXR0WlLxeqHJUCtzc8viPaeMELbXDe0jFIHKn9dNM2sY
qnlFi0kH/yQD5VG6dfRK56v7A7rV3TeH/zlqFunNc+vOLLfsjI6/g7FAtl/55baF
kMg0kUnoGcARAWFgotF2Bfv3qtjosoGlle8zMphbxCQkJZdfaHZpvugSAmmNUQ4i
2yiba7g7TKdPKggO748cecZ42FmdwPcV/62LyWZo+HyC7NNvAvskZF//w+daZwsj
LTQyOcOOfbLSDfRJF3xzir+2kT80xjK2MpXFcHOO3ydMWMXj1xSPxUHJgVRSUU5/
m9wJRyDu9VaEGmdOwtRNsAn6EjDj171NGT8NEYARR3jJln+x7Mbqxj8ZX6uWPDDN
s+fKXtWCxIUaP5Yc/EZuMnQ78LKZuo0Jkv8zkG8jKc7d7JtN814hmVGuZT9KKpUo
GMUCd0MYZk3Gmvf1gywSgjebvMjS7pQGVc/Zbm3Q0ccQeP5ZNwOhoGPHZaUN6o4H
zqLPkd9W3fOY9iai9lHDaahN7MfeIsGYdwRgYNLnojJt9rqukIxWMDjw7+/8U+oD
4vcDkUawY0I27uVxF4WSsvj/em1mDikEhjtIPvPJkdV5q94+PhY1+nrDPMMKDyqm
AK46QG0W/AQ+gLkZPuhoS6DqWxcZbZ8QWaH6AmFuNxMph4Vusi60pi9EmviQAe0Z
cn7pkH5x9yCcK6pvIDTNET88lW9UcN4sQP7B98k6EywEpA0LJ4oCiYaVzEuaCT8L
1nKmYgW7htDcT0r5QPr9MA0PAD0e+Rcx1dpRUkuOjphBazYBhZfrgV3qq/hSiMZh
uvdiss99Qa+kPWxH1OGPRUWTvGuXwmSE46+v5uyeX6YatsqSvyPOWgZOZtBhzQoM
XTKpqH/8V6786houoNz9y4Yi31v34+gocawuBLKU+SXSyHQcGYg2xfuM/INABzHH
NXehhJ6XiNI8Ny3mECs9mpixxmhE/DoIqJ81qKrKGxexcS57fzYvg4flsf4hZGht
phSe7hs596ApMPrCvgD39KDwN5qMuf5bWoGNlFVtgAHIvjTdC5PtmZeXN03e1YK7
Pi5N9DyHxZBhqN3+qWYnuJ9Vit3hC0TYs/KmReHQZoSmEqKlpJHUTfLeKwqJCL93
0v9a0ExAyNfhMHe82fUVk11C/acqFrdKpkW984zcUJib5Aj2kIUU72kzhtAewjYo
2mCVD194lFoa10fAcZEsn21uLEyXoVtIJnRO4mDbWOLIET0bkLrjBvfR4T19LoWd
Qx6DSjX7HUgnjmOM7QPzAZEZkHxzq/7dKk+Nh+D0U9Kf+MBlwTbs+tlZsndtwsgF
arrSO3VHR2FhFCKbKYmRv48T+AKxJ4AECaOSx0MJu/YYsU14ILEvtP/zMIToDd2Q
QDfRF4ggf6/rcVldklphsHbI0LCVmJCLTyKPBw27VNelGjsK0zm06L57qfDaAnGD
sChHn7XPi92uxsNYAi9eUbYqn50nv7u04ZP87pEaeFG/c270Ryy17TcDTPF6Uoro
Cd4GDZP47n4VHviDrATIkhwSnZVfpfl3Rr24n0Z+LL6E/p080vJ50jDhfLjO/CzX
44py9FUYokAkr/5iqsqD2RojMRRROt+RdNOP/fs/m9GrK4QnvA+tem249IfLBLKk
QRAYwSPDR94u1lQp6v56blZWEAp3kotd0xG23OxOOpIGwYmC8wPj7dkqq3pAZGtF
MR+6YiAAYoYws7BMfb3uDee3kwjSZMdsCskTMrzc2QfFggeXiMht0yw3/Az2Vuv7
qiyhtUAINGi9uczI3mLscX+Il0IiWfjnVbnInemd2Yy0Cq3D0QWg+rtGtUtR4+3n
09ksgfjC5SyQ40ONPMyC+zGUF0KN9Tt9DOyrRDkocA2v7xwmCJxf4UyIwDc3BGrV
79JpX7FsFTh/7lWk5EzEHuElrLhvqw51utUwtwqf2BfBl7xM/ktuXkVlqnDTwK7Q
I463cdVxyDDm3QmONCOHjz1M0zr5Td4YfU92/y55CbBq5JWSwuhB2U4dybxZsgQC
mHI96es491T4dPTI9dvUogL4rqc11/iu59jkFgnhT3uRs18+30pkiIr5XUKLAdO+
MAcujl82itBVEmX35ZCW5u/n8PVMnUvSAIXdFT0rZxq9BRCPsFLjc7MtdgstWG1f
I5OmEQQTqkGPFT3q3cIunvmXSJR7xI32m3L/gF848V3DD4drecYdV2T1oGGy3Lui
wpnXwpIBuvcL58P14owP8qLFg5STUCfWhU7rpZFy9WMHLZr/HG94/EjC0EiFWglS
v4/SUzqqyJ7ONDVISv5eGYv6WbIjV6XuCVyosP8IRmUKOadt6P5d+eUG1tyBK62m
K8cCpQX3OmB/BxAZd3NMpQohPmg3wLc2TgR9kfrnxJyxIB8y1iCcH4E8wLfwubBm
do2pNrICTWjyHkwdgwa8kcqm7SH//xNWrdtwsSDlBKgiZZaczoAHjYqVgpW0+PB8
hJ9TJ+0q2oce1vNaFhBd3gt1cq0bk0ah83odkYgzcZuAhuqrhw+EiwDzYsrWDcLm
ya+x1KgNGCciyJXZtQDbG7OkUODfGiBKQG+R7YRAxjnpvfYSsg/IhJab8lpqIOq1
qigPxVpZFYtzLPZHRza/tSF+opshW9hwaXfmQ0aNFYGijiLieaOwqYVtuCHiV0mS
LtTSQehtlTzvQF8bydVsskhNe8yDdkyp08rCo2w9+4oubIp3cPzHQ6lisXjlv6Ds
lGXo/VUApCC0F+jqBViI9zEYcmA0YrMjchms5M3CaVndhx837hM9YQDdm2xR5wCT
AuYFYYaMddaWYu3b7Nfkq6Wp9+tQ3mUFCZALt6kS0bvt2SoAXCKyJMcy4HS3O2ai
jm3UpNTIbMU/z1BZMRd9ODVB5935rl92P842kvMD4IIPR148W/RDhku/t3e5Oevb
OepBhbrJ9iCwP+eQI+OLDnsaNDt/YUoxW90/vrY4iBhBEoF3kcdspRXK1Gvucis6
qqfFJosfEu32CzMTC5JhgPMNPBF5Kw7LJjLXNmqHTSLM3WePGwK0Th3S/ZybfRXm
TCU4tk1ECDyujWkRHbWfhSocF2eGwkbN+uSVakpjvcM4GC7By43BcFfNVVHUqyYI
piEVzf6a6/kZavJ+5V3zqNMOBjGDcNtQ1JEnz5KFMRe0AXjtvHdfD5jrINNCY2VL
d1Efw/li4AAssHYmccV+XWn3g7x0wNSpR7NR+8xDyTKqzZqbW6hBr/lESpbhuZbV
ltWaW66F4Cs+PJji1SAWIMDPdZrx8yACLq+9T8ZjmmNTeoAKq3W0/tNbj60O3i1M
9FhycFJwLfaUJ1MVUkXL5ThzZkF3+gNvtgVQljyLldcWFLpMo3vckbMHSVhySx4d
cBS9ntP909e+dRjuRsR2d6KoK+JE8Ji2jiwNG9SaPU+bH3S62GYn6P/UBmw5dsHL
rqyFKNLCzBldqTwXW1+cfdg1y6PMAv7ZH93oTx1bjhEXJiJS1nB8Ab/+6Bfq/0E8
cUSLmiACo9kdBv8PhiSTQ11qtWh5qolZhEQn6eI27FJMBHq17w7Hrg0dT6Kh7Vy7
uXV58vGdbp+FqkfuDTsl2W1DOTcEGfngWYnBKOqybC3c/2oZEqEA9DgRx5xt4QyA
Fk4PHBeITJsKFw6kDoL25lhmqsFihnOdNAP3i5SzWUj54BBil1minQCz+a8hlsUR
bxXOAiYhM4MTi3LuA+69EYDLrZM9/dMZ8RzRavxlEhC5a2pLy/AK+5okzh3OvGWh
iqjd3V9h4RcrMig0zrf6ZhPNRDd5iSNbVM35d1FnT0BrPrYLLwghZKVFu8YdAoHw
KwBZHaqeJz5JZC2xxvpBVvNhIcM1ceWxsuDrYkB8BSRFRgmKV86gWDIbJBUIVy1k
XrJCGz4O2Le+im6Tb4E4SWfAS+FEDrQaYZRY1jBlSU5KJueno++X1gNWgrW7wc3p
6RTNMIcwiVKJliMbipNoumdOZmP3IoHkN7ojsKai56H638xZC2dVL1s1z8TetN0H
ZDaCaOD+dixbf0MhXGkCPILkzWUxQnQCD4CK7ulPZE9hjYgopUxicylFkt46Xa0e
8FG+sNPR9gK4gq/P96vNf3YADTnfBXTR/8R7Lxx8QoHHst1LsrLtCNP9ne3pLNLR
kSj94ONzAEP9RYlQjrQqeAVjQ00d4kNWNwqR07T41qSWWJM7Mg5G25vvpkbCrc+P
IFiMkrH5eJU8CtNCO1wjooKf7iwAlAG90WJlfKdf1Iu4wAt4+GcDtB2Fmkpvl7IY
u+bRTFP1E8wLCiELuYesyHlhSedrL+3xCb1kwyWZp4dolu8PIz71/BB3utHthD7/
4reuRtP6cM67Ri8YdIry5ojREO4hmkU/wzZF223CF97xrfTGOpmPEvvqbVUfYHnF
eYkCWPU8+HlheLFVJbxEbKGv1VStByepA10Azm6EBx8itoklMW/T958fw0jvvV8h
a6xH5tdfzghOCIodxk5kr0dnFwhI9jGZRATwMcl5R1W3z3pTJk2BkRIoi/9MAONK
x+vzkUe2z/GC6FwS77dYfHb8JW6GeOi3WHoHQOsCh8AqTX9G9TSjamUIxHPmxi04
8ngt5jGwo9RISniNIwniT+j4hlYKXud1vUSoYU5othoSP7VfAT3MtVdnLhkDWnxU
v2ZFHfEFRRfuhXW1COuFnT7TFbPX5T2afm+Cj4sf+32bgSh6e2F2x/W+2CDd5Ik7
7tngZFmuASLjzOHdNmpnoKuTOXTAXFG7dqoTsUO0/vDXQjpsdoM2Tj/lqw6HzQfm
VNHeOrKF2eFcbgkPwcikSVvG3oFYdH6XeGZ1pWui0F6/8fV3P09Y+3Kph6TMhC0F
KguZHCieEGHHRdhZgunMac9G2u9L4+qtifGUQ7W0LpM6rzMuQ+B1aCjCQGUMcoIZ
wY3pJQWKvVO2FsdrTXDAVfl6Z0SToHuGliSsD+uWqON0FBK+8CVv3GXVN27bA1MV
CQiIp3ALV9MOhbmu27c/HXieo+ykfZIDa7tK7flzc+z/10V2ERrMiyCKhS5s5Sex
JjiBHMMBEzG0qYrWhE45gQzIvKQ+i7Itf92etBCGvPGDhmdBAki4bWmwuTMu2ScU
o4EnKKUMxzZo/bj5NOnYyzL+a218CM4ATgM11JfkPkIpMZO4siiYN7ScAbx9ke3X
QCMbsfK+ryoF/Mk7q4y5T9cIRRkbYBO0VyIXf+lhdmIp/6zfeZhmNwFzNT50TlpK
fQn/f2JGU152WRwLrIhz/0gYBqyuVQNHR/DNJLOVzDkrQx5toS5fUzoXCx2JFN0J
2jxSxOIS0gP856/jXrjrCgU3vayRDhyiWlq534bB32yQcl7JAmSY7E3isgKUn04h
QX2GQUMHfQLp1yxI5Ix4Z25vX7vRcN++I+SkTsFa0k0B5F3JJgI9Ebn/fKW+UQ/U
tKydBkVuAZIEMpqp7DdihAVFDdsfKm8/cFLavPjdFDKtONMDkiSnfnG5kR+UFHPv
O0eooxsSFREO0LHuVGAMrDIEblxN+c3UYZLuUgGx7V5XuWHqBBBR6YLxUhb+KDL7
SMUY2dZztDMsggivtu7LupeVpkiv00EAplCr22JCLIGmcll5Sboya4ZacY9L0L8o
/eicAywJ2OSN84Ynln3vKclmUMPG0Pz7ZKfNl8K3ntXW5MUx0Em1Haa9wiIweb0J
ZqZl3ozm5G0jszudeWcYxfF7aUSPdztvId28YZ6zCsU04KY1WaojKg6cT8FpBtM5
dkUtJyFm6Fixafn7GeyBz+2PSKNBdRSsNIHJYkl9a9XNv5SzAYE8nlI18jWHrEAA
HL0/HGSCXrFxqWXivk/4ix0mW6rQnWfatbWAOuJPyvuhLnkZ+5wq6OJcODD3zHtb
A76g6mWr5rJCk3o+31h6vh0/1Xp9wmVPMD1asbmpZFPysISn+gGqNLBsyfcUTruZ
XFBQ+H2gas1xQqH7Clldpp11WUc8dVYwZChHA3PJbdY/AwVR79QFFmnklsWH1b8c
hdb+zaWF26VvfbS4ygYf6Z8fW5RsXdqcWTfHgubYH4a3d3gzZWpnfoNcONo8r/Pk
x04jCAG6ogCw+wLNd0u7E4HBwFfySxjXZa8I5E29wUl+D5BNKEGoGVoIXcImgO3A
bX24y3wAal7cVuDCpSknhx4suMgeS/JufR6Uyx5igVvQ46bDzgcRypxXMfPVsxcl
3zIw8Cd5aJ37ycSVpP7c0ZXdASq1nU6n7t4TEin2VZ0QTTvTC2arjJukRwirfph5
0lzVbSaJX1PZku+bO69bwaMq9SF/M9QXhyd7cziXRdLiu+PgJ0lgy3WCDi9cVA7l
gr+V1MwyenvFonfiL4BCq8YiTZsuN3bTvCUdPRRUYQv1ZMspsuYINsRkO8VVhfmF
lGbm+3q03DbBn6uBWfdWO09FJxcUUnRshewWw3TN4nENrvURWMgHRImC6E7gNEBs
c09fOhlFjEBbl8ojlRdYoE75Fd7DTkgNsrj4Nl9gfYIIoxelE+G886Pndhlqm8sA
QDf+KpCT219SP6246xd2EjGtozq42KMfF1/QkkGq5JElCtZ94uF5uNGYHGEA4kRf
JwYI/MdpMews6yNG2d/Pxfx/I3dL/4yjX82Ov4U6LiNKRKHlmlF5rU6jKVCEYPxs
sOkr7ggIPKVR4+V8RMNo5OnzXO7/JuCt/c05DwvVPvik+kH4bCmFjIuhHtBmqL/6
lrdmysqe1phaGqUlfNlu3owO8w92/cDHRq25Wn2kdz9fdzCzhHsEYEq5EIME9J1m
xKTDXO87vy6LAajv2JyFb+Yjr3a4NQMpiXbGaFTTDBXY95PQ0UHYYrTMMBR2v0mN
QfEk0jcLiF8TUz8guVIK1g0hwc2Kszc6tby5g8QPlKFqihR9GkHwq3eFbW3uMW6x
dcf22zc1J/xWk4nuJ61QV/GWOT3/GfDvW67nWp7v9aKmKv0Q4d0dmgTX1a6AxY3P
udt3Hxn/1frSIXY5pWo5r18rPix59wBYIttp9XAGZGsvXoj77vWOufJW0SX8A2z5
VT7STRTHU6OK15hGCb3YYSur/Ku+BiESEP694fdJQeHN7vS2LW4FfW2ZWUb6BGaY
oKaT6CZfIWTjYaM9js1c5M1RHM4pDd5lnZaxI+TOYEcDApuwqQ90dMlnywCvmCmS
hYWrxcEK9fSIb2BeTAwxQvC8cZ0n2V+ZE1Cu5Jzp0JXGChVd85131ZiV2iUqJcbD
SsYQrtCKZbefUbDbXIL+otegpps73chSmexc5jVUnp79tRqPgDQ30iXqvm+iaEzV
Q3pR+Mrnjzke7fQT3gFLTiMRUO3dInhKd9bRTpGuXOEuSvfuOCfteUbqsRnPV47x
508AUm4HWfVCo9okydi7GnMXLc1WfR0JG5uUW1iyv5NLNGze7GAy0EVN8b09Q5YE
CoRdUXvu/qO4vVfWQ9bYeYUNaw3EANuj+V0zvoCxXM0XgxPlrx/S8g+uZpd41Xgo
CKvY+soCeidhpnzcAHery98q8mLG5+3vXFIxsEH6Ft3Qgvn6bn34pX1xEsJPCqjC
ZjGirYu4huqbBg4HlOjUr2G6gPeb8/qb4iERX+25zj/t3uFTckWn4NNDULjy9B5S
tRdig0/WxVC4WjMGlgNQJDWCjYnlnQ/W82irSAb0qS/cNnXpeRkkta6zsp7Pfy4C
EIanPFi/EDoRSgS8DG5vB/e8hnVVWje7VUbo0SY3bsj9qb/whE7YoP+rQaVyx9Ny
gHKIBEauXiM+Rk9SVXbYD07Utzd0P0m/CiWZq1hLHwoW9ESrwf7TXua9WWderTuj
uYowSNgKKWnPZiAn9BJsApxXyp4kmkEYuj+bk+U6sj5N01BH5/JlUhPTrgG1LAzd
p8JGDGHG3e8ubQm/zOZtKPVHDZu8c3XhMaJZkUMMSXMOML7LXi0a0+2QrEmi06/c
TEGRSUfLtyDMSd9WWQCICNV7L4Fbytm7SgBwHeBkQ07PbRfzbTxCC2XMQZ9khjAt
DE7o7osr3cRtECSGIhcb0ma52tLZsJJzeTMPMybWTppwvu1G8FR+H9vigw8zQgQq
bKJVF7iwyUj8RRbyjxF7oFNYjArLWm9YOWCzoQG+4s5xE8T3oz6/FoqXHrRh9WqW
OJKz/yS2wmqHzPbIZ6WwpRtoCVND/wQBrxLBv4oC/Cfod6xZqvH2zXd2dgs9lLDJ
9flqtTCR9GU6z7GfORzi7bv457X56kvGIecblOm9ORaL55Xu16GowungyM5y9ahj
UWrM3hjlcnxBOph8+9IsnYnT9Cozxv8Woc8EKk+46PUTiPFCjrM1BuiCHTJYTX4r
79MTC2eto6LRiv4jIoCm7PXKMVnx5W+o49YOK0z+GJY0ikW+S9eO4d3beYro1m4c
mXbEaC+syOI3N0xoiVWntqc7Ouq5avnCekJY1kcFRw+y2QaRkp5lkor0QavSj7nu
/Svh/gzpT2I2Nfwroe7cL3uovBvrWxgrcUkdKN3FifoGKsEcoKwZbeI9+OZlCFHg
0S5y6xulzPNAaxxUyZ/awKsnDWj+XpTBukTFUi23oCpsA+c8mNGjZmcCheyfjmIK
klN25M/WhtpC5aWBpdgJvJVPgieN66alV2oXtnGR8WPBYFe4irSl66GyBS1LRcqe
IPUki+p6ZP/8Oq6GocmpNYmfCASHH7LKkbeBY7iYI0SF3YnmKvRVLHEJ8cwhm1we
fR+IfqGBfCuzFAcZmBFgXkwgnlc475X5tKAFtJ80uQKDPDVppgWFeDz1r3SbVodC
EKwnlBNAbCQa06DS4jFSwoUHXy21vURpxViehZ2Blt2GpBs+nUb+D3bxGizGPlsC
FWTtlIT3CgVt6eAbeXEsjt5x51GHnU8r/TMIvWEpdEngUliSuZK/z1jehyei2AN5
WcXWWbYAssIlp1OAokBVwNVF3GWT0RBDKea7S3rCy36aJvcQ1PUz3YzkkIIcQd4Y
sjEbfkD5zt8+Qy06yakmCHEHAOvQR0y0sDEIi1WjW6OubWcQaBMkgYFahiHqr+sT
Dj+bomgUIUysx4vGjxwYOsbahMxrcARmIS9uS7IzwLKZN41DI2vMslaFpyYhPK+U
BcQsN/R0Nkgvh7o637aw48bG8qgfC55OA3d0n/z9VJEoVHGxwkQYCDeQQmDLaKBn
lDQKuPLNn0XnilL9WGDm2ppR2rN5vPBuRiDn9oPX4X+kO7Wo4jo3Ic6FnMUTU1TH
Qe96gCbx0o/iGiddALuY92EXZgzOnwDg15nlptVZY/zyIIfQVJcKobZIpJKK3zcO
bteOsovUgZMvkv4L+ph894C8bIJUdyijPqiozv92lrg2/jSUoR3HHRnaMP2p4x6e
4J4CdalPAKx2V6Iv+LXqrvTbE+0Pjxx4Y4tA88BWp6bx3qaPPaQ3RK+rYnu9SC8Q
q4MY9mPz+L48/J5Zd0jrxok4oygSETN7wK7L5bZ/skTG/DInMethlEfVy4W1qcKQ
fJJJ51yYNhMSamTYZzccVoolPh4ovKYE8oPxY/t2Snsds5PeCsDn60cpHWSXY7K5
7GG6so7ZGzd6clddw79VjM86oy9PBkw2yRhZSRnSup0eJoHrIAC147vhmj6TdF7m
8+WOK2sVT4T72OdiuCqXlo/TYPx2Coa1h24ZEdQ64bhWvqGJFCgnKRYiY5IAcCUS
7YZgGeXous2YsEmQm7JiZ4Yp7E5cewTWPeCVGJUcRJO1UEFiGhFrsI5j2fNwdFBD
lCE7f1t1qOCRRb2T/XNMo8n13fIw6dFgoyXvhvydMfhXn1Xzh41UM2LwGjVbfkA0
vP2LNeaIzKjLCLc8RMkSZV2Ujj8Ch/toXGf0NYUeBOz+hjF3ZyVMOm5i8/TQ13U3
GTHTfa4aZKMK7Qfz3syT3zlu/pp56b1rWOf4WzcfE4bFxwBm7uTPdhQXcfzha3tS
HugJoW2Y062N7Jp0mLtFA6Vu2J2CIp/nJdCBzC1Y3btamVb9EglTqKmPYDklM5fb
26wVjxf+dunjSs6pQTRWhmKUueG20KAYbLebbVYgXExMHm70cVdFBTjFZIlNV2y+
/fHQCDnBSO/AIzhbNYa04/FGPHclUnaehG9JB1LObskzR1xXmVPofhVthb6T3XSU
cvAZl0RbYMO1cmkudLi/g/QIejwqkK+9Exn0ihSCUoQ=
`protect end_protected