`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 54880 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/9huKRhRMtvnNqb3Z+UU7TahEoHV+T8U3P3ufru7l1O
3DlgtZzb9QxCbOjthp9+wDkjygH0eUfDrEl1ovhZG62GK8cwMf8vCDqePVMhE21L
WUpXIEZIPDJg8xs6AN7FJEjnMEpleX2Ekw+lVJZyazbOFQ0G0eQUhYwfyzPDXKc7
wSOIrx+535PCZV0pPBCJnmpJw+ZJ2jrzDOIhBLCZmORWnAtmhFdj349/goWP2UXY
tXUyTsYKRhqkW05wdzuuGFNLGMHIXMrwVgOQ2QhLZ/ENdedQSW9seUUnG6Ph0Bzy
DaiogzoUplXvNfRCWEjOSHwgr67dgSRhI5zjMHkaHcWqHv/iwUyh7JUibQAfrmR3
+WXCSSoLNudyx6jPaS+PkebUptuYb0sKrjihCdekTGQOQV3e4YqkIIHHRjpX4WjW
cZJjAPC8Nv3y0u9a5wXpTYk+LVEGr9xVxQdUeASmHn51D/T3cbVooKtCJzaB2hQ5
sTg9uosxb5AJqNS+aULC/CBPrD4cyMu6vKjcydAH2jkmPi71xZ8gGBDY8r+L9rpm
UWY98FIn/sQTnislxd+OobOEH9u8HEBw5UMccsdJIW9DbvCP5yaPTou07aEOh/ZJ
uofDF+CnN014zaBDU9Hb1AYPTvhkvFBAxhRJZ0GzasV0nrK7eYFVQ8KmhD/1h3PE
aKg0MCLoreSHMOgAecfREZEhrfk1qq1/b04+Bvgl3C5ot8Is6Xtr4VGdJCGXlEAs
tyqIJ4kMROkZZ+brcf1oicJ0TmuS5y86V9hEbBZWmcLxx5dLDAJpeSfxl5Y6uijV
7GmtBvl5c9GhDGUctPLyvsr/fBrMZJAvk5y/Mdz64lUTTFzYuvbGdZN4R53Fasy6
ueQzCMLBFGKJ0i1sYeCyB7FVAYTIIHL4RQ2ZgZj3EXrSPxxhmEtUgtilIg9DEId8
A+4yGhGxCLTuuwYCtldtM7qt0QxujHDg7kB+xLZ0Sq9J7aARqktoMHCTGWu7Rv8l
8Or6RaXQW4ZlxrwoC1QWqU5koYngMVYVURGV7Lseh2XvOF1p/vASU02EIpAoTame
DN7Gk02C3QDM9AlxHPFzut4IxhPa7p4k6X5KPGAbnHSOU2foczp/Y3gxRxvS254K
s/o02HpZ7GOFPQsh+1gdgt5eHs4MSu+jI8/FyqYdZafk8hzJI+Wy3NQFxlui+rHN
q56xu788hVfxfEApnhnYs3yhFJGo17DshJwNVMTk0vYy/qyhvvL8W4aVjF6GFfyG
LlS61WS0Ykb9QlVHp5lVVVsdImUCLycAiD9OCvMlElz5Y0nLEHGF2jGmFBS6qZYm
TH5PrvBwaLw73+aaf6WJIwdqsV/fVgWGzgLkh6/z7cfd8JtWR9Rr9dBeq4ciCRD6
GY/IA2NG7Vg2SxnrlnucgwTBMuTTX5gEPwR81RIR7ZsqZk16gKgYU/gQjcIcylUX
hOL4ncKGrzALXKnyC6/1u8wFQ7+Gt9BPudtmGZy/vc93ZQUSnZu1M/V6nrHWu/3O
RfAixNWIR84tPpwsdrfa4kSsNcsiXY1kddDuuI3JF1fCFfEbHZFph/Z37pqNkfEW
bgD051+k/8oT79gYiBJ0n7sx6qnJgmERBQAuLQDwI+2LVA3EjaSsWJ0tTNkIGoGF
pBrXMMb27AOPmWN+9jbACG7q6rlQ5kfFbTrAzQR8grYrPcsSVKTxwvw4AiaPn3T7
GLE1I8AjKTweOio9HKuXuVjGrgHZwHMTJzA96IUMykGi8LO6QlZNhJee6x/EmP++
XIlCGZ4ukl524mDguf9OKDp+yXBar8sPX9UzWcFs+Qnr6Jk97dok4nsPwE59QwaI
f03pItO/vAgesu13UyPKEnM+zPr8X3XdF+euI6rFjmo3d0wq3045twFSN2tNnANJ
ORaW4bFKgsbS3YOQrQaksnhdhwrTanFatbqaXm5lUIxpBnym3WUk57YC6fO7ivAQ
T676qspGka5xtBteLG0ujYNQGYY6Wt0iAIFl3Dwpc7JjJlrNLUBuI0bWnlJ/txyT
Fdq5XaCiHb12Jbo6o+sf+FEZHzvKqp7TCr7JwVQVgsCrriyz2dvO0t4w8nV/GO0Q
5lKv6wPgXvgW+OKxgrpPXmaa+SbTdBTF8e1PvzF1RuVdKDlN+9PWQBQ/8EhH5vMA
ON7bE0cD4GfK2pHtE69yAmBGub4XnHvYM+n7rv6VED9SbbwtBD3zs6SceFjoj4U3
GXaP/ZCiE/LjYVqc5NoOGOvokKGE6+UaWjNmFydXBZeIfCcqIcnNNVerG08mNI42
pTg9EhO9z1FEN4mspUHhxIW6M+gI37VFicA/MHLjjx3+yFImHZBo4Uezk2JnsGhs
87BQp5lbSh1jPyMTjYfFTaas1g5AyPGtS4A754OxHkx9nUCBfIDIbIFuSHzmHgFJ
7hhAfHf1iKEVeKdP2BevnN8EVAkd1+GBotrzQKIuQBJOVYm+gq2Fsx0Dt7WMuY1p
om6Nq8o4I7R2Yseb5b39atQRxXdOuqTLG+1i4wjOEyBSSVH7lszmqcVA7bfoPqZi
vuQlkWf12UC1boSJqJmeqYI9QmB2vEJf9/D+Qkh7xNk7/lCOi1Ep3JfJK3Vq/qWx
YAhzqcAxPDAUMuq/tfcPK+4H/ZhPLBWSBojiTULF7dXo0FglWzHWJ3izvFtcu6In
hk1uj/utaji6ZvXkqaPxzAANrbiyfG3XcmulVKpOsWkG5dt/cAz/v/PSscdUcY5i
1lopIYPM6j/vEj1EFIq4aWhvKzj+4rys5aqgYvrL7OJfIsaxWr+XOR8XlHCkhktH
g1lavl9CBFq3ZElbYOl/9HDv5oiHmX5P4uqLTYiC1tDSZ/0u3LNFG+nErTFDg8RI
dx1LDWJG96ibpgen92w2iGjiue9AMaKLGNib48XKop3qwtYFcPAZmOm52T8qF6CY
TfqnTKEfD6PriilmSmI5ZsmoEy0RxE6uZQwHada9BMonIjEDFE5RYpNAA85jM/OX
MOyTbqVb5t904Qc3FZeyj+jwL5A9AEClYdzU0ajoyrvXVk7zOMAF98jakwyorkQs
WlBEvB0q74WuRNLSalPlgL7CTXE6FPL8/tm1tc+MmxnvO+uQ/Y+3xaqLPCfWUdgd
C53DIrS3kkKIsQK80PEXYv0CT5ZYwKApl3/XVGMzEiHF7Xwity8l1PErbMakVzbM
coIED5rGr6tANx4O1/bvR5pQ8iYj8C9oq5wZ3SBdHb9O0XAoeOZEhOMafQ52dYyF
UHF8sosh9yKEzxMTjQQrzz3ajNVcvceaYnPyp6bd9hV0uMvocUmwk9HCvvdOtWm9
mUIHYxRNzyG8dVqmV8Jw8/qIl7s8QKES2ioiURyLzSmnSLzpRDxXvp2yZ+V9mzoY
+2fh+JK2I1IwZ5relqBjgGJIbZ3bmNLEr3DEM+0VhtJC54QlM/uGhz1M7Dd0reh2
PrCdLj/JPRPJ6rK5NFl2pM4rdGj7Tin5ffQjTumROYtd1ldZZAB+6+VDBPFMM6QO
g58CKEntB/nBtQEPNN6OAdQDqFKWxPYcwYSOwkQFImPvlSACTt/8TOj/wasaevSF
peXzCwW0YzEf6U7AV4RIYBsGjDSkv9eu+kw1D+9sJk+QpAWSjbsg5A1jdnLI+ONe
PxK2aSGuRllhrkVN1eKCVumwwUgyGSm9vsOIKv4mp+7tN2OVIaGJSUtBMS5xX0ms
VHrWt4QEp/2WVag8cnt4mLcpyLyrk01lV9nB0QDGWNx6KWg06gX7B0kAM65yR34l
wK6Mch7Gj5LVXFWwPDArPB0BvslpPMKWBFAGVz4w1MIprhIUnc4f3ihfu8fhwUtK
7Zz9t6qzEU8ModydPdYxoola7lEUbm/7rMXZsymm4JiWGUPjlS86zn7fuBc6ussI
zbioMe1KZZIzKQsI8fXeRGFiQ4d81eX+JQTSlxMqOn0DdNxpeg66xEWuXOCVIxlv
o275a/DaG9TVbC3I0LCoMybA8Ng1SruCq0pgCKaYw8s8VrgQTuL/bWnjU8ASdPCi
+e1JaYjoOSlMPtNGI/dMo5i073t0oJCpYmSwEY+HcAXSz8UcZMp7vfDPcA1rDjbg
J1sVWkS1Z1J1nlDpigYF3IPCDVV9m5QrJBqgf9SqvX3C+ut0Hk6F2j5THi6BQhFD
FUGpao8yLISum+vxzDXX4O8CMWTy7E31lyrNWbhDhwePxXpknV8kBlN0I6Afx3P9
lT0B4f4gL4fL7ZiiMRqpBb+luVT8YMPnM+n1EJdePdgb5B7mYpGv4cNfLExANPs9
sYXVpDdpxdnRgoDjd2YLfYHImM5k4AkcWKV+xCznjN/xknWBYSVLmo5SkQMvnKXF
XtyuqN6z79xf35hgcU3M1Z5kcmPRh96lKvQtX+TsHREQkDq4B8szYoIG0aD6nwhz
EHDEn6tZaCiO3gJBQuewBlKMbPiZkWFfKkzQwU9DVCFIiOZHzz/kmdZzUldsmBzP
jyfqbGUMACbrW/L8X2u2hF8LP5T+Fx/T3bQ8Bzq0wbzmQh76CsOjk1n4PsQjtZk+
2mnx7+ZSsI16Olxvy63Jy+mYwq8qkTNgF+ww7gRsQ2CplNGiXe3NA5SwghYZnRZk
hRh2rj2zPJ08zaduLPuzWvrhfTBPwqpEnCu80Azl6dFzivK+XW/Ozq8MojSZb+/A
ukeoR4AHjw6BgacHe13+BeyBdNyaDpljreUD7icbM+fvV0aY8887gOkuHbnvpEVF
pm6b/Rg5i1aLQJiPYEJpeolw3MI687TMpLz4fZHCLnvip9eTlPE/Qqioo0vrU1JO
E4cndSbg6NlxfbNy2yrGPm2ScSeQz+B983AV1Z3OFWwyvz1nDRuKU+iiMKimGmAG
AU7QXe2n1JHk04SIT+oCcllSig7hmaTZUZ22X/tvecbP5rmsmBheAh/jODi7lqov
KKbaq9Xo3XUxApZCZD4TeBFIMmpMDPoNEygdRQL+yYWwaggp3OoWqgNWLo5VG9X7
kYTMrMfMlUDauBEOOLpQhgwIQ6iyNykWiTdq8Hcp+06IjkRSEs5hYxrwtN2Z84jI
J0VTTFFFnUJQGX23HZggGDSj2WdssI902OL1KYu7QmBUIyh7Qop8IfL3oSy9AjmJ
/Aj8uKvie7Y9bxrC1RAXOiEL7lgY0hNQFlQB44Cf9FeBqFuclhnizORFqpSNcklZ
3g0edQNGSyQvfkwWOX18jPXidjuJ1TOBYefIOKH/IDGjL/wTX0kLcVlFf6BYmGaB
c1QU1mD/ne7Q7krAlvxKKbr5lfLBant94TNZIIK5LTmRFq+WoKkXHs2OH9zxM+Rf
/5J2idA3WjW/mLOv8osVqfOVVPMADo3wH3QZODB57j1a8wzxrysreo7zOqfhGwhM
xJqDqHAsf5VLTNaj0gEoTQ62Dr4vAbVxK7MhIJBjUJOwIKEYOZI7RhRpfUrNE84s
OWb5jP5E6LgTFJYe6O8DuAr7vp4Ay/TZjE7CErxn+gJ8hc92qZgAtUmV2roCFQ16
wfAkDYJE03Byyd/SFlQ1CXbe2m2vN5zd37/SGd5nzx+bnrus1mZRZM2o41zrv3On
asmidAsq/ES1mN7kai3pw7DEX6bRvPA7PBBnCQ5iwn4/vfgcvDkel+NfBjzomNPv
CiN8OW3GADlSz8EN/U27UbJsbCJwjeSoeWlEIx+/Hc3QYoafZmE9WDvTBcemYjpQ
MrgmcvV3u0yp27iwsXsLed8Z3FEGcUV9PuCVgL36L3WPxyZMufeE/0VO47NqJarI
qnhpVGj/NlANKF954bWL8LFMtsVB0mySCr/q1whcBYXqVfYZoa5LZs+fOClVoVkj
M7Sd9yKGC7gOhM+9sVAZR3jFcrXap8bBGRcbIvF5WI1H68yF3MbzbNtH+/hd+xwA
3HCQXZfnu2/W1qdywW0DNbSvt3BIsD7xExHS8HgfnA14Sk217FObgaOcNSB8yQeg
XBJ1fTpyfWbwDvAOL/L0hE5HdUPUVlXKays82V6M29D+Xjl1jWzP9z6AWiDc8cpA
qY68Z5HRprlQKev/igR22X/EO4kAX2VhyHC6RYCu2/xxQNv8wRW3pg1FWRSk24xq
IFKYAFRcZoOeRs3xTzICh5GOMrgZhL1YlTgGGNajLu9stBKM74nCITBe+0im3q27
CMmq2oFoyV7ko4YJXUf00GZQ0f9M4G1sPH5WRI73Fz9IQrdc/vu3DRDhgSaWvALx
/gfPZKaaP48XqNLQyT3HXL5z+l3axQSTCpNM2lWSrCp+Os93VG7cI1BiRksl2rN8
ubduKEzfC23qaC0U5f2SHDR73PbK+TjYyLscwrkCLC3LickPfBOvqfNm8/eIdvtD
85MWzaeaonCtqtNu+MQesKSZJ294ZeJzMbeCZ+gutCGuVaKH+/XubBZB0jyG3HpK
SC6Jzeut2LRFJ/YK+/yyKfBp+SEtLAPZodRRqr8cfbCS2lqq/uWMzZfVJhyFIMuF
dMmLE0Inl5FWm4kNS2nYH/hQqGvNLGmk/Z6a94LEzh32Yn69wsf+0Fykbwg+w5PM
mZTd+aU8UItnLO7mnwIFzhhrgA8/do+OYfFE4Fav3PMUWg7m9Wy+VTslC6VmyYjW
aYSR888JI3WLRmlH3lUnLM3AJs9hKlVZcqQUiKUQRkUzLxu7Ydr3hiJvMfq/xPu5
R07v/wfp5bmYumVn1rH3Lpi5dOKps5ZoT2ukbGDrtS56EknREILdxDbJEL7usMs2
6iIXaIFBo1Mf9XYkO7LgJ8SRrL4X2TT3Yqfvx0T8Y6/ChkmwGCz9zQaXKOYCawTd
wM646iH5I3dBXUB/hokvSw65sBclz+gSZmGM1lq34HfeyGpgzbO73iti40jwfJna
e8GzYAiu994biT+qYxiPfqK7d4vBGofhEYV5CQ0kjToMxRjLSTjhEsyGqEpVwhEP
mCeP7/L5zzIjhkWCJZ++qIwDJoL5Wa6dESMfsoRZKB/Un3b5gUCQzbZayH6L8I7I
h/X7Qnu12Hv3bTFH6ruqtpTc4qgm4lqCwV6p5RNMxxiMyayOVZzj0181vFYKCBqM
Yks4REdbB8UOcfntI8+vohbv/ou17GsoJg3vhxO+f823K+0Te2Rx3nVZpnpbxK5y
4JvqT323TGqOg5im/mLFabVXNJxQLYt+Pxo9G7bWTKjvaB9JuJ8GMrjjp398a+g3
H2FwFLH5ARa8iXj/9ATA5Kl2P0Pw5Kwkw1g/BFfsbC9xyWgzdUxeDEfySN9JCaMz
cQ/Hxy5qN/YqFkdpRiXBB6rH3xh4qeoN/LrIBhiyuX29EqaGnfPZfxuV1OycVbAu
SD+R0ciu4hKUPN/czsSjTItNf472koF/Dche3S/wfr9oM1yrUyv6WXPxeyKlbNfj
pGdrdyHlKp50RncaJQbp26ZyCYlTlLZwklpQ/yE7VlNAfc8JpuuOLXDlDHqJCX8K
+ZF6NMgwyiECxDgqGmIlBNvInWzTNX9RHko6+Jwb65qSWm3WcFSSDvd8JqFnCdYe
far2/rFQojb6L1LJC1xNgVgGD2mNDX6qihKuaZwyKwQk2xIE7SoXJuPsxYQg50BG
geSnS6v+qderH2bQwWyM/2xudIVKd2J/9t7L+zgd3RujIdAv1+iJmlvoLX/EPm68
rP8iryAX8+Wz7JnArEPd9EuDyiVKFZ8IiEQ33WLsFYpvTb0SAaye5NnhXsn85saa
grGL3UHdT3DOudyX0S0UIbaHPBqjZGjYx8MrvyrIsjevl3hfVfP6KO+Xz16PeVpz
Yr8jKP3cP2K72SNqs3j0aYHrA10QbV2L27zpFjf7Rp2TM1B7HlfyBYECWbZZZPC+
/2K3Ujl2biuT/r1ePQ6iMfFMpf6HLqXf8PHznX9hmKIDonJSqjruqfKbBLmMHMKk
KyXmFXiw/BW7bSpc+UEeVV5AniTnw4iMKDj8zbiUC3CqJyAckkjlYG7wt/NRcGxL
WkOkxJXyAdy6JaTCADcnke8QwNWxIJ6L956cmt8f2/YZ8botJTEGPU+6aMqxVydx
c3k3+iJJaClH1Qn4INxU2xuql4crUbcKJk1iQWrZT5sBJanCtP24P9JQhTzEwFJB
5LYT9+IoYgpZYmtF7UYnlf+at3+dB29StnC9gWBJN4bRw372Xx+hO8MyeiY+2sit
Y8mntgQdxLJvEeNBrJvH1IlueMLzbVNyyQMHxJI8l6nswFrDh7W6BU9wYmx5Ybt2
TBHzLzH2WQf7x0x8gQmPWeSRjamvMotWRt8hMih3eKCsWfKo/J2U8MhOkNkHHM77
P2EYAWJDcQbOqZPhQm3WNljTyd10QYRTTDlL+DxazFDlMTETI5fKgaDsrCluFba7
/ZEdDxUHAgRz060GB9zGWfxeasszGICdZC9DybI6YXtsy76TqWjsm93NyRx7//Ne
JcF+SEY1aMMO34lGCyYJkSAOJ0lHNFLNkwt90ftEi4lObMw57MG7TYjY9ovkp0Cl
Q5ZqkaNA/ujcabk3Rvi8nu/gf2JNqv5RID67CbiGZ2t7WgGEFxeOlJCr4fQ235Yk
Y/e601dkMxhhyYxaaWf/+kHlftgqgCKp8QpdnypnG4+HKH6Nxq2KRfw3Ky7Gl851
Dyn8mWMpJHPUnWn5Ig9lPWihUDA7+ggwlfgEF+C9anvuOrfq65kE+bvd0iECklvX
Q3Uu3fWQsr62lT+qMmc2DM5RQ3SU/B5uJzUqcz60FG//TuUdQH6ATHJjc3gmdpnJ
3Tmeo9vfOmSQ+Ob1OHuevToor7p8Mz4wn8i8fzw+JlnjW56ptAZYf3htopJINIQx
t85fIntgMdy1/N2toE4PCQgnZRul2ygbNyhMBVgdZmJkR9Ny3dEt/lav76/CLlhX
F8N7QmMtc6b8VjP92eib/pnWUvtDa1WnLXifNNb69dvF7MrUw+e2Q7zh19dk8tVF
FhhRCwAseoAluXKnod05SAqfFtfpdznMb5xbeJpHPG3l3JbP5Mr6LFvQRwMRj663
eX1rrj353q1FXYsOiaavDh2Kz61hVu87aSoNUPIbWvMaOCLV+Qszyj50Er6tsKdL
bbw9llkg98MfdCSNuOa9uZ9YaecsoXxeIimIjByO7/rzBCXXHgimFxCY1caUbDY1
eVWkyHoT39Fn8/dsEr9ak8wXrRw2rWQYIfAC1qnPDg0p+N1ZG1gY/Seyo+Llk6V0
mvBLpuolEai6gc1D8lgOQcK7/lR5sLcvt0gBQD6WG80o1TsE2I3D3ZCuPWwsa1Nw
VW6P92nog+1yMHVhDG89wSFvkiN0KhSPtb/spd49vF2DDQ7Tlg0tmUr4prprtKHA
ReedpcBNexDsKmHdFsHq3zhU9g7FhYPFLYd8Hl/1trFy5Ojyj4oME1pi07YHSh2F
Oc740RStaI6bHGA//Z1/YqHCWueYWeDYRVMWlYPTbG0aj3W47uqHjMrwm/KSo7Bd
lpA/X/frwaCjZsCjwzIK2ffKL0NjnMQjnokX788wwHxDZCunbPOO6jcgPsiqnCdL
s52SjKxUfaW1Ie2Xwr9jZPqwDiFJY9MLiKDWmoYpAQkDQZjcH+59QL6+vADpw5w3
eN0kxs4C1nL93yltybJTrGpmQfYtmnloxqVjWz/xB56qAsBtusqza3OvLQcj4bvC
lQgb1aGLRltrXFRj13TBod83CjUHT695Lhp0SWOKAitQQF5uLIm54Mcaj1MUWB1S
gC2+ChPimnvGw0FY1Irj52MieseRM6O+/9+d+aarxGedyViHj6ukbOp5pZ+oVoA2
89KGjlT5i/jVwNfq9DOhymLWcI5GqZK9Rrdl/07SdImSFWUyv6rHWDjFRvtN0KT1
1c+/oC6aGfjeXHu8ukbtSkAGAC9NpHn8AWpyTj8pTwvyBzKDYtlwVcNqAj7XP72u
xJcCgczrVE6HCFCeNlxfXRabfDW+48p+NZjz2vm+oW4e2HSgrl3ao3d8ZCWcAwLz
WF4iLiBiWAy3nXReDMZo9cLpkt6r/bOLUU32NBs7tDQB0jsd9C4bRFRNlD/CFYxH
94oAmHf0aX7/dBWmXcYCxjkV1sLQp/81c/ih529cZbXJoOTmPMeeKc91Xerb3fe0
sX0PcO7ITcNIOTQf1qHqFy5PpboOvnLiwIZF5Sg0iTRPOG+VTW83aR27TcIFWhPG
L4K41jEDtThBdha4xIi05k9mCxq5/KFYg1xGoxDz+Ph9OBrWUXvazwCOn1ll7OWa
kQkreojYT83WijqvL+luCkq+Zbtr1TVRmHLWSl5SaYg+gr31//GCQLlAeUaheI2L
+q/EOUJSwsHt6A3+h0MrzEhUCRkNQysvrBB5U/gODl6+6cZwrrS5dmp0P0LsPzb5
ph1d+Klr5U8/ufJjezC3H9KH2JGimqeeFi/ux5XKuL98n459o3n/F5624b2E+s8x
ndoYL9On3AADuqJ+I48zjldddXTP7MpwQjSp+7vJPB9ktMRqYuSuY1jhwU4NxasZ
wCfPnd6YU5KJfsPeOT62UYoZXKPxvWKwgDr4AGjd4NeXvr2iIXzfdavLZCdOt8Uk
RtY3jAt36KHovENNZKOwAGTRVq4vygGzDW5v9Qd5an4Ti/WFro2SdwofXi+S3QwW
fdpkixSzSGIVplOyl8AY29i/urKKosWWRLApEaGC6cq3h/wsdTkfXP1LBdmqKXrE
7oW5yXgRcYfyzgXfFMR4foxrfY3oQ7s/7mpp2W+DQ+ujONH2RxP2VX1ZlCxJIraU
rCoEpPhKCAjR8t8rYAxw8i3OZFXyWqkfsSMjLY/WiAl7wpgaLuY3Ry0bcbBtDnyS
DfLVTuLMS8ABxD5qPuk69k6UwWoR9/TAdxEf5P5df31VYJIgEDZwdqmkEfhkQImw
WL/jTzKTCB+bFemqH+29Nz9/V7UP4iC9Fej98Aq0iXkMzarZy6tEQMQNa7Sx70S7
08brAY/6NnmdAIziVLgS5aXabzPWJCISHzUewpKfarMyYRp+RohEOGWrEAfzOjuW
YnFYkHn0vHCgxW2PsnrzYa6GyIm5LQg7gTx0hcB/KfNqKQvVJlOwdRYtWYv5sitw
kjsrKBV7su1+D8GqfSfoXTHSc5MjB+aiSS3ieHKHcwMFuuMwIF1vmKHk+nKXTlLE
neQ6/zxUpfc/4m8TaJBlmuYDVcZdoZYV18jSnGX8/u4UBGWJIDOvDbQVythIXUew
BtYyjctdCYONzkLgV1/2whIqElQfsIZvKqGXN2PoFkNnxjcI9fd2Wty8QWRxWIBA
AYN4tpPK8+2m2D96LHaOM0EN/lYFP0q9+AKCJc8Zna8WWkATdBvZVxCl1Fc8LB+O
tVdVJEF+22/6wKBzsOsnN6oUTEv9nPCvb9befVYSWmm5phZxISTIh0z0uWgUgcN2
CPEc2+rGn56Iq4UxYWlkgMXurTCacuPBkf5dmmBIDeHawwpL6RrixRyWJAhLsAn3
Hrh002yslWKDvKD0nmL20gUy/BcDPT7c1C3GwCJS5EnbUYZwr/q4/9KtG+M4q2a4
akwx95UZp4xNzkqR/U9Xikel/4f2ZKxFFxmTTTEZf2oVDo10huEjRP0BTpfQcuR2
TUDvrUYHtAqyYs9fN0f9w9YHzuCM1A50l/6LYnG7p98HlLqPH2xxVXm5I3aI2NyU
kHK6lvV1uIex94IpGxQB0iMDAlCC65xsdFwLOhxgdPplxfPM4khi0EJSZupJiOcc
zSTKw+JwMnzbD6w8hSO05v26C5z5PTrkI89Gssr9Za+aCQi5Gm7cvy+1GXgfRyHY
I3xKDMP0vAynVpKOuKXpuBWEYRJwRcP0HwxzPlEZVHN/BOy8DUN9sueFaNvtfeyv
SQjHLOg+pDz1yACApMEuqp3dukAL+1obAYRhUw2JXEDaapvkhVK++Qy8A6D0z4dN
a2RfDr/qKiqY9oH1Mr5JA80JL1DBKhiuC3WhFv8b4TMVGronEd/PG1Z7O5uGkG6j
X4t73N18iNnRbZ3E4Vc6oabFpNNREOZH7wKI/LzyhBUA+Ai/sHHvkWyOfmfBoM3A
Lx3yb70gGS/QMhqYpUa/klk6QiIUbwJGHTqnsUu7ybc8zDdSIWd2iuApvmBah8pz
lupLVscKnvGrr94aiXPsGpOYy5i9PS7F9a4tjMXkqXmyxQeazQJ+YwAsIxoBIjjG
mC3wLmqU+5WbrnN1KnWwdnrUtP/mQ3nViHrw7jFtVqsYx0ABCm81k2IQyuBe27dK
G65YNRFgks8kDdyyiwpThuhWrIhbujYGs+9WumxEKc19L4+/dyvdZe/W38BMOzX6
px6/UplmxIMHnbedpTvpSQLGWi65zpSvcDEwohEUkkZNZzrNuli4xyzCx0UwJofo
k8kYqlH5qYJTcLVpEPL9L/aU0qYogN9oSV5l/WnfPqA9rR0JkT9d/+jJFLofc7l3
Fo5YU9JRnKHCcOp6I9MWs55syGb2hlBCK8vW7W5oq7lJl8dhad6yx05UI/sKqI25
/uso584S13wO0jjRvc/cxIwQ0bDYvyq7V9cZszt+qdH7KnJSQqhtMezDEVNU1EV0
oz3tm3vW6FAr/CbUYiUTOmvvfLyIjBGi5tT1NWnPkM8WD/vJ+YrSr60geVDZVALn
NXxr8ZvdOioXnCwrPic5bRvyLNfkW/4RDD/xkezasOO/xtIjxwnyXnSJoS6LLclB
kZ/NQIoD/q5rrlTjala8RMwvVWNEmMdIvIa1GmEvFJ/ePfraOOxv52VZDafaOUz2
u+leRXc8gYvwm+htLSRSUn5e7CHRqmPk90mK/xnRzubeCoyzK4teRYE085g2kpdw
UO/gwtXeUFVx218MdTWOODhb/Bb5UvXmsS8ctMNYvoAd7uh4o+qnKNDadJRWKdFy
IFBsbZG3QPkWXIAUoSKexUMT0uX4lWSpmqTAtgHKnJp3LPFzL0U5xGnvgHUvIcmN
FqxJoL97WUJlHo8B0cvnKcZm6pLiYKL2uYPC0BYvVt6cvydRdTYBnaP40Iep51CZ
bNntEyYDi8VXCH+aek8fOCbOXCNGqPLtHW0O2Tp6T2qNLs0YBOKxEO2N/rCVuLt2
npQOHM6pviMY7ZPcBD3DGKMJK/CoM2AOsNsUCDA1heMDC5bVwfEgBAdyvV2tDK9N
lkjauhn45b9oIKUIEDr0VqlHuPxX3H7OoIFZuIrDufcyi5XwcaE00a2g142EX31e
WvoDLI0QAQmyuKsgaR/oHC09AQJUP8hB105fOVOWai/pFMn3X3UNfaCtGZdi7WLf
Wh9eZLO8iNuBW7p9HPGK50i3RF/MpOeuUT9hEgALQnC3QU41ggKouNujo2jF9Aow
+QJqHIDXZOy/JAlqN6e99B9qVTpBvNimfFIV7cz6ucOZPuqigi8oVAUO3534rExa
yJv5N2Qj02y+Mq/8ef+Wkv6XsuipXKqbkuMbn7ZksAGBDhblhpOVISM/RbBA71wb
DYHGULNe5aNz5UJKJsdux1rL6b1JMMzlkcdqknhm8y4O1aKzaNpPFQPFTqFEbsEf
EC/y3oRahVwroTaA+JDQrdGHov/piKJebSbg/vbLgpYiL1VXJoA5P32SPBE/lhic
bho32BMbhUO/EJ0NQzK0LMpAL+MEYCWs8Sub+HytRYzjh626mhxp2QfSfLAXCW40
GhcKKfRvY1cyXUYArNw5l7wkxXjsWsO8kqdUqXCZl6CYbnB1tvtFo4UbTPOjEcF9
NKS4YlzsoOpx25hXIIXALrBcNf+tbNQL+w/TispwMQVeyD7DbpFsaFuyGb0YPFw2
o3mYO9GdwLMcg0bWLy0qtpWEWxUSsgE3evqt6dVeO8CYl2E3MsCbjpvfm8ybOmjK
+OveZVIN0K6nr09yBLPjKujJ6R69eCBKZMQyjScT1amCtuL5HQBuarHoMMeky04S
ifpLTSXJaYIOlzr7iAINXKrlOKm/1CHCVotkRenPGCDD/6eZ1KCdmo87M6u5Z9wK
ak+zPxazZMMHiQ9LsvdaXA5gTN9E+W7gFxCZ4Tp0FKsZR+hlJ9jtbxwYOkkRJY+S
4tKDyb3s/f4uFyncsmD7TlniIxc4nAeofZcIjuNeefSSS9J6ZguYSGIOwfPmsNLm
h2EfDtjUbdvfGCBepGiDJ0GRStK3G1B7M5hpPuT8nfFswnSY1sfsEtmoxAwPn2z3
SK4N1id+pTgpKxfS3t0wJTv6D87GfW7xmrXTw5BVvGaYhPDrj1DKJDxrd2Wvn4mC
Z65c3xNZeerZ1rYylss0WhXWRMNXs8wmLPIIg57zB3lRYroElXaDgBaEPbfxqYLh
l9pzXa9f9nDwhW2hFs7FIisjtEUxke52SdY6ckgUsqn9p4+DtMC64IPIR8DOi3S0
UP7cTPrBVQwqGrOvRR8TDn0mwDxUuKFQn4HOcIu2B4BOu5AOcrJ2JkXvWbUdnHqU
7BnS9Fx1HXt7eF3vUQQdLvP85UzCw8nNy0xK5OgVqp2PVIvEk4XW+ekYWCIJXzIX
HBvpGDuz1nIoVa1Fns1nkHiQdQBgF/D1bFYPLupfmfeGxWHvdDYazkARoN9wi2G+
uT2I1CtkH2jQaravjAXDdjWvyd53zZ9DtCJy1djbPCtVU76UPx5H2bf75NrbupyX
xSKT7bXd8FVPXBk4JUfjyPkraZbNlJYPdT9WUomzhjlTsPN2107zi1drfbocCFy0
09HiNhDoEGUMUG2Nye2bN+EopOfvtwHnzlZyQfNLPfBSDx23PG/ea2x4ip5/Qh/7
zdFCpUh7HJ5DCp9EdQ5E8yRJ0v8F1BDiDqR1G1Q5uRphFRjIsFIfUAliKZIa5iAu
8ftTkuZ5F7EVizgIbtVurR+CGQDD/FZlGT2F2ZqV7Jy4VgDeeWj7yBDri1Pfo8YU
rHrm1bRnF5oGVWoE6y8f83x63MH8UAoyELFQ5Tl9pPRuUTBnkS1pI70egJo6js8p
4O1vW4m1TpU2aVbpFJocHhC5SPGgYXeIM2BAKGWvOoEtDhlWKsDFacUBvOf6904F
/pQTu9G4huTx9704bB1q5TpARoZcKEP/2YufSdp1EYPf8RKoYgTHa9Zne2A/39dq
WrI99UxWS9vrPb+Yy4DMhB4Qitci3jX5pKFK98uWAavDigYVbtG/Jp0mM8ux6Nn8
okmRdLYVHvau/6ndcImLpb6Gz9vI/RsivzzRlkNqj0XGmVTi/w18nG/tbNYQAcg5
K3o+EAjWdvvYfjIl56ITuBBNR4+zvXSs2JLCzRxw7pUfk0kXv9SqNZHPADNIdyzA
RCP8t/ZSTyrhA7w73VCotUU3rbXh1ZdfyavONwI6ufVaXz0T/sMk7D32L5EF+W97
GEbAO6NpTGTbm1yvKX/NnxWupquFWW8HsCjVWzKmTqRahaqnioQ76Cj1VeRdxofg
cyi+xiGfF1PqHzNjkMEaxVt4eat4JJZjFc8oYoxOWrVON3KMOM1+42YiJiUry2KF
MD5wOFcbfrgFSbfWPBxrzpurzvv7X+elQMgFDuJb3chpDzqPR+QwRGa28pUlJLmY
ihPPDBJG2ZzLFdsqt0rKTeJxQdp8XC/m8zLt1DZB9CJpwhV+pUE0lYaCzW31Y8Bi
Ziz8efvTyT46nncFcgFu8tz/kH3PczRfJuJCU00oeYtJ4FWC/81tJSuKdJ+CyG22
K/id2UXPeAh70SB/lkCQZFEuq5fAN5QFd+AicwTyOsTqX0r48hquWRaMNDDAfWLF
ntVOYFL2EUh23zLmyc7rMYaTpAXOo9if9kqMmvhyuZYeMcmZhoKWD4ffXjwjtzcp
WjLEKCNV42uyvGobNkzE8U1NuKaUNZxytHlhbZMOH1Hy38MXIBr3jgvd779Pfp0B
uBftnF7kGTulP2L/0wzfrb2Z5fVDVv2+TtjUG5CA393cUMtsy6eLQGQbRUXmMrrD
V07KvmKvP7HSrOpT13dWx7Cxzcc+nwo1ubKMqRnRQT4pxuBtrU8b78kg/yjQ4E6s
ipBNeK3neC1OBNfVC3R5bhYizbUOWgjK9Y6Szf9kGswagp70n/hjCLg2grtz3XDL
BvOJgaGQa0/Y8LVCcydggxFYVfxXwj6piDgGhDY1B9IoNeLXx9QPbzdygq8kA49X
G9IsL/Q6kK177BIpvSBFUVji78tcFQK0nHNVKND6+dlPcF2YmQ7oNVcEEebZK26d
Z12GhhrgvWCHVNuIMKnw0GFzr6SGeYnTVYQBiijOBgSN8JDcRsnCXKK9LTVMnuC/
euY+eQPhbTJq92Wfv54qdtHZzqqhDQ9DWHWQ5hJSnwJKYlrXcdhqm7a1bX8nEI4b
X4yzklYNKFPcKqvFkWeYDPoabLDw1blVzM3QTxUtHpUN0qVxlHZbrbVDM7g0N/ow
OqXJCJCRTxFdcZDDywyBH3p8Kx6X/PgV4M2DmdQmdtBsP1PfcbA3w5lXkGTiMQBQ
/lfRHV596Ys5tFvv4LenEPb9WvvbFA4FtCyNKItGkd0v+E9hC0REhhSYZ50cgEoz
5CcWgyf7leSRoFm8ezQMni/hb3pUAuL6we4rCtCB9Oj3XNtw4slg7ikYfSmHhCJr
Eqy2U1/RWANiLOdtgyWP4/z0vKGgCuh5sFihRUnRdxL1660jXQbHbcNMvFbJLaOX
YMe/6m7MDsZmzKa0C2n46AFMFaWgIulgEVxUFrWGBH23yghaGeC3FgN8QDtJU/J6
m38hxcO1cWTALGtzUBCD3P7ghH8Ybe/UcrbAJL1gWqZlXKFdCXM7g1trlIc0CNcx
nfnzv12DU3kQLl70tAz5sS3MDjYyTJgqPSvmOt1f2wFB3g8KLc5mC2WVYJ7PL15I
D7qr9QlICaR5adDdfTGyFH2ZfuDSOC4qoHcPifjBdEK+hopApzCYhW4+Nsc36/ht
hU/CGyjoaXq6WNL0YcIbUC5gO4O/876drQJxl6EK7pdwVAjpuHsDXS9659wkH6Bc
lUsVfrrGVqwBu53AX5yK/MHPp/1zmtEadoymGK6IB0V6Q0kFilcOg0FGx8sHXsnZ
RQQai0Zd6QCCPyD2ZlALbFoqZKdM6GN3J8yu8sBuQ03e4NLsB3WlV7agijw5BK+b
3QS5NgXBVjyEu6RVf86XvjL6dlsaAj3ldAujRk/kzNZTLbLSdtV8fD1sN0CXna0t
cvJUMXhfRV8nBNQlk7YO51IUKBRAFwr3DaIXUbgU2/NZzLpRUInz22Vp9XOH0CTj
nUC5qbmuI0Diwqc4ykghZ+/Ic/egcW2YEy0QgSr5nC9bOKrnnCG9An09N/8UVEmk
/1DudcnI4FBXJiT7K5fVVb6VjRfcpJRwiLsEko/Itj9sQHsGD08lw2Dd5+JEXqPQ
8yX40vzaQFp5KurdMbnVGKNVOw+g60CG1L5sgssSjEn45o/Liw9lT1MnkcAZzq6Z
KQk0L44BSE4XOzz2LRMoPJ1/zTXgA/CDwX9Eon2rq96+5UGfqW4/bIGqSxygaMDq
+cMLFsMgusdn63xFW1cDcGu3cs+CoDcKSK0HgE5kQ/DgPayogVAivQ+ABI0zdR7o
aypRTNyVuilzLdS4O5ByW7uhIOUGMu3djODyGr5Nx5C3lf2aQgCPcFJ4Dr+0YwsR
jsRx4BOu0SRLYyrUsDyT6/r2um6Q8+wK/Lc3FgA7jTrZcTZIEvvueZ8UJ/pFIJU3
SGhBoLKSp0RwLYwI+YV0i1kW5HJHwvmVFLTBgdeccc1Ht44iO7Za3la/SuUDppfB
ajUxU96TQJOuTw0sMnC/k1WKFqFE/UZYZfSSbZJOECUtu5whBZwdZNaRCKiUv4JU
MyENfLLlHX1eDvSy3uEt7PWrWJoTR7T6mYnWjSrG2g+hx2znV1qLkArGfuwRhUC1
CDwXqCrxI0ZAJvm4eEHL0nZqi7t4jXB+uVeSIv+lDXD/AtLVAbDUaE66SL36u7+K
qz71oGiuEgC2w9ZKZXfqeRIxKhwKFxXW2fuUbcyZdsmbzwO7/e+f3AkUTESRgSNx
oJt5IH3foWgU/9CagZvmloUDn5+oBFu0N6cKujqVlje/r9EXltnCZOdxtxwUYA6E
O0Aq4LDC1zCrAvfumqKInQQWeCEN24os6wooePS+MBly6U3atELgYBLoW93pNesj
LZsY0wDL/B9fJg5vGnXD0aKgbQHLkSunQ6hIKfQ4HJrnazuy3dVEHMyXqMT71BNq
6r/+LoUNOclvhzM1Jzu1/OW0c07Q2EcUdibyV55XmO6vt5Q3QgjPmspqRUs6XvxF
cTbZLkuv8IqgCZahq+mhRvwcQon4edl3jaEeWSomHVMwt+SwfBjJ/zuAhHC9GMzq
ITxtNY5w+wmdCjVVxavkUc547+vJA2QMCGbL9EmyfSLABSH+y9M+flxkCboD1y5/
XRZkEigV7Ao7WEYeZCM/iuhflEoD/oE6bflk0nm92TVd3kzCPrC7pBCsFuLYKv2B
DX9OFJojjV6jw8h9E5GfoEl/Ptbl5rhz+WE7ezCiE2AVMdrYY6cNt6FYFVkYCfv/
8AzqJ7FiXDEEn+16KbbINGfRs0BiExbBkUW0iekRM9aFIfDoLHjKCTW+O4rEV26N
FCrkOHicFPK36bsJUf6QJY/gh1MNp6C51foDLWCPaCtIOxqBgcOHpRpfXB/B/wHK
icDGc+EknZzRkeNqh1YopX3a4zev1jwcIZShyx7TY00+AefPzPAsghVNgGKa/1lh
7aJb8svsHU1+/HroQtrVfg7GAZxfonnVwdp3T0pPSEeSryOvT+OHseFRJvi6Z47Y
BEFhr2hz4JDluhK101EfgXs4X+Iq84KcIY8XMIP9L/+ffb1NiK1Q8QilhISfzVok
HowUstewhHgVCFTk6+uaY5JWDBdbfm/tzujOD0GUd9ZSRv6Zbm6TJK4hri+x81bz
c0VArpZRVs2Lm29YQNAYpdHFJdj/9pwRxUPvLwoYPUebfOvJtoae4ko+3jNvv5ya
ENMV22c+Vcs+cQDMk6UXhoYtka6wSY15JIP4FBMvtU+iEjG8eMRuCSBrClUaX46G
GjtONeWwA1svdOHJbHpAa8LlkwGuYlfRHbkFBC+4PKW/4f5EqNKs78ACh8OAAuyI
rPh1yt2IH9nwReR+yWti/AVrKomQXBCPf93Gi1oaNvgQNtNB4UNg1zrIh6IjQvzX
+vTDIvySLm8i9eK13XEHtmujzkZ88rKlh5k8w2sS5fKJzlrJNCE3Fuyz0TZXXOzM
Y1rp8rTLL5eCYOfHu/1ewlN+d4dBHmtBX1u5bS1iBHooLLavNuJguT2fn1ciLJ/h
CLJRa/JirSSe9j/j1QPytI60DLQJZ68f+fSjgDJGecKjrbMi+Ugf4WFJn2FzMol5
uGBa6v9qPsno4oNB38bCRq+rJMhwfb7ecQtBJ5426UvI8r+w2yGTwaIW7k6BUiUX
LPp0g3dmYfhBZQY5Fkqrg9qHSgK2C1iR3Je8F7Ira8CJlXO7rVFJuMbRI1r7GFyj
1So2aB/6436TgiHp7I9282OJZK4a/yBmQnmlcGR0PKWXNdUniS19HmB2gAOdzB70
kGd3bzFUeAz95t24bSlgndaewAdVk10zI2eq8GBpgM/Qugh02NN8NLqoyyQvlDVV
AMKAJ9qFIyF9SOaGqLU4zxmjU+f8IuCAaKRex4+k1es8gCqYDhLMkNs4UNHC6AP+
uJE5M++3uJ/STwbm7BHfOvFT4cuB3GZJoucl56bUXelgdbbKLHyaLD0f8qPdUTdB
M5SDJaO8LbJ7JAJls6jZn2aqgKM6av9LDd3hEP+fUK2kSWx4wOSVtwaOudYc0Pb0
kl0Y91RQsDe0lQdUDtm0392mETDaw4f7GWCWy5DGWCtIvurP166s/BN0WJHsdwXT
5592oo49LiGqcLgLz89xb8pjMwnoHi+VXMsVXIgYYjX/n0wznw40lroPy46rP61U
qVulwPjpmvA5pstb6HUs9PnzqEcoGMaXDyG/6wGpvFq0ObhGLLmMwl1nAhw0w3+Y
fjH3igQqtxWXV6LX8SNSPtJChqLpTz7BBzMmG2ZxmhiDVYUJTFYa1pdl2to0fWRL
FreduxX7SgFPry1x1xaUlOVJnEEDvgDeBRExqJrKFPECuljIGB2xUHz6B3LZj6o+
RpZ7N9w0xlmtr0WPbIi30soPS0dss1mRB+9OiiqIulcjE8nxLoh/qFi0kfWDWrBO
KujxqZdt/hvghzmuwFzUp0B9RpvluJblhpIo2ddrO4iP7rggMK/CsH6BtZQ3RBMA
EBhWsIOePsgMADoW+9xriKg8Dfb5egGDAbKnoUWzkp6fJpVwLHjWzX34xxIoGjoy
kxt9JBNM5k2TFlpiBb14E+RwvEdb5SlMSvTgjjbbbyZd8PkIfrWWF3lV+4FdzKQP
D5pdg4u4atXLMQeNiKavU70beP/A2/7EhRITu0iAXbM5x40nSSgzjAYhR4jBMvDZ
9xCBvO0yvDtkafiyoLtWsDLJLamDfCv1aNSE72DLJqbfW/zcbei6wyBeYlaPLTwZ
64/geD/ZBb9RTSZPTMnaUBYDS8v7r4o8PxScFoOSriBtmShNyJbNINjvDQE2qbAk
b5/4RUlDFzzLzHEf/clBpMF3Za5LWW9yIGdkzFkSSrqUALhqB6mi6u9xslvcEsOn
xKAgU/yf/NjrvIEN9E6MMdRZyqR21a52b2YE/PpRz0tHl8ngrh+ay0bgsXaScBRt
ehddeQwIJljftbMoGPqfxoSR3Vf6a5ZOQPa0xoERJJ4qQ7zkVLEKWDRu6HGitaGN
p0sUvc27BF5MuNvNNJb2ffFngl2ii62KbNWZyrrf4CTVvYQWt2gGA1y1Thk8awJD
u7tIQ0RIvVct42ol9s2EPL7GUW6iDjAtUFdKL7Uvz4+n1FWKWSXr1Aj6V9A/Yd0n
SzXDi0zMueC/cQxiiah6l4qFQKBSedLiiUnfCJrwI9r4WkDPqy9XT6C/G/QCJWZW
QwjEdmhTlJqiH392vddZDuyt6L/27yRwNVJbQhQrRgj9bxIgdcUsxMfObO0SfuhF
nE0ISp52yXYys00j48XX+UCYvd88K2Rcn3wHDLzsbQgvKNpeVR3Dyz1oKYilkVRd
AkSNPKRClALYay6T7RNNfK23pL7agnjJm4pV65CFLROJZMsWvutbhyqqvAtZjjTy
7tQ89r6tw59tIbF+CzNKUcx1qWyl7Ff/gP7EoqwP4meG3ws3xGyaGvt4fxOV3mQB
Eq6Bohu5vptGNRnJSrsnvVj4WTUcx3hkvDHyfzVTXb/0+qwdymwkcImAN5l5ff3v
sq5Fy5SbVkpHTM9jsz/GhQH1PMYr3SajYhiUd6LvpC2E/S6CTf4vEwpi0eaZZyuB
l3BXxfuNbT6rV2PeIRNVDqXoe4fxSzW4jTMZ6PgH5yWxVV37q3eWgMoP45MX15SR
kwJjQzb2MbO6IbGWLZL1VxOg0yRAatfDyg/ksALRTIwVTS7PD/BAR8ISlgSe22sd
U+1bqIAifueLczLy+5BLFLW0YDi1qk05FSrYVZc9un1WB1AMovM+El747oNvHmDD
A4EMcqqm6A3YMYk+ZkD3W9f9gfgM/5CW58ia6TaHO05o2I/2hnvbu1PTP1fVhQ0P
5NCyv5lFtAewx5pMNY9rVmC79GVLJ8ebaPNRU+JYv9Av8cM2ZRdfTPCfubhKJ5vb
rNZ5s2YWMlq3cPl2FNrITdRCPtjHVJjFvzDNYDhmWXHdugH8JFzlWyxfXvjrpglR
cEjcXXf5xeK4ayW6876u9k4CI63hI+lpZb3GbOJOM13kZmxopuOrPwpM/3zXiDF/
bRmlmYSD2fD3oHRD9BqRYzOvwGmbYbNq2BwG6eFGMaOe4w+tTRy48XCPND/A9DsF
xHQKJlzEZC/nTUNr+wpCIHTdcdvaNAgzM6reSIoE0MU+97sjLEWcjmwcHPx5E3uv
PdK3e4jy3cgkAj1XdZ76utTIjM4hD/t1E7NfWE1RoF5Zx2RhCqlsL7GXPXI7zg2h
8DyF88pRhn8I/0Wk/678x8i4EXCAjUAFm92dbWmQoLXL9U2W4gV9lILYj6lDUJ/c
H/bp1wyTwA2AkSHGfLp/OMXGXTvlvoyLxHGQ+7ZWkzS6WJgXvoszfr6hcknRUbrw
nCJCrKVVKjp/mrRqoj12tHoj8QaZ1EfDQ+Ar8d2UQQBmhE+QPQ+/nyFrlpIY8Hja
ToobB7YqKWTxMYxhxoev7NvW1NSBsDohkpamprdmjYO4YNw6exzkK0VIBmc6PFJf
JIiS9q+yJQIYxwnVOYbiK4rqba9vRiB/xwfTFjDZvmHQkH+v6nvHc+AqzCTm4k7z
hTNvwdxB2zfsOZCFdwoV39KUzfQdubxEKtNDfsfxevptQWf1VSEygcbn+G0pQsn8
a+Xv7fG73lfMkOFCjVlhr2uUW+WXHQ0VO2x6o2KOKDJswo5k2ZPbgn6WC/EBirsH
tSpu+bQz3iN3fl+ro66B1Ntwd7PjBIhEO9hx5m/FqDc/PzOr+vpC7+Wl3k1FuMFR
pzuvkqsOPZ28UjSfwWZ2XJ5ScbKms4mTrfWfWb0h7UeA/ajJa4ypMug+gjPwbIQb
sNwlTLILfGLZXuZv7n4irlVVXV4YFPQRqmMaJNuzXmijmpNLMiKBTXZOm2jU0oKL
aKStCpD+qbk9rlvDIf/o2w63d8j7JIvjosWnWaDvxDC8+FdJZ7b8lYlRJ22ffLx9
VmPvUtYsFsQ9jrFw0jpcqvc6PS2TkpEfVrbFw7IWXaj8ePU31U0aGSHrC7lWp1bC
sz91MhLt1sUFvip04J0bzFOyhAKPZNI9uhLDRB6B3PFx/b5nOcngJMC0eQfl8Ss/
cdL8vJtkQM39S8QOERxPR9N06SopNcBPVA6Y48DLhhU6OEiibXK26s1A1SOj3W05
4ZD0Jb5Qxd+w4I+ZQtviftY/PTBW7FQMjnfyjmQEksRu/kguLTDXPrPcgZGiEkgD
j+Tgkr0ribedP6ANiPT0H+KAbXicIXnV4uaYPh5j/3rYF1lpfagn+ib/Hf/Blg8v
Z0byA+1dPAAI1O+6EW3tRdSTWIghk4XUlxQe/x9eYJsvoBYXpcQL11zBcokGK5rt
WaLOLnDwOGwlzI4fVaj9s4Kb/NLm7uV3dGhZd7ttZTdnR2jkB9vnnm2iZAchUGJo
+pyLgQN+YvKcFoJj0fdUkVcFG+lfHTaaMjqnR+wro9Uza7gbEoatkNQs0LxEOr/B
JdsYyQTJt6Cl9/hb0KRlHieDn4CbkHyXDw7qqEfVYSEEj11IdCZ1VUczPCC8eAGe
xLrmd4JbUn+Y2oHFa5ikBwQSTviLxb7xut8wVWbkKwwoI7Q1pZgAt2ny4l5fbn2H
aWjk9cLuaNpRd1l2qRAXCptClzecpDlYuAKuJbara9OBmUqhg6Goq0k9q6P/HFp2
oXo8qCW5AQwv6RuRpZ8WwB8KKDquymBgin3es+Z1rE1uHjBh5ksqS0F7hOSNMVMA
WEK2L6nLd4tP9gegE7MbKp4ELOS+cybRR3gNhgkzsELiwzDwT73PZwNcxgo4yHcy
e19bOcN+INY3wkGr4ii8HjU+Y+4+Gvp4uvBQ5n5xohE1GZz2kV+i8fV+oMwX+mqj
XrIxiJW52UrZrwiInewVBMwHVGaL4l/Z9mcrtVYkQp+8IDZrKre+EoueHBJEByMQ
W+6OrQgo5gbRJvvmLmxBPJgGvQQtIkHod798sZiYllCmbpsWt3XzsEET7m5gZ5SF
4FMvqEgJZ11Q2uyRzF/eBkurlSKqqmFSmM8cALUptrI1Hg5aNFEvlqA03z0xiNR+
ckSK507VSQ3XAZC2hwV9ijReOhcimzX2/6ZURJOZRo6kKjpcRfxgUolPqIrEhGIZ
pihwCVvZUbJi0E4y+nXm8kcyRSJDT1AbMfG6oVMMTSsrHrTEqFHGO8ebI94TQij5
Uq5HH/DsQeLVwwyfrGo+JrsXjFhpyp6nscymxTt19Kw/CQwqchyjXe+At+cWtfCu
m80R+8TScvqLP4nkxw4oQJULpjadsbPU7ZFaxJQLQQv6Qe+C1MC09d++NArvbGOv
VPR52SgfxMrbg4O+rug9oop4Q+NhilLwStWkTkblGRZ3e8ykzCqjKkdZd1dWZKqL
lfQYRkTVBBzvIoaiArrUm6j+FBv9kF+nbrefBMZjakLoDUOoc06TaISZytbDOjkp
vCTKjovx81L92A28aYsau2bAyLrPjpz9xR2HRCWPfaBGTHNoi4L9amm/X0HUpyVx
jhYKK2bTyVkcuSeimfAVuuGdw8A2RUxobG+VNFEQ5iCfHRprnb/gDOqK/v2PBxQp
tCImWipB1ihniCxqbsW5hz8wBVmCBBahAQqSwmWBA0A6r/Gh11cH1UAs8goL91Qf
do/3cf8EZFYRNJtMIvpYyPqPlglXN/3Tkl/91hMJCbHg/hmIRkIKNuuGOjNmzydl
xkyss53MKgio16YcsjcOvqjupydKZ0o7OgFgemf+OilQXHU/otD78VLzeBhYOg/u
jN08urVzwYfYQW77x9Rtl6hfcCRpjgNA5k3EJa/PFa1jrmLH2bXZdi9fOZZMQirP
2vLzBN3zgHXgJqg1g18z8F+pb2BXHzBrtJsaC7qYaKu8uHLPaBcMJe1LkC+l9ih9
SGviPNDR++AKj1zZUV7W0ft6GeE4z5VS/5h3kjsEgqF1Ha7q9cpkvZChPHYrQLX4
gjxyn68Ju4qC/lI/qJ9F8XKJfM17Q8b18mw943wT8FKgwtFH2ORHNPov0QEYaAqD
Fb5o7qFCv3m/c03DUwuanWuYrGE89ZgWD+c4oaOwNRxjYFR8bJQfx0pru38lHBBe
Jmo1/FfzkC3cxl5wyH6eihXJsTc1zAvi0qLT6eWqGF3lb6boOo4Pn5eScK+VsP/p
GER/hJLz51WNjrYlw5gL+8Bd4RPe6R6X6Q1CBhpiTjooC9rcJAVqwgRzG+h55+CX
zKDj8iB+DFrOeXCHpSHKbjkc9FLL1XxQtFCaXN3RzviiQriM7Mtmp+PKGJz6A8/Q
28OQR07agpg6/378yUcO0LxdKRtPAstsS8tHrdF67/V1CbowZF7gD7a0yUgo4pXk
eRtuPEwWUv9COrnsF6Hjig7K2lvKqr57uITTMAz381s4YZxrzyjdVCQEWlDCpq7E
8KnAqVFJJbH8Ynu/LO5vqETy1OeQKMTIjG1vQ6o0rfQ3cpu26oqgZAq1dy5h9gqE
qUb6fYpCuWPs2RIO25u8uEIgy+HresXHz9WccLlPJuXt2sqe88uXQKe1AptTyj3S
pUVjl8V4c3cI4jO4vFFfUeJs4nyQSTuicBi5OJd50Ikw99zXl7ZZSf11Au1Xt3YK
iEof5+nCVHJtuBEzVOnWAHvOj/YcGDDu2ummXPU1OcrMdMWsnDq9aLOaQUlvPk/h
qlKhvok9XDtXDFQHI2HqtZeQvsZHfeJbxqSh+RZhUMP/jgTPZbvjfjC2jvH+XX1h
ZkYdRm3lsWjREHZJj08hGYQM3h+mspa/UdxTiApGRCZsuY6LhCrevy328zzPtCQp
fgDns/vk9oCdtkrAmYk7hfvWcs7qHkrligZvdl5tPE//YwNM9R1+uPATHMhnIhJ8
qko7SA++azuOYl6V+/vu9Si5+NO0kLI/NthPwf1fHlAVQCaJ2gOw7GxgqBsWRPCv
QHKtjMCTsaYSm5Ql7l+CANkL5CSH4ITjcc/ygHzELUYBbeNsIft7cHUebAxqeHoR
uuwjQq5hTbDOD0b963Os2vxJhitXWii6P6nLu1IewH/ceFxEKyhE7rdBLjg9AbZg
Qh8OoCo2wkWUrKkxvwVF4gdSO66ZLqjER8ddhW4mZ6fIvXCraWv0EUcTWRFtG4P8
gAoyg78HZjzfi03NHkmm2Y9nQj5AjyhMMi5rNV4KdK3ZEpZDfJYfckBZrWe9gpCb
oSoGv+zrGAPhx6tU+VCGT+yX3wwqu4GgqpY9ve1M7sLjr/2uu0q2r3w6wOAe4Zsz
HJvPULsw2kyHrRnXfS2oyb1ZUWB+9ffd2ErMpphzqh7PbzRLUIf1eNxh62KWFL8/
d3OCMBR+s6d10WxIRej0TIR26299noVXHf3m4LNDYqy0Ydn/4/UGCo8QbTFjFTxY
Aj+lgXzX10y7wI11MVegSOOtuFUNe81Thq+bo/K7XYDqL8cDNbkBp8Uot1CYuaCW
whjPpvcRCWu7pA/ivI9NZum+8XZ/AjpRWj306hs3BgMY6+1RY/n8bEoIP54zoxES
RG2D5PzeVRgBTMIF6v1dEcqB4BVns9GAuDztXWVhXvEoVJ9N6WxNyYiPlfIWkuX8
fysiaxdgsY8AozFzZztJJ4bPs9DSDEg8SfHit1F1jGWww2fcriuXPkLyNRF5q1Jg
GYnnAoKYPmjUMbHlPSJU0GG+oV4NPVARFpra7whSSV9TKIuDAJ7zVW0Zf54RTuRb
XqHQibHPffck6bCB8GeT0n5Zc6UZ9b+RJ018VI7wl0rLrIvTpZ09eObGj6mV2Q8s
ezlZbpHaakAwRNqbPve480e1aIORe1ilxsb2t/fgahvTsiIdouE+Bypoy6AV1BoV
MHXfk3uuKA1vC8G1mmwEAH7fLgZAWh1IF3cKoMqVmXGtvjAMN4uVDyRCN6gKUGy5
d2TplVO4kGbOTnSvGxbHcuVk0JmccHI32Fo35ynxu0oVHPaHZQmB2r9VQfPNvuc5
xzNXo2jsOXevxEz+Q5BPre1PoLzJR2ioCEBMmEklXSqyKyBNu91JNlxJhZXnDipd
0jnQXyopRwJOs3nF77eDKjdrpIfKHdhliYgzcqfTpK4A0EwJ8OvUa01Eg2pw2v3L
b4+3VipcBsbz1bRMy3wIwAux5FJ8oAHge2G3UcOwZF4XgNSr6aH7bP1S5sDfI7yb
XyUwr18vDfYbTtK9vDNV2KHyYHP7xU5T36mD1ip/jmatf4MY1hO4BP/clShEYHON
dn0x3GfL/DLkY61BmH8mS/Yr1/KfiOcK8cSG4tura6h8rTq6aCaogP3NKY07mu87
Nz2rxK3a+zOJzH9Q4X4nnAEVwu5iuoxVyiArGW/JATf5p+2jo7PgUtvuub7rZ6ad
kTQsbu5oVaXjKieeM1Sl3f9g6A8smREJYt6rlVwzxn/6HmrJh2YeieMRlryR2MSK
GnoAmYsEffDpyOOUmmsn2X4iQSWG3H9SZ/IiT1hZXVCMSNzjX53xRXeRcDqcRpgR
fVD9NfE0y87w7MaLoZ8wAxsV4NZunGSD55Tg1NmhhhUuXjFOCQyF8omfTiEaVI4l
z/IFc3EnjQqokM172k1M0sb469Y7rPKBrySLMFpG6zpZd/tG/9vZzwUKP7LTxZn5
a314s+zE4FYGnPVvfnLuFkavG4f9EOeXJz+S/RLrIGB3oS9N/+WXpHdivAz6ieqN
ZUGoIn24zDqH304wnG9qcIzxaFDVwPMqE6OsMIG3ApYX49EmTsGt/Jb9lX9KzZA8
dzuCcsi0h3mOm0eqkvMnfkzXK6Dj38JFtcshq+Is8RqP3uD25ITrqF3L3iOQGnXG
sWxLARnI+kJTfEepIVg7r1kWLaN+9y41KbQI1xGPF7afVIwWV3QudLYh3dqRwWat
ojBtMxyObt2XiYOur1oh4bLBIOjRdvkmL4lcnlOEi7OhliC1goy9gam+EiJ+B+OR
qTtT0bBGQ+Z1WSKdVkvvDA/Iv8Oz0VktcN2GnT7hMsSJ4Ys6LgSPhJhIWskEP2U2
UD2K3TO4JSqeFOq4Ccb8ufpj06/bKjI12NxSVflW/8fZIM1VuOcZpsOxFFRrc+yr
j4KlVFKfhKZCMlrKkQM9GqHibLTuYi+aERgH/IoSAYF+QOU65XQNMF67VOVWGEqG
lP+XgJ5+iUDaU/54AbwH0myvmuxjvn6dDySPfAlzlOAsfFJrvr78wS3w3/AmzjTS
1bjvBbmf0M+9n6EfIQ+kZI7MyzKd3E7ouqzR18wcwbRmR6S/5MpsR+CTMCcK4dgh
7R0wXubaGpV2Usx++POIaj0cGqYdLx8Kw6/pnNnTS0m++VNNAjiaWmmgTjSTaH5p
rifzrCC5QSGsHj97g/67J5/rE9TwAlKDIxGQQ8v+H4DNdRJFmkOZnR15pY/7kMCz
UaIMS9EgvRAmCe76dlv0Ybi77iCSKBOjAwvSYy0a0S0rKpDVXN5Vs3STrm8q9jeu
nJ73twCr14K2BiYRIkP1rXAWFEPzwb0yj7rPn6PmGg2FMmrErHzQk1NldCJdLKMb
3o+xt8rl6heLd3lUcO/DE9y7gRqMj/NOPPnTjVHAR/popIFEWtWMgXUKF/+uX7id
JoQ2v2G8kYTbCxrqP8ZxVShS4UtwMReVquYN0yXa2GLD9fTA2Ew4CcQQUHt+cQvp
yiJT2lkrI612qv/4PI9E7pqrRIyIbsbBvuW3qsX0sLN+Br/Tt93KRGPThQRXJToM
PImDvbIVB1W7XvZ7hqwYuaGpNhoraTBJu8C4DcJK9EXiUH+3aw0fsfFDpedG3Uo0
/nrAostAXLoAK72qQnG3ZlBZ5e+GMRtXJHyqpsYZ33VEGFSgZR/kQgwmkRkoZo3N
CaQtEva7ZRrg91lqIo4cTLKC+Is5XRYwNFMmqNWcHZhFrOneUKNClX4GfaJlER/g
FeI/5fm7vrzzwVFbpD2NLETFHJGTK4hkegayQjTDZLmpdBiSkfg//Za9GCJGS/kI
9ExUX0SGy0YvEVbOmbVcvlGanI/HY4o2RHw8KHZVtEXDucz+ibCPV4GJHR5Og+fV
RClnJvnuWkh07p7QmoC3DmGd+Rdt3YMrIljuCLOQEJbmMqma9vBgnk4x+ZRAa9W/
143dnZw5xJjULQo5BwgBJHTnLhoF5LmO8I02bTUAFMkjXB5tboyvNc/x0a+dNxwN
HMDA8W0/mERf+skit+wV+fjaoN/23F4xs98tY9nX1eSqJu9yQfNJ0+/ac4JgMbTP
KdxbjHH/cAIQaAIhDgtIg8NJt9c9yfh2+Yjvehw8RWHSj/vMf3DMC3aStOjSdJI7
Z8Ioz2WaOPslqJkhcydS005eRXJFhwh1geYwtiX40nFBwToFTdG6pE1v2Qw5K29K
+wKVkFVgCjN1VUAy4SG9vxsqfOp/7aDumAByEnJKw/eb9ydwbv0y1cmq0lwOzETH
cBXbrI2BCQ+AxvFXXE95OzD15pA0ce2ec2KojuNeS7CAUIrX8WcQDFf8AXrGJcfp
eqiP0tIQLQfZEh87Ti8UriOfC5qolTNrvxfnJJgmuYukNiAGkSZR4/L/Ikoa5u86
uTC6giizhOfNyqgCRme9lqBw2/1QQ9XQJHQZpxhH7ydlHILuuH371nfxdEdD8O+f
uo44CPJCczWHzXHxeWQz2T81Ukhj3/Kpg2y+ZHa2A1pn70JCZQ5pseosaMpNhoYU
wdnMFglsge3Dttmirylqj5noJZSX0w1jlN5ll3ZMbL84dsfCp2KKEYV0wcQeTI4l
8A90T6cHxEqypJShj4T2pTFSvQh0zcbUOLG5FgBc93gAepRdez9erOwlv9l12Zj8
+X1Ch8eNOHq2eLgyJwDcaGGeZFpfg656oMH2aU4cpTkwBWt2wDx1on5aYsYDD4x2
YlprZsNKDONuJB7kpx1Ng0PhquudpEgEk4FWZIO+MqGsALLfXCtpxNFxHoZK9B0w
ZMdKsLifKgatc5BsSuJ33MDXH47boF44UddsiRRHXR9ObG9eI4OYc6qfES1xv41Z
5FlUwDLYSM7i9iEb/phxdi0b4qvrSiDBePUZCpNciOUZgjojB/GRvuQVRdV/BZy3
Nyl93CUFUrF7b3op9wwnvOWPM0ndDFuVAbuE3j5aILSCuPKXpEuaD9QyPr4C1mrP
u8kDRM9rTOLTyckegS5SaymU5f53dGlpCLH4/pAeWQhtZuGHQguBsCr4W99Uq2dF
R03v9p44eHYKpF0lF+kfw+0AdXizTrxlRJZ9AWZVmTDs30HZDKl9y4rDTM2yhuOA
Rfl+I+HKMlj+eRT+dyKia+zzu9kS00cA6BW5nfq6mc3Qp9udUNbUxuZ4oeQ8YGnu
tW91p+wNS8a8TX8Whms0wRki73wcxnSQG0SkEqzqQu2KAxb66pxgKQLaF3WUuHsJ
B8mhXgh5JJp1gNL2aAflrzzAE5LuNYKkj1o31uAG9R/fFl9RQGeJ9aU+BSaEwp83
v3MNTbsdwAN55S7vdzgqFbAudH1BmhslE+2ZmTpG22+Xi1xpZDJ+GssnLusItpJA
y/8XEOlkiZcZz/GV8uSRSbW3Xe9qwqdJQZWqmJj032evJfJdt6PMRp0fLNTDoE/3
4ZncSBS3WraQgZx9F5poGwVP+iLSRxNR17/f2z1vY6qynG/ZzXI+OBg2dmc4CfCS
rdOaf0spURGL4DdtohxNof7wPnQ4T3qSef5C/hN+RcVwyRIBeCt24tx3qNWuMJ4Z
9cEcuE4cnRSvDsOJ3SU6pcoIwC6Bix3lQd49D4V1XpgGb9Kh5H1OO+zxRoIhV5/O
CIXEXUmUTH21OFyKDfGQu7ZL/WS1LspOSOVDLoU2DJBSlw6tRQdT3Y2gigkJvK0E
pR5gA+iuXfZwxwO/4FZI/Ly/iKhvFhjBCD88EQM7pvIaY0uszC6fOu2uRbp6wuzr
azi023N2vCUjU68yTqO8cV84l52LPAFJjVKcTSJlruGwXLB5bTx/9cSFf7y17wa1
XnqNEmEuDD2LC/tfzeJsghi4ryI44B08l9O9Hg5AqUX2vUbsXvujS8OcWFFeITTi
jXxP5edaE8HyG3/dil6/tMQOClz+A8knarmVt52MFgPrShLtia7Q1t5xgg6njy8y
v96SOutcC5S77sSjXoveXtIJYia7sQ3+94fwzc7/7S3sqX2aQKkjh9mJ1vsjZ6w/
UYQU6VNaoU2m9cs1HRJiXNS9gnJB1bf+NUXj1qq/vvRYiVeKxmZHvnX4cGRR3CHd
ZYTJRM8vcOjHJvIhNcPHVEsAa07MhTVt4yJh8k93NHNFt702gxEIyTrINOXK4YR/
MVyT6BJ5sydf+7+g3of6XhopnPZUww2fM0dNcXQpixviU2NobtU712qwGPzMj6hy
UISJG/IlgJ0dz0IxBeyL7a99E1Qk4uLNJGPH6QTJcfe9JQL8/Psh7zUIZWuZSG4D
VQ0ekbCCgIM68Vpa8BlYBrTrw7FYKZx2UTrQdQOq9+Db6lR2fndBT1HZzYCRa0Nr
lpRAnL5Tt+zpeTzcbo6hwan0+Fk3m6h94Hjj4ct39oHZ0mn102qQXhrIDPjluflp
BF6lHgBHeXfU2JP0DHXytEfDs599PKTeebiH92iSeT2ITko9yav0Mw5BYPzynikA
iMQqJTA0SCEpAc6SORqh+Aux1Z7wwo8cX8shl/gdG+1mlkTiLv1fYFhFMN2EZLTl
wefK5olh3onqRuP75DIRfPeR+TH1QIZahy9EvfkulDePqK5/IrbNg6SEKydX8ELN
CcF2TxIKhGC+RhWFO9/DCJTWzgA1BE4oWT0cHAYHjLu9nqc6kBjZd6U5w+aVqrAm
PgwEqnsrgDLbkSQi+tFVwplCcFzFivNJj98uRcw8OQRZ1/LM+Tz8JZz0sw15+trR
hOXLcOwdXx0U4Wy+lAlgKB6/FdbAKXhWdR9NLwtkMbQTCs7BaZ//3blyP2MeTCYV
33Z8X7AMzVoPMZHtohAy2TX9MoxRLt7y9E5mPYdZCS1Yu2k6pzEUewdbqtDJoULt
PD1jpYAoIQhjE3JIuC9N++7n+2xqzNd5udw1xnR5ce3K1OU4u3ObmQrk85KZyACq
1ZuZ9/vlqWeTgohR46QviIhbcg3pW/ZHGk8w8HFbH98O5i8UI2jUGa9umtYvP3Q6
x5kcLmCRxumzVE2axL3raR9AQB7FlJaX4B6r8ZuCYksPRwaPY0fcX5VzfdAAXza4
gZj+F0AeVAb1ygwWLxvc5W52gpLkC4CXBNeyGoJz12fwPyUhfJQB71WsxupzVi4k
qlKv4FEZFr3w+vXdWD6/XRsDfk1uHczpR5eiFkVmp/Krc02bjGp4KHdI2uKXV99R
50c5EM5bRjCXuXKWiSuU4v+WBrvMq75NDnbgNUL2HQl6VFnSa67PLvAOOO3UdvC8
eXS18hxR1FqIduPvdZoPqZXFDQc/KIoe3MsbeDDqOmPbw7GyCtY0AUzwM5pR4dMn
qeqS/ez0vRYH9s9gA/R6yhhc6acj0ta0phKYf9civkzGTJIhaHui8o7AhfUO85Fu
ntFp3yrO0BSXrKZakbvYnXTqnZyUwU/NxCDVKh5E+m5DNexoI7BknB7ZvpeypHks
dxp8F3CqFHJy5ZzNYpj8RsGcgiyKH+Zj6/uFF0INdDmgsf/gCExnErXCmGe1DjLZ
gyWjPDJpIafGIxR6y+n4zln7bMEVhsSThbNUL1r6ZVa94ANYqb6PVeu38PRp+P/y
b7XMvsVExe7JCTOzMt5sLOZ2q4KvDLLjOqzUJnTqTc6Gj9763easyRr2XbYStk94
fRvSnj/hgPApxTUMZnAgoteEoUVUKRmNvXgB57kmAT4FuqKzXPFgOdErDp9lw8PJ
jB2lNMc3zBRmWUzBC5orwv2LeqyAyVfqj5+GMuqaVApwlTsuZqOFtZycDuZB3TYz
aAUeGgw7zWHRCpliAbIkkwLfKo+//PRC8EVE6hGFuhfMft2M63DkRrt7tonkvKQM
u4PrS2xHiL+gqEW+Gcu64++rDKxCDLjjbjOQkT2Tppxp9RZvjQmtfx2jag/qteAx
1mRa9scem1QpjqUFV0+coouxqvGjbcRPkd8U6A0lD4uBGZ0ZGzsTytzJfqWHjTmM
WMRnD9WwNGmnWRL1EdwPhsC16WfZ6rNU4WRxdILXsyWW+19plkLcgaDVk2AxXWgO
Z92/PUXW5058nsz48hNWLsMosfYclKncqmEIxWfj9O5mBh6kC54eBnL7qJ5PxXMj
E54sxyHNrM5tJAGsIMd5tfKqcMGnQ6aFBnch5G8Sz/VLZkpB+RiMDzSZycj7f1Ib
jwmBDR5X3EbDg9lStwp3vw0E09Of9ovnS5hwAjBJOm0uV20nHdch8BPj2Isime+v
XXaKxpNGdMk70LxMl+yYO1a6kGmLVvCaiwLkCfRFqMWRnv3yALY2vWPooxIkExg5
gdgv+ZWwCxi/zDBRowJmfiB458nML+gl/SwfAEIQ9oy3aLvgqymWMWCp4FVB32lY
iwtOxJPDP9fCdocr0amG5yV/toY4ko3W5T+vnJA0XJkQdn7RN9iGEmcSdBOgNC2q
P/j7mtUTMh7Ae0GGmRUMWfSDzA/hkt4iP5t2xmZlWyQLBphspngb91W/KEl68l6j
rqygojwrIshyU/MsJj7AZ0qQmAEMnSoqEo0qvDUc+prG0+6uvB2iPv0vGNd3Z6CQ
UlKWUfKqBCMpZC85Ey4QXNM8IcWBTeJ9GW/QZmIcTYxE00LkoyPlx2FTYiXmHilI
N1Aoe2IvLBNBrTYIuFlxF5OU6ck6eSQJFfqESLXo88Oplxcm40RLs/Yzi05mGwFW
gDdFeeWEOcav0o5bQl4uFS2FfHy9Zz9QFwiRQYJxrdFbZd6NGnZILVc92kf4gfQH
b3OFSkPmfryic57vhxexvIOx57UKSXdLi13YcFG4g7VlIsEUNuXhqYqX+xQYbYDV
hBSoFHmEXXWVaoBsgAYpgt/WSOVTCq39hyE11n2QjjxlHzagSZZL53gEXPwGyLxN
J+KW1zAQIfHE+j2wVCMer56U9iDwdsWJiJvw6JXuoxCfXWMBGL10t4RBPB9D1yv+
6u3B+lL7cEYU7oLhIpR4UBVpBG64bEosjk5fjsb+jNdqd91eA1gWolEAbbECv37+
FOiMUtuT79mY5TuQHuDNst9+qKXel9d7PC9VizaI2Rsvuk7DeIJaUQ+SGoHO9nHu
52CPPCkS9YU04xVmi6PaE7EKOgOtQop8OcmyViAgGurpVA+gwrAPIMiUMWZsGf/t
3wCwcuyRx0pKWRQ/ZuH2nhq+/XRYw2ytvXOpXrUxT+JItv6baUZmdVLXG8W7OT8v
/tzHfQKtbKmSoKgoWTOE7/XKie48icxFnYLUx5f00VMWdHir1ErkF1SWeujPO4Sj
565skDWYEQkwNQkoNU4pUWGSJsDN8jAH1tJrgiXRoT13Lm/uc4N7nYtOHZ1ndbBL
LEGcOy6ey8oeeNLYm02/CMWfR1QmhrjmnHzgppXuNkXrMeB+wPIFmzh1TjtTzrMw
mEMFBQR9llTVdkrB3NeGMevBvs8/DNHR/yrezcpF80EwqZNy0kd5hiBZL37SLBVw
E+gId+pTNTK8X1ddx9qtI6ssx0qxQShkA9vlkKvSpqzDQcKNvEFQhaDpP9Tv84eY
iakI7Ls/xx2TdOnKKbCMiBA8OQobU6I98y3gRJa+GoRn1iAGb06qmd5nJNCQ/Hus
m1jrFxZYgXphc5AIT3dbvfkahWyenhI9vhCJG85GgTxizX63/UA0yVumrjt/3nIn
69GGopGKP+OHnxlCVyaIz8RGUYcmYqaVfD6ElUbntweopK2iFVl7ajYsqz9AMD1/
DAYN5ZaEcH4cAu4PTHLYA5NHzNapqQ6DyKUNOKcz3YwCJlmBhKbHDqdDHmrI4Rc1
23Jn1f+C2lwelg47AYTwAblMjGhz/os0qHyDumnt/2eNyklb+TeLznxOK5/7OZGJ
Mw916y+rlff3d6DwQpeuOp63BLXzQRu9V+Nv8Jf0Wao0D4cccqVoaYwSgC++i+IQ
PpDbRK6hNb/f80GaoEElzYuwfKCs2vXiAfjDVxxBrwtRlDxGWG0B8vaZDVKngU5t
/LCtNzhe+N6g2HwOYjkFzAexRTv51EykwZVqsvMrpQJWS2SD6dUp9yVcpdu4cgC4
/VH6vc56Gm2ZuLMdk68UcxDDMQcuGjLMALBFyauRIg8nhVFq5IjUE6drB8tDXwvw
lUCmMETA/fntSU0s55AEZ77dpmLSjGPs8S5DEkMkDeeErkZ3hQ9SZUoY9wX2mqAC
ELMzior+pVFWbOw1iSF2HphTU0/COAEbkixlcE25XFZPVJ7jt6xeD3QPjJLR5xJk
H8mIV0BwccOMfMyPKdl0AQQLzoGWpJ6s/+QuH5luOTTR0+fUyJ/Ued0Jxh4C3PWF
jjhtqOxbYhduqZPsqX9vzExbCi43Iurnnps+kuUkvWeyWATSSQTEmxFuDw/bmyFv
Z7YRzyJujiG2Yeg/pZcc/e1TicScTKQ2EeeqpVClJghCxMlTiJ4X+bk4jkVpiWKd
DwTJRG0AyQN0kLAQmhWHce5g6rHQFyJbGl9qqLhdc+UeLT0N1o4/tGIl8jBIpog1
JYab0z5E7usOG+KiOhp36SYQkOtlyBvCwkuhm5smrwnu3gPqKpqXt2Av+lm9NhWU
vS2Acl98RfT+8qdNEo7ScT41k13ndptU77/GYhona7LbU0KZNZ5M4m5IzkfUXvrP
W4uKYbXcYVRNT8BLC+fjoxwprNyL+0X1qhcLqh3pg4WILOvqG4Zn/1KJHl2BAyMI
rN30n7d24cwPkndCNjBDuW1F9Bz+ode1A2YzImKlPzUWui2hCl9SefaZnurfxHXN
YDfr3pv9CgwonXuT8u22R7czr2mdKEzo61NcRBdf/Xn4hzbZD4JvvWlTOjmwjVLW
983O2daT19iIvQARfnNmv4BjEL6/GpYn+lePc07BCtC9tNM2W/MR6VOzVuW9k4hf
JDK6Hpm9v6SbOnCimGLFyU2uLeZZCEsOuSOBOyNVsXG7iQRFkdEy6FZF9l126f4E
chJRAovZLpVTqVSdVd2HAFAhgFmgiAEBqJZsFPhs84LyWMLsMs+rf1vL3lrJEKB4
nwHQYEK9IJKOvOl53GUFw2vvr0PFnQfeIKCjvdzDhQaCa3HuccN81gRzyi6wAAyV
nyKR/QpOTzDrTG5V3/Ze7e0twCfzDZysHr39CLsvvYUzfRzdr8FuikKvJCeYmcpO
2QV/LaNrH1l2xQ9mjr+9YdM/ibfWYXoxFbrQdHSblZccUfmRr+9YdEcCdmJ6UXQ7
vLhRdsJCubb6FYP358NzDbjwQqMKr2Jkkgm/en9x0swox2T3s1f0iyALYasxo/KM
xTQrqxAWqwxNKs24BPlvcUerf29g+7L6FZEvWQ7dUi2AOv59Jri9ESBe/pTog7E6
CWIIA99Kbf5Z+JKC2dAt0JWipEz0sS9SRGbOfsOeXMe4s506lIqSkE9WTVZS/fNL
dfuVGtW4F1MiqIvuEJg73SkMNCDyXxfghWTQwn1R5Fh/YtiPyM26uo/z5cj3+LaW
S4F/LSJ6I13wR/Of7lWCphn95kZWmIJEX7PrgESHG04FdAPALxTQ40bP8Chqemag
raNsJNlApl8iPCM/gJDAPLr2NQS0F2dwVYpAEpU0djpOxB/LZ0Mwpy9i8rfquLRA
CgMgyUWeNXhhZMlt6tE9JlEJxfoUTgnq3K0DZ8V3OnLohukK1HTC4/xiv/L4Ua6i
PukJNevRqVNBSnLLd+x+yM3nfohCKcqFT80uDYsAt3WxjOvhmmMk0D4PcIA+nP8F
z11z2j0VQYGpOEdZtMh1nXY+1cMp2QKlsHyaIxH49yjF83D6vcOcBWQxBwkMa7hd
FpaHPax7fxtrH0NpTHCOGVda1ZinlfJKyScxFWa3Q8G4ZM+3aqjb3Me3Ym21AC6S
0yxuedu8vuVvRKnUd0/JpbAuDtUC95TRutWCth+hPy8Ufj87G5qKcah3+X98BjAW
iJhFTWM/lkXqKusUd7lAY7Akr4cgRUzY0PMBDAc9hkEy1EgmCHOPvJxu6Cn/eacW
YDjx3m1nT79a26TtLJ2hV760tfHiaZ/6sQxrdWjdfKEz7lAIu//5qnynMr+ym9VC
JuWj/JbWKJ+edb2w0jIUFgiwVVpDOLYmMjXlMIfFO2Nxp7VfU+Wldtln+N8iDjmc
BYtD/FcQFyt1mRdhD8dRcCVYl41JH5lvW+/iwgfykRTglOFfI9gG3CGRZlKwE6Uo
fijWjDSWHJg41ckGHqeBsBlj7ybvWyeHjI0x8uT3+3wjv1BbHrg2zEB+FScKAGpY
cV3IVXOxmnQcDd1jPyywi+t076NoikomXYL4TypA+20aDEhjsmGocAqkmoaeqBg3
oWSWloNqWCkFyICWP9Mtijbmbx7sPVwNABxznSC9BZjEafQCI0d1ohL+SN17jpmZ
peHL3O2HtqFeZ9umT7nRJu2Oh1cG1hTNT1dMHyOC+HHcCa9xvBh6RVWDkCHLJ/5N
LhMsgqDCvAPKuq/JN5ivJdBMgKEVy3PqKPbbcm87F3r7L4sKdpKbleouWEI+aK8o
bnfudDBZIUT3etOBLzDPfK9EkKZSycbnKSNRjT8FqobcqOEVw6nSY/gKAQkzmrUC
gfxOErOeLX3fVmSQGmSN8l6ptQugYpVdfiOSWa7A75MwToK+Eq510f/P9+i52vml
NCnjbLggFZcgQkbRmWG3xK/v6cxc37iZiA+4VmRzMpMWM56OsyYKOyM+78Bv3w88
7zwYoI+5CsKDX40bYMOYHeOlhtRztepjSIprGocHDN4rJBMEqqvdT1BjyUeh5SYK
xGjSkXTpcnxXqFI1jtP4uM+NCldiFzBoN0pCaQnqyGCTZ1yGPsyWZF4qllityb8/
ctQa8awTMSf0e7WPcQFRH5JBpo/keDZa4d+HDdogYpTvmN20CVJxgqlzWaK3wEKp
YMLQn/FxFB2gEbMTaVOxV10mPe7Qq7avVd48n5c0UJj77BOZO7+CU7DD02wYiI93
5j29UemYf0nH4Etq1ardEh2hUjt3/MTqrCVEviBJt2ku6+k0BiTMmxKcj/t8aUr1
bzWrj6fUbDqLT+Z7145NXd1U6aVQaaQxT8cFph/Irg12zDD1LTi1zJi3CqlFwzVU
wnVhl1IzoLRP7DCmEwT3J75z8KJ+CsOtOSmix8Gx1OstY1bir+YKPcHL9suMsymO
6giEwzqi5x43yAlrdxPUdhL8ZjUopIe8D/FWjpVKEng3Ic3Jr6HvxRAzxfEUMin5
XR2JkolbuEPY9RpJZGyJMjAZgpd7y8LG09hFgU9GSggVZRxMqnoXQny21DPVmnHT
Y9Ig0kCTFi5xLzvhjGiLOLCZ160+UPCeSAxrWPrcKg04wD0eMcR5MRyy/VaN2dC1
7R5z4om7ju98CPtRDU2ElQfiaUCH+nnqxdqJFA+8QE6d22Hu9Yg7RlT6zwycdQD+
Ie8c4O4rRKyH7HqaaFcH15ISv+KjO//Sb0pLmohx0KaWReMf1bAj5tP31whD43nT
2A+hTZpVScEdY1WX7vSTqQvdZJu12DrMQ8zDRKU8cLf7llgIqlgAdS1n8kYkm32G
8WCry50qEvhkTr4rlwx6u2BOKfDvsnBDTi78fBibXdcDNOmSqxMoeqNID/PNwiy3
tAKZewcRWv21CKsaJGM4NxsjPlpjYWgqVrZnhB4oovPtTk8dftpb+d5ZMv8+lnH/
TDJDUxh4PQayks+FUZhU1ggULYNM/lSmJLAGy6lL8YCSEl9deyvLJBi0dwXfcF2Y
3v69X2lfab6DIcWe0P7NvcHpq+Kk7OMnEE3kv+sT2tPz4I4ya9c9GYCzjvW72F5e
PuelXQ2iYsVsKgSBTMi6BzNOUFzdqiSRj1BNs4yS4Q769Csb8BqTGCjzhTZG1RsN
+K9T9udd53ZuOZdJOfopgM0Wkm/uGgyA8u5y1IQW2eBQ065nqVBRiy5CPcVPTMSm
ijqgRHFfrW2XR+0MT6eM1jwaeT1u1YLL3EmRuX9K8clv2u6vl+G+uNBW0eME/of1
QHn3pxeSuirdvuhjZVbMD4wlNVKlNeXPWf6JUI6mOzWv/0Z5PSYFohgWV8H549MT
mC0ZrSCJ42g8gMFZH4N2wCAjIYaMyJoiZkZdI+DXcJcP8QG9YEVoJY5+lxxm5cZd
4T06BHGx5WtsmVi/gp/GLeP8b+WQbz3RudVA+I4rC7PH2ishtHBwFiFv2tgkEIm/
YCpQdldkyuBzksht8EWTTYHoTJAGYoJHvlKkevcECRWCdeqFutAeZ92ja8qBXij2
xcO2qqWuBl3l3eajlzMCmFFbbisQ1DV5IffVj5jA6TZu5Pz52UG0uvwpKxugxYtS
3ZE4CQ62XTQRxOyvMCDkq93tSTdBRgu7GhtL7ipkT2TTevdvq4Uyvah9b4LYhNLY
RyBqL17jDtIt3YToWk1ROcGlPh7lc/hgCw3yYcq/3xwFjEjbSYzOpTzt2PMCjZl/
7daB5t1dmLrxClW1OfDPp4JTKa+sbqaFggIVqdRVwPh6sbtOdmPOnNcQ3wcDpOy0
GfaTeUA/e8ItPNy6IGNQDruyAp1YbDGX5E9iMgF702oClQKvwlc6bFJ8YF34imIK
bq1sefkcTC2wh/FAB74IGtX9jK7v3zRGpAC/2vh6HGxjWx+336o2B4QI/5UboREj
13HvdGvNdWbOq0cIEeGJpbXyRIrUd3IDKhEhYYeQwekn5AsSKY85gWmIMj9OpExb
DyUEgEz76hG3PocsylhldsO+6TyrHN3hU2FtouIwwkTGfMsAPuL0Ph3QPtccnIqE
zmCCYYdGxK6Hbw7mzgyr1u/0PvMPKo/7Lr2lMIJ2SBMfMeEM+uBfT5hA6NbZmVle
TDdHOgONOfFwiQRs5YvBw2GTIZK/5SR3rBDkpfqWwVD8YKnd8ctxfUPosxzGhR7q
9CP5UKgmnPWinUut9I+3bkvdYAxRfL6bBj7UvLo8vIjJUm5r+xtrYzmciJ3JU2HA
6d1UgC6vyz8iSu5SPjcRpNOPa34sqBUfwxXw/4j5f4MM4QrdzCnVvzCsFXXHMFZP
iBz9x4DD+khK6c7a6p1KRgivvy4VrQFFIXsqrSXFLND73cH+NXPdulxOWpn2BgW0
x/L42IG4OcZyCUm9ns8TvQKtahFSOSl2KxFOHZ7wnkMieeMx396uvFrll977l1XC
bdM4r0QDqn4h1r1li4H7RUfvVb9s1f493Aj/BkM0JeYTUARnkcqJVcfKXAOxcnj6
EBgnmY/3gT74Wn8cDjqsnJe+6gwgjw0K+FS4Kzze/05iSSO8yXGTesvANq7hdCte
2YjE2ehdgyNWQvlVelhGRKuJTdddCH/LgAqw/n3H5NV7P8f57QmZAyFcuq1OrGmr
HNvFzE4DENrIMfYr1SgdiPRf7P2FvsR8NYYM4AKgFH6R/nAd7g0fR1w4x7SMg0hb
F1Kh0mJ+5TZFBJSDGU4PBTdt0nL6LZQBUfJA621T36+OJhSBJvDLUXnYY1ME6Ayo
GPbAzZvRj5Nl6WfI47G2WgvuagQHUXFNElbOerCpycKq+OVEBZufwu+rVwDY72Lv
1/vDaDLbdUUh67TZ0IYTBHYzGBdh2pr5EvSFehCOwxG2qhGqhnAgaXn+NKZKRsYn
ZlP998f7RF7mhIWFCtfGOmwSL3TluenKDgVPn0a226XLv+BRvpXE+ldeQMNdYjtI
G6Gp7i2q/y/LWEusH4odC0rqlJ6VmwU1dJLAlgPMELFhHe2L7i8oIb0gf3TWmX3f
5JCsUDphpX9FHWp8KfFt0bS8jboB4LQz/ObiUjsisW4vgTQC5QiNJW0XCUfhFqAc
EjIUCoNG0rzxgsvwFu3f9Jsb3PiXPPssi2XRPh5ffLGdCJIupATuWifVaPvcqVZf
NiUWMLvAUl8lhF+F9iCrluMSCZAsBYr8cdp3DxTX4yndJy94IiYyx+QRoaVe9O17
nTLX56UaCOm+idqLo+9FXyA69JBapRFW/PR23lfXu7Mjpwu2WjQZ0iROl7Z+iw+3
bXpRNuNoVmj2cuQyxuC453LZcskiSBLdYl3kFQfag4QtdN1NOjMFjUQjGChnPWrp
Jrl8MFcyFAjfXf83W84lpjMOOHJao9FB0nJSi4QJiE4lQK/lBFziikidlSXdctY6
3eG89ixMc9FwxWiyrMKC1ZnDzS4OhcFVe3yPi1uybCREyzi9IMPfVSdQ70xDXGQs
Oexm5Pie0+bB6v1ljCvXV2THl1yq54IkYkgTVtjNM2EGsysD2po78FGMUAatcttO
7nT7TEaTNuVTTNhsp+/3RsMXmEZZG3IWVKnaCdZ1jXIxb1B3nRvWw8SgdWkCyJx4
3NHdAdDFWMl8r5x2TQ5gksHPGZfxAN6HcWltCqLPwKrrqen8VduE6lGl0BgB44NG
URz/QksifAw4Hp5e3tCInhkt/KqC9bM2lIwNRwkJYr0SFdYNJyDxFfgz6Etg/VkU
MNuWz1M4J4gD9TF9dE7urpuVjhYEOrPo4evhscbSpEAQhyzwT7mmjvCf+Bj1yKix
+su41a/OSbcXmZ/mgrwE6y+RaSE7hCTD3qVTbCaHRV5bpSTEVq9hcEBck+pXrbz8
kE6KuODvkkh/TjrS9lKdosnKLBZk4nUfcjrWMt8cWmsEvdzzFwLkjePPuLjAi9LE
4tdC6vfGEQqXA0r7v4nobVugEy47IhG2lemr58RBJF+Zm5POg4offDC1B5trhuB5
wUTVdhV3rjrJmIJOo9VhHf8GUFKxqzrxHan0eH+utnOwETXjZcpZjX/y17NAfMZf
pK0A3FovQFw39SZ7dHz0XUNe/5CB8xETHAlFpa6htKCaQvImVUV5tcyzQedLP07y
gptJ9bJ/LApPWmLAzU1KQBOMdnahVGHjcRC0WM8h63KSnLUNJ0KuNQJAD9GA5jFj
VeyN4H+ZSOkV9Csgg0Qnm6FpG2QkuoXfgw6A0dn8s7kSd6ZFhGFir9iPZQuhB1gb
zPRoAkcG2H5PhAMj1CcSWsj5Q7bqx6j8FNwjDrkps9Bcp8uusiXwVkakM6dN/ej+
6xvwTbYzxraQawFjZqPPK0fPlulICMtQA725xNTkWfAdaLLxsuDRLNc5jBuVSdtj
G7uTm3ZxVlUmCCQarD6ME+lmLBpeaboapJ75qNilsLPfnx3jGhVlU2ZIQfgrSOnb
uy2WqiMnibASh/3cLZS8nP2TJCFZmwjIsjt1jPhqLO6p01NVlpBQJqZn4XVLk1Bc
GyP7yJ08VfdL8N20ojQnY0WqfjvP4y2DKMFUE/B0mnvi+yk705wpiX7Nyk92UZR7
OmOKMKx2pI31fKezLvDRlHXztDGSPzcIxieSSJNj1t4v82Pp6MkpRtHaSr94RS2G
APGaY+cHQRR0EBqSpD4bR4elUnh8hRNPp9ABVcmcZpVHjJ7kjYNJrAPOXo2MthT4
iDSZNH7LNXfE9MPq/o2RoScoAnHAFK9CBF1Oq7drUZ5fFkBAyT+3InxDjwGz2B8g
fosQz2d9C3rKlwhYUXGlOMQx7UL7BAM68RZZJS9vaO9D87ppDtfvzflAraDmkIcL
3I/AfmoE6Si4IPfZ86XuKgCuz9cwb9EVMpFATnsZ9soKvkEPLBCUPNqCVdo8jA37
9hhPx0mRKb2Va2+/ZFKEWFCt/BxXbCWo/8RsHW9cufoYjARVFOdEUorFHR7ycBS9
ZqpQiKj1PcDKkGwBr0TQWAl9hv+D9Sw72TawGV1sktW1B13EFKiIf7tNDy54YYvA
NKfnb+et7pLQtNztx6ysyl5+1ssx1d955olw60gOFAAK+WGgTF9N/Fvm7xa0sceL
eFOk72CjCTksYb1oj+vOEktKfTJcjYDUbZ65/IMUcDuUReaVBwHm67byW3zdJKG9
1OS0j4lcFBPeihv4mWUbMrhbxsZUv4ze0UHJ4o9UEuLmDCBzcsO3JWn2kiMmmdfL
dTX8lWcCOkYUqGsZm6zBOEZ1rlX9YXh1UwmTebNr687cZ09l9SiptQGXTSjrgWuF
sg/ExgBePSfXIIzExNWEaX3/YSZD9D5gRtRyppLsk/6tCd8uOu9iPB4riFiqnimg
PjybOVw4X4RowUJeKYsj38r32OXtjp1/Res8CDkUPm0K0sdO1QiW+1aIcjmbMQIU
oacNd2pkHgsnxIpyJF2LJ3XHSM89JD23d7vZaK+Fe41fSDbc71CgGyZXPaYKVIy5
Aj/iFHSL0gLTbe7sXGAi8kskv4TyUtehRUlJn7uqci1kX7iw+MNNzNI3Q7QU2Xgy
+SK/fnlHBC40oy+XU/o/RYiktUlKfLgGpaI37AJoNSgk2JsRSYu5MXeFwAp/PRc9
O0NXN2QdfCtlr/NxFIanBvM3PPrMkDqUSwibAWdOR/3TlQ+gAojTsMep5QMhcqjx
1/PRVuOWtgnXwcnWlRWZ1Q5myMBB4zAa0Bnqto6li4UWMzOgQk696OHl58PjkGZe
KN98KzHMwpE/zVp+bhXIfe90SyuXMDSrD9pLDy0CLIm9QUyy2fgxG2CBCYsHpGOK
RlrPMYt4Wihrck0ucchHT1GYFq52tLMRiq3jz7uGTsOjZ4IW+DxSd4AupPRSy8po
QfO+f/imMO37vY1yhEyhr5FOgqRY1RzFurzK4O0f3nM1vf6ypf8LWm6Vc7wXBux4
i06XSmc2Mr5UISi3Wmt0d90/Cz3pIVH/xgJQLBTVObpflC3YYKbyOA0kUAdaViON
ryaKk0kM/b/jmXP2kxoZMBH2iIKajvDRh9u6RY5Z89cLJkb9JJ/lE6G0f4I/gZkT
4oHe8n3/GTmGZer/gLuXhTRS1u1f2Qo3DInwQZ3OMwXS8CTGVP0mI809Aa3Tj7e9
eLFe+rssqiANaGpWPeBjawdfBrhZoV1xyy56tFSYnZsmJgrKgCzIripzVCbF3inI
HAgg3sahoysnziniAPjtIf6Pg7kYNAdl9XGFJbKUMZ8uLPyFmxCwyECkyp0/8YSE
a6a+EXix1I4bAaY9bj3yBr+bUOrDDdKQJoaRas+a6gOBdJ4xyR84ILex+uPzCY3e
g/OPt17jXsBn9AvFrlMsx2a4J5V6wJtrZebJz1uMVsLIQx/OM8WXqVQJ2XSJzoss
eVUL5JzeZRdEtqFfLNtF6i6atKsujCzlMu+czrbkWO0cITCXf+Kuu5PmMIWN3eua
RhAOT8aAc0dn7yqw2EvWpwEyk2dUtj7EGThONDn6y413ssuHHdtguEdBclL2hfzQ
u75kI+VjLSUUZLMuCrdWVd7W86xr1V+GFPlY5vX+DFSbBKlIe5apOnJsK5FWJA5f
Sr8b4r+hK/9+8yt0NBAt43Qi1M922CM0yZClW9tTYFvUtXm/f36YRBOPs30wJ+GU
cy0viwPyVZ7YqrPsqBqdlwBzXY9ICHxjB0qtkAMNa/CQPSv76azMwWjCnsxXDUEK
gXERV70GWWDDHZQliZSKAnL+Ii6NP+x8WbQNhfTDDgUVkCLcCUeVwxkjrDX4GAD5
uUJz1qYfVhrVZR+nSrdkeREdn4TtlLCq6vd7fOQjxByGL7pvZtypAjXZPzHQEPp2
bJN0WwOgci7w6KEYxzRFC6ADx+oX9H8bOR+JDv0cZk6UZuVrRN/RiGtlEGIiQPof
uetcrjw6niUoQxHep3w1lf5QLtTKtwfs5eZS8gAODQVTrZb92Y/DDUZKt4IcgvSo
EIgDsCDupcfN16JaYeEwo+MRy2AsLMbRATj+3/dLcXF3yKsWPi6TiCLYmo6srqJ9
d6svvdoVnEwgp0DQIkmuNFbKFSrAsAyDMi8zkEcG/ti9GG9Ie3Iq3xxTDK9DVutO
IZhQIZlNnf/TtyRe8oMWShWVwe4sI/vX/4hmJz/QPRdo3RwfkyglCSc1/cHRegDg
LUAcAl47MOZls/iI9k0jSbfdcuxOs1zm5kJS3kUlvvgFNLQ3LutAg4NsQp5Be4Pc
oT3VE/iCedSLmSnDsP/HE0nQpznm+asS/70UpHoL6Fk9BCtONDVxFlAQ1a7xK7jL
/7egc+zvY2LMb+UmSjmvXeufEQNPlZsj8MKGcAORow1DufxMmkSf9LfoQDVgQuSR
ykys2qDq4j2OsGhboPnbLw5gdWYTGpeLozcN0jglRcj0uzzHo+UcH6UioGLXe3R7
fHBaO6Dus8gD10nIbWmJf+gsbe5G6j3vZFQJsT8hE7ZLmH8IB1WPefL9cCm//cc/
68BdS+X6os+XNoxO2O7dg78Apg/QbM4eWyuCrq7C+9wPujSUVvtSwec9ohr8plMm
IO36bsun49SLA+WRpPQv8l3LAf5LoY8xwzJyn+CPtaIdb6ACzQhFqWDtdRWbHmWA
XdQ1jW6Wz4AoNPrVM37uokINnDKSYZ7SFl5hDiqfpNCsc9FDirJ2o4D+HDAFvNAr
nanT3qxV++olKI38hyiTJHC40MgapOwgwwEypNrNRYZURGdGP0ra6hPe5hgwGwOl
xFMs5Pv/f8pQwYFDjToZi1W4bGe05z5SI2nG3vVX6ByjZpOs44TNqHa+rzUAXBB/
CpzX9i/0bBoJXPLzzS0yXal8z6uNyTBVwKGYMfqu2s4DSq94D/5SpxCyGZb8HHTK
eXy9CIeNiJCz8ZtTm/8zDZphnesOa5odR9es4JZnFC1aftZ37TLVQxnZx/Ao0Rdu
FX+7G3HxSx2T88KI9v7MzJ7CBSxfiRa7Vs7FR4hyduxoOWhO7C3ePNoFeiNIXtX+
1FLf+WLQbhHgq/elLT5+PbNQR6kZqAY6OdNC5FzJNW5PRetnWspfLEER3wrtnqnQ
MT7sJaF0Sf79xL2yROOd1cFRYCPYcmsxbJokHwe3+J0mW2QUbcZlfF+/oeROWF42
pW7NWRMXsPamRGZoaZ6uTtuaA6LipmpDHuQrWCAndEmNCtiHZSaC8D7pdXlLPnhp
48oK3zEkRQp2oFBb28WO2Bfi6oJ6ZgiikVRbQu+1JAsPFpaYlmjwH+dUQrYdHB3a
mL7uy2f0lAcMAFOlQf1moZX0hSKNcSGwozPDNmLpQKzMnnl1lauaKM42ZB7/Kw6G
Xr1dYlwsMx341jH1+37y6ZbD/onj5cXnguupprnHw07bauQzadkU709kdu5CXN/F
aeUNLHTJBVsExdqhdYPgEnpF3YHzHRzj+mQTZIeYhmtN6YCDjNPPuj6ecwr/r75I
wNsAFpcHFXVh1I+blQbNF/VgskCvLWKHtIhNduV0ZrzFn5ulKXLmsKyIFUG2UrvR
SzCHTsyjqF2AXuKZcmS88kK4XkRkCl5lrIWs8Zc7UDb/BQ8US1KR9O90v0Pf2X7H
GqHPt7uPGetj6qBmRyZTUUc3l7j7cXShy0qTdUgCqE0810epv6dZ2Xje9rQu5i6O
whArakvVCUv8B1RYhgzv4ty6jH+YDDGJTQozFivV0u1kaMWJByIYfrmRKIQwiK4/
mmAuglbNam68Y/KMUrAUgW0T4+QArIoBASfAURNrOshm5Krbs1pbIx8BQzqa4P8L
jP3cvNrvrRU1LGcG+9sXUX5D4V52v5NLJ1fk7KUE/mcgplMzwmodDrge9fldSgJ1
t3EnDL8KSyYjkhjc/+XeSKlcv176wf1G3Vpw2imS881hDYeBWz+7a1kDmIgr4pJO
SCHBzuqbauabLj8d5Ff+gGCc+zFu+590RZToR25sH3iewij9bpu3qzHqgrtj7IKI
uQePw2zRrEeihSlDu8yZickPeTpqtPTaL/cpCt6zUiRGMJBQD9I0FLxfJYKY2Mj9
LU/LjtfcsGzsVM4jUp4osRDWSJjUJw9nzQagZdS4EBEf8a4cUqOy6z/DLCcxN7fj
hXrp6jsSCs/0qy1ocPKwL7U2YHSSmdx//ulN7FMAdJy8POgcT8TdSCUMpyd34htI
uEylI2qOJoYE7PFSnFsEa7fMC+8xDBt/YoAXuq7hUMNMxwIO4xKtOPF0HD4mxi7E
6Eg5+iCQ8qxt1dhUKlZXSWDB5PjncXRJNICgajxC2mPgC4GVBe3DE7nI+vlzVki/
mc21Yea1+jU4u6zVclN32+1XPiluUPja4tS+e2btEt1FRBLEJpmVBojZs1aAcDLQ
rLu5G/xQ96KZjc+OI3CYf8nUhRat5XiyVIT+G/2hz8u/UvxbnadyKrZLUoKZLQ9i
ULPkycxWABUglDmXr9RLBEp6zLdonSE6PE7omk7POSN4nz4a9adMJuwUAZEFxUfD
yxX6s8EW0Usf7Ej3VMCHBp7m9+SIYMJikgFbI09A04fiXLeiYJsmVdvyADUw8hTy
R5znNlIKMVCfuwp2nIQqPMyxKyVswjjue9JQkvg/mj0XZYEwof+VevXDGkKIKtpv
YneK3mMkaPPnNFWpqSH/QOdId2/fM1B2GqbEilmLoEEriw+tIRlol7xpDOiMVoEi
4RQDMqoYkmIMqjHVaIBzjx55ICuH57+7xbz8zf6sHhPVD3Bde2wjXBNxHKlOVbKc
UTVb97u3UDxF9yUdjg3zBZ+biO1HTB5bCf4/bAQweuJiITN/Yym+dbsetMt22CUx
uGnd2G/BsRNfcpfumSQ55VuATKxduxiTj1kjbpNuWIKVrc44iMVVvQB8vHWhMAvb
/XLhKDnv9Ge4ZWsnDltvnGZ31yUfdPPEZKH8qC4GdHnhOfpgXTP7gEdXuDD4wJr/
/mJOyIgifGzN2LukbhKNQXqnvlRg0wOO5kJAp6u7/zFHOqpbrXcok9hu+i768CDh
qDVu4/ntSqMfgAnt1/ji3I3jaydLIbHLN0GidbqOf4Fv096bUXNnwyCEq+8Xnk51
7UOWQHQSArrc6F0B/MlnkhGodJagt6ryhro7SRgU98sb8nM8IfAyOb2sDtyFT9YS
aHIQT/GWEWEaTsHk3Kiecza3BGfh0zolwMkuTxJ+2rn1Vd8LcT1qnmU+J/0w4OUw
XGf5+dk5WlddT6qLklwMZWAJnIuWGiblJ8ceYGmUPEq8T2Z2+gZmwXZ5Fn3V5D4K
dFVYSoWvQ6RdXXKWs4QXhIdOTpm+i+IK5z64W9TlSLJnazHj5SpAMTKrDH1B3OiN
AVf8kWQXY0YwO4bmQ0VdTfkatHHt90L4Z60ByxrcqhzkrTYPNwfjpLmYVT0iMPp5
d+py2Ot2y3S9H9XAL+KT6LeqC6uH8WODAQSEhh+HCsc+fBLI3m7Px1AhVU79ZZ9g
Lt3lYKM9hM8vSc4rbS5kMYPhgYXuiJG0GARi478t2SIKB01ucuBpfdIkfSVJ0k4S
72Y+XiV5MznguNMfN2CvrXpvimbm3k+DvZVsQqg8YObUV7Ao+wCyzeVBZaC1uITL
lqrCqFqLyR9rM7gpR4NvgNvF+FO/Toiix4/7w/6mk6jdWlvvYq62bjsos64t34SK
wYOzJId3nRXWH8ZkyQMSqgpgYGcwO20qJ+Aim9QN+c5Yn9gza50Wn5ajmBc3M5Y0
3ZE57cxKF16PXmfIf4nawUOhtN0frd/7XEUkxRlz2F4sW1XFRSVlZc8xySxoPiJ4
Beo3WwDP9MgRCJItgA+zHxnP2T+3MoDk+mFXsS7etkxAdXW0vTSAIQ5SkJ1euIsC
lkde/qQMLKuFxTFWNMcaNueIxT8yi3DpxP7xuWU+gWbyk7owYS+00oGsd+x96PGX
3IMqVlCvTHTbzJqLWAaPE17sEBugM87n1aXZ5663nUyJUj9wMQ60fQeyz8mhzZAA
bSNhDR7l+IFMqUtF2CUp8KbyEiCCUgmiNWaNqNOvkBAURm3o8lH9am3xcO3zVK1v
BjHTerrzPOE8yzzw4FfGEXcYMSXEgiaJUUpZvogfLE+Db9EXWhbdQqU8JhDroMfh
yJXEy21aEP/Tuc384yThy5vBrdDGANOOwIJtsqg7hNmpKSeV3UhOyHwnDck+2PYG
7zve/knvfm051QwEIAv2QmnTgoQkSQWs/+BrpLC7PH9UyZK6iPvfZDKs5mtD2TFN
gSk3NVHsFn4wtp0rkXQCuKn8k5tw4F7YeF7kaRyzT+vVAsFRNLM9hEpkv97iOwl/
9ygqaB7uIltQme56ICD9gYFaX5fmTxLOdBWJAvfUff8tBZ761Wa4UGawsWpq0vlL
RaDugM3hSgwNp4sOL3e9nE9BdJ8cRK4l5xiphbjjOfA3+2MeQ3AaxQm7lfnXvZT6
Ygb/tnsRe2q/8Nc/zioajQrWZyR0gpifRlsEI7i4+6suj6yYsaILpPuRQhL2s9IW
9bNmoRGUkyWfwnpodFEBqWbcEUcvXUCUMm3jo8Qe1hTbcssUlwsSn3B7J48HfL+0
pHngStmkWK4lnve5FRzsBx/M7bkGkmQ9cRnIviHSCyOornlVGaI87pFM1Pl5er3x
UZ0LYzBA6xuZkZHyWI2ijeKoBuTQBJGQVDu8pM2ykVvYoUcO2Xw0dMsrUE3JP9Zx
/uHOGYIGmdTET20Do7W9ZWlHLKV9Cdx6piLJwKisRJfSZ0PrEAmtT7Cv7udhed3i
1qxanuH/gscgSnuo4OAnkS20ACXT9cYJ4NWjr3ORcx3d9pwgZRs0/d3ADwpb717e
GCAjHOtUhfRXF8hlRwDgji/BQktREPDiAcg9yosr/3FsrPWhEKPicIFykoeWL7Yi
ILcy+vt51CgjaUpCCZkw3xxegpkeFGGSDMyEL9WDf6kkHhERKNj0tHEE0qZ5fBtU
M9jr9H2tmuWBHDiPdkKZOA1AXWSSs9YMca4VaHxDjiOTIKuOTuwzuxN8tg9BNs2C
hjoM3F6DPT8/fdBZpkLHouzDCXSYm4d3jlGl31bxZWVfvu2HJ2XM0tu2iWbEh7uW
2jbUgKNw0sc6eymuyBY2o7PVicXrij6AdnhLL1ya/bVMyIsOu2djR1Emuc39rprn
pnoYesOYcxKtzAoiinDUtAUQxyekDUSu9Of05AHuiVqytUygHQhBuwwO080K6blW
O65JmeOEniG4j2+YiPNrPjqcoaY+48wo8IAbDJEAp9pfILKLMNScAEZzklQCAVht
9bNt2ck/9uEXC8xkgtjC6eNAjzk7ex3sb0wbX2Vbdy4bFa/6L1xP0pu/EGIhqYtA
1aJA65JLka6S66B/s6PklhtT3WYzn3mPfR3XDlkHhlRGwBLajGX+Jyh6xYA5rp5p
pYnECVMgbigynxrOuVnGG1LyHvM5ilatMQkqM9rZuGHzwknYxa3tSC72miHvawhC
iqlPRc9DMJ2uvDXuM14ZC33pQYX/dfhLHeIgVBi3zqF/UHaWzPCMjXb4Z07+x2O5
0YQk86+1BsApLxLZfKQOU39cjThCQ2qVnB8sObCK53yAsZK8cM9sbQ9mBFzvENUW
CC5Pbgwo2DPklrhrfDWwSkcJK1/4E9Td0uvsc1jgcXDa7UCqhuIlRDwNtxI5AYVa
TJcm4UBQzkD68uXfGsngtjTQSlCXJdlrz/tc87bHURvqdbG/ar4f4UlQTUxlDAoU
HqTJwv5eLF79eIH8NLVli8hm+WKDoBGAt7sLUzJ7wa3wqzGe90UEjYdk8u6kZke0
OXkFQxiy1ZgW79ku5htvrI0A21Tz3re8SChXVyVoTpim3SNnL8PYTd/DAl63vTxq
C4dDNnFuYUg7TIVbYykiyZrPiS9lCLSUtmKJAilPAUQwM7eqJOQzmvQ3g7RAztYf
ncuIe909EoPC7MBGLuWMK3K9tvAjnbOvEex+qwmK6BykOXaainsPEuzb1gDNISWK
RcrbGTOVZeS5iArFvZaDLmHYYNxDirePqEFhE4W8MyMUqNSQBZkTEEOcrp8btC/8
1x8sxnDFlENdDMgzK3d4AroWl9EC8YjszeREuIkB8oFjk+d+PIYYTgGUE8GObYRP
oQOxHgPqXP3HXNPYbMRXiukbWWVNhwOLcbq8ooRke3/lS7469hmOhEME36SPPx7t
dDQnS9q+ebGyOcVMVDHsaFdEGN7z6yjsNZYKHV1kozMLgPZDn/QLZKj+CugnaGAL
pIIBu256iU7JmZCLSS+ziHD0VYTZ6EIXXSd/Qgf4R98qsskZdiFkDvy+1PVviBal
eSFcgDDRcd/tD/k0kaPM/bhk8tDDl9ziRuBbO2s9CbiXVSBNAEDg3ckQebeOE3hX
zd/1mIwHp/5aCjWKmitiT5Kflz5/gehMlpYNboY/OTfJxCnx67uK/9N7vKy4UXYR
if18NlWiuCl1voE1Ok7qfWWrpj73LKMSfrfbfTyiPTVZQ4tzy6qm/YFGJiMlo5BP
Qw1jH/Z9djgzp12c2ynI4MlsQtqhJDYr1ydB5FqbaRWnNCh+T73THhAyMmlBdm6I
sgvf1jIYDigortgACa0aMpiI51bl6KHw4/7WWMEf4xgGn/fktdUHHPj3uiKlXEb4
Tkz15FkJCJH7LVeTE80esn01zihV3IbxgDUrZdUoT9gL6ddsIea0SWmxqjUDR1aX
0KOVoX3tbs5UVP5+RgAMsDUWYj5hh47uDj1V1lX56uF0hq6CKRyeNEQA5erifipL
i83F1HvynAsVKKT9xVGRmX9lH2quj1fGZap42pyvFpe4fASPt9YLoT4KtegVNwEH
B6gw3WG9e6brypANIP/W8ZSLj7MjliwMMwVBOFtRnRJ13k/MzS/b35UWjkB1W59k
nt/QQukZkA6T2nS0jPl+01hCNvISrzGDuXne3IzXruslO8GbDQzojCQMu87LHC9s
KAG8Y54H5vaOGA9Hw/ueLx/meXOr0AQ4GGWXaxQuikqvaTbshe6WHkGWc6LEaMGP
WLfsG2t3vwywFWo9xq5DvOtJC5fSLah8tS8LbmLZSPF5BEzsw7sbbfbZUpe8G3vl
StYVztjUI7lO2SG7C0DFGRBMy6kUtA+eiTAPOdxuKrWr+TtcheiyFFoux63IL5sY
g2cV3I8Wd8IEFaIFnKVutxWg8f2z24+MFDioF8PAI7kAK6Y/4zjblpoJs5b5WQ8C
69+4+ZpHgaoiLp+JqImH3Rm/YK0EA4bhoi7FqGjDvkxcXkS+GS25c5E6y/qhEofu
dHTeqm2uPb27DRMWIsRftKbo6WBYLkiZDitvQi3NPMJiOQwr+VJ+OHSvEggBg6fL
shlGvDMbU/q9sObpNFDOMC4fLzSAcCMxY05NEV5GlJ6Rn+HATT2ja7N78AxpZCrw
QARU+/YAh9/WTLD3cvqG3cNeS+mfBYzHDDU/6iuJFApzrbw7xUXxW5T5lUdwhWIg
z7sJhS5cDeuVuUXuTc0Xc7IHKwUlqdWpk6TSRx+cVAzvsaAMWTDa/xklNzfJl9Py
62Okzta151pIkREQ2UgZV7YcNE43mRSFXbsAEI7RdmWmikQrNKnolwAbgpDHoImW
ychatGN1ZTroDXQg/HFjPsv3s2/m//Ro9Q4NZ5mgvLNU+zgAGNvFbiFpkjm5vTGO
MtKoINFjT2nueclx6mAvPFglUUMpiUb1f4/VbTXDdhCCJPoYpPpk9uP5CFiJdorx
6J69G1BBiQezVh67NPSbzULRAX03RnCzRRV9L1u/QhogW874uvlJVcAOQX4y8Mvv
YEr8a4Z3XK2AU8sNeytVG0+FHP4qV6uUqT3JQwbgcoEyS3pJ9HtZp4q6pzGbneX9
tmjRg6vkFSgLeNYzD9sopyN5zI3JZkUc9uDEAa05+Oi71cFGcDBFlxN7QuGMd2Dm
NT6yYGTr2dt2kFM6U48f4OyNtv5N/BSQ+3eZlrVKp5Z4pPrPiMfLZh8zgjiS3EA1
T9cLqkcx3e2t3h9Le4JogrKt8YCBqQW6RP+OC3uZYCvAQqUn3DNebudTbE6uysZW
ZiAQhXQmyJLa+Mw6AqExuPQ6AOnq5QVgjqKZc2qUKKLQgngK8x+zotfvgujNpzbi
6nIwHsnVYi0Bhyu9Yvk3fj5PL01KYl0HzzeVYD3PciVHq9AXKPfL2yxrLbGPPkIX
gWzSDe8N+BNPn+bOsK1mb3bAjydhVPmb7E2+BsIqSPlJYqyi/e+czWrD27RJswFf
psHsobmOvCtw/DXdjxmfXlmBCKzkRl35j2wdysBTKWMW5Hg+Dk3/KuTBdS+pkNXG
qYrd54xJjGJok3s4lJjmRNsrZdrTftmh5sXuYf7KL93tEJLQxMnsSVWkBOPAZ0PN
LF/i+hsgQm5V9DyoUNS3vfDsgBdIubBchIi/XkXrAncuW+iiT/DJWSHsNcXGn/qp
/ybVYxMZxseMwOomVVQHjGxrtpfePvfbVdvplC8KUQNpynvBQoCSKXYiaoV2nhg3
/U0Dfuo9lYTQTdhy4uUKfO9DaWLLRr+LfMWrLzWunwS1EiV+OnQAze/+uXsaFVeh
jHQtdmKjHOR9bGGdlo3afrzGZMthpr+OwNRPWBaxDPoktEuNdkyw5FmHcGE5iYoz
VZ+5svXsBRywinW6uzTexWVtrVnu8ibWPaYuPLfwE4eFm/L9OVslFXVD7B7ZEoTy
zB6qr/hqv+ogyBWXBEuLhaZcyIsXFdzpKNNn4S/3rM/Jc3MzIbsrfDula9awdg1K
eNFAY2XXdW04wSAeTJh09YrGtJ+YlVqucuPYXt0rJRG85CU8VGCtR0/K3EJlX5eq
mVgGZbPmYixM3snpk8OGzPgMGFgWNePjsCU/Gtvx+4fQDbfhWayw5V4xkNGzFeKi
GMEElAPP5IVTCaUVk50vZX0Ze/jRI/jcK4AGMqu4w/mRYENnp6Lh9U07QUMYVK44
XhYOHOj2jS4soCHZhwfBOLOJV9zSUb21GlC5jeo6GnMQWIg4lzgvcNEyNPa+0D/3
jKLy22J7zZLc38ElMcT6tavTr62XJQYTdpJ9q7phg5qdyP8VKT33nTQND3BWZi7o
KqIiR2+I2wJmDzLPYp26gRnfampXoXAIBSFduHjhMU8rt1pcEShrRG+co3iRSy0J
BaMmtOefG23Pj7KU0REmMV1xJUSxDuFXrhtJcpi3Oh2HtIK5QVGNVkbSda6dGYKW
SCK19oLXbcW8C1zhow73RKz7xRn6SoaFlcMGpPKBAzmWgbMLV94mQAi1R7lVROuQ
OkYfsg0dRicXCvQNCKUZ5CJHXtL+tCGJ6zNP2xlazzYbbr7IoYh0M8ldEKom9jRi
tif4TKeSah3Y0ave9Vv3YPdAoVhbulGGCPsqU4kfkDBaiYj40LcoGSMB9yuxssPg
X5Y3D9X4Gvrlq4U4sV1yEv+zvaAPVceldEMxKeQN7Y4+7zciNlrW5z0G6aRM7XZL
UqVHJoPqhkLSSPqOXjhr4I3m6PYRPKce68fy1IAee9lmxH0FVxb9mEi8zByNm8yD
Mw/WsINDJAfCbrkXdQyJeoIhK7dTYiethsMDyg/Mjc+e4BIV68Xp6QhEi+ki0wVE
A+o4OJrEf2ScEe4SFRTlIp1AMBu6rshCdbBqgTX8dZ/gnjlKCYpt1+1WLr38EzIt
CsKn7juj04FTUHLjYNwTAW9L7u3C+p9frE0Zyzmy+fViqHNCXtusqdW5VhDi/owy
ulMMXWRTe64uQHfviWUQPcsWPVVl9c18EQZfdG/93Imh4gA6niktfc8q3RqGCpeN
0auPph/J1EBa83hE/P/LbFvaRFeD9Yi5UwCNOYJvjW1lL2VXlvpYBLDg8hmT6JrP
Hjj3eLPfzAEVmOTAiM8HdkEYOojRzLpnGSIM6S4OSXhJmzwnVaj/cQMHayLfpWa9
deg4eHAfFBBmhZrVHJs+7/CMJXZsVny7AouRkQqjWtxlIdfSq2q+GnpNvLk8TE7A
xDNPDK2l5ztN5DbHywcoiZ0+Lg9SIsLeBZ5eZJ++AESLvav7t4UB2NdN0mbUVuNt
IN+sslRLQjQtCpQQgVRgOSxUmbpZR9Iwh8Zah4qHQrppXCLysANYRBhtB1qhqPOT
zRNEddvFyt83vT4GLhzBqtx5gNh8m5T2yDen0O6aEWEsTWyhks7AY3sQL0UZcJL0
cdsdYOTxdDiXbZx8G6dW3FgTI1gKiDnrSOlmBwKfrHB6mOC5Odzokm4a6sATu5qn
9gIYBp64gN6KmngJqrY+LpIpHSS3PuFt109CTpQ5D1Nb2vQEY3IiMiaDCOP9FBJk
5W7ZJvNCwFi46/DafTYTSidtO5ynupxpE7kWky1Bw9r3zVOQUcMCqTyAtKJ/sjiS
VcnQsQ+buwKwpPEOU5stw+PLBSzN3yPeQYSbM20mrp2kSWxnthNiX4yvgMygKioI
PM/kRInaubT0yc+TaG8JxldaMo+Z9VKQH4anwxfW3f0XSkj6w6VLNal2ggQ0laHb
8RNqRTnIwWH8//kcRifvAyHBfINjR+jADw0q2/jzooFR5i+eyq7BBanSvt3PJg1z
Ns8h/RI+wD8I8yTTULcnM0NTligjQDYsZ2svkP9toVaJS0kYijACXQjDTt5EfRnR
fx5BEqbcC2BhimYe65IEW3XvUVgw9wFIY2mV46HX5JPlfvdWzNQZZHBWZ1VjeVvv
/iOBqEScyC2NQ3MHyaRtk3w55KTPKuPPJjaVCi+LsgLd8+nKw+4YqSLgu1V/iBq6
P+gEmaPcHXzHjUnjGWvXewudJHkk4R/G60eNCN/+pXzg0AlM7NtGZRQgb343YAQJ
ymJjPCNTUPIFe9hvspWvLgqIQU7bxH0HkQhtSSqIXfrEb+LtwX1YpoGTIb2bKBN4
Ht8zMaytB4/uirRC9uHyPEcBe6FrcRZLOiRNvxriFL2mGqklZtl5UiW+oekxhObi
UzJvYvVSSve8cMWbinzkUkdkPH1dlXyYWfg9kDdh3BtyduMW+iewXn6gwZ+sjdzC
3XA9H4vTw7gJB9qlGbf6D5XymPszBuU0M+BAoAi6AO8cCEILTzTZJFtUpqx+W5IV
m04jWl0vTvdJT5TAxBi7bLfOjzNo3mXbHF/aNP2HRa2loqGrb982RXbdOGNCn7JW
K9X1ff4U6sL2ApGHpFVUsA+euh2aKHspnhzTisKNDpGXiq/HMK9WDqiz09dt9wuk
X3l1IXa8/Y++B0KtZ0zhdCmVwyAcPIhEB3HeuS6r97Pd+/9ZDmaYoEvglOT1Ep/W
YwtrAMeXNrW7tmRgqH3Ge2Yo6J3nO4kQysmgXH4xpcfRrvBEhnab4M9Oz/vLn6e5
KHPEJHfHmG8xZSqPMaxKxBwD9UU5U6+o9s6s6TgR4XM7xjykz276ZKWO4Mvq3fuP
2rOzBToADtfNbqD6YwXLF9XnXQR096LCApt5DB40vCpwczp3Mb1OxxelvRtvCvuL
tXWcPIW2ZsSiI4jU8kYKM49f0Bx4XY+oZFV2vBr2OPSNYLRLCP79DYYLq0+MCqPa
fjf+mQ/MvRk7PmBNAPY24bCpbmna2FrLN9W6qGtIECSv1q5uz3iTvUHU4lv1/LdR
8sC+aY88+VMrtoPutUnZ8zAiB/Llllh6ybowu3tcYqlBnI0iIw99RenhFhOkT6Lc
XC3WUiyxUk04rXk+5ef4r601QOJ0a048ZUatmRbJUgXMRiEi7sYFnvzycc8T7k1o
4ptiCdtaCi8rqyeLYvKhov2thVlmuem/buFYEDu9nydtsZZ9RTSZwaHM/9BXuvK2
V8t37qdh1abS+1YhhZv4FNPMS03WAnq+QDXRz9JfsZliqynN3+WnXXFjL46rEeRQ
LnfHe5PaBjGYBkFxtH4KXnbbo5AiA9Bb0bsFZIfQZGOD0isxmcAzX9MdV/86rC1c
VvV50QPgKMPFO+rtQO8KspP/RYyhe/qImjmXXaW3uA8U13ygNknVORT+Hl+bON25
cdxgAOPsz+wzAftB3NwQs4kSjnvc+Xfk6qVbQJwXROcGfb4LWB9MSMJotQjbkMXg
JKBHYG3pVQ8PIRxFTDA1+cACMk9wGgE/9OP0GFEWozFu59BAgsNfczpvwETskGPJ
3IKR7fdY4Fb07aFIetGdx0Y5YrxmkOutfKMgRgGlJ6y7xPl2ipvtwcZS7w7XixeK
3IzYz1J5r3FIVdmPMhWJLGpBRug+4I/d0PO2LYNqdbyfcPXoye8oDEo+6vv1fuUD
PPibWRBhwHD9629kmDPTxmpecWC9Z0u+0Q1br1Swf1Ds6DCDbYi3CnPhLiAx+pQM
z9l74NCVttPAoAeu6HJSNvABb4dME6zVO8iz+cAenXLScirLsYh0kWKoo/IiZYTI
nMApOFhi3Ug5qUZMHWfaGH8FDS9TZiJa7ebS3Q8bdV1c2EQYRWxeaIlhrDB2kcVy
EZ8xxULYXz+GDtKp5yVC0yVYOjXHbaf8N+C2gLjHjpueypPmClq30DvTChK4ZAvX
ZCXnChDF1ZVOnyTCwUgx0/ACbFHs2YstToIrqCdjjPkXGXQzptjlJ0kcApfjzWHA
KVdLEG2U86RbT8RTCGaSDB139aADgrWgFa2rKnf+Y34cFCxxvK11YTGmcI9NabtZ
LdEEJdmE4gEMqMlKeE6bkkhYgiLbOV1QVkoigSJVJadealFErm8hoDneF8XLq4jk
vcFXhAdAOIjk5MOQS0bog5eKVMNq+5fqmVW8s5FuZo+FCFVu/axZDIFER+0DbbZu
PzSI+udXJV/+J1ToIqJl5IEORRS7dxg5jg9YUalL4JebB45tRlUIHdSmFwoU9/qd
sMupsi6B+qDVN1mGATQiWIm0ew/LOkovusuedCQVlgm6EAqsfB3y5PIb8zMWX/Sg
aC0GwTg4dBymo2lb9L9jjwB7Y08EkHnrg41dnrcUnoygAGUKqVviIeXpZF3DOm72
V9HKjsOMgFi1qZOpMtkiXBWZU0xx443Yhl6ky0PGgJ5d5V96COjnuJIBv962PXp8
2WhckltA5eRBQc5OOXBYBCTKaIj6TG8esfBeYMlHd4FhBDkI9/2cBwh/Fw8QjcT2
GIkGpd7MEF/7MIQTIhwxT1OfRGukxCEuPiCpVIAYWLl25ApDYBFIe6/enaKGSkKJ
3LZEC5EeKD8sFnntoggYpaz/P+/uu1xpjTjdvf8ajA85pRE5unDOwwWICA1lBgJ/
k7dTCOCPw+Oxd/Kvs07ccDfVqFzLFGvuhanknHbkky8UO9p/FmPr4rI0JlBunPDc
tx2X6PxKGo9/IXwFJ9DabgjRYhVYwBpvYKZYLHrSf3ZW25JajHXTV2pJ9+Yz46Wm
E0TVU52mJmTiZ+68zvLjxMyEk/V0mP77UOfmQRf/YcBTbiIgk2hgPNVH710zlvKm
k90CHf+9JI0igJ/d5RIvU3ysdQsFDSbMJuUsPmUw06kS1OIDuWhgMd9rTdM2ZmxX
fUJDCfPlI7qucdBv5/rLwbv1FUWL7TtQ9Y/5LeDbMQdtv7fxB4sM3eFxZUaz45WW
lyWT3xYbDCSjTvkHX7UaOaqCZG4tW0TDZXY6KzmaQMKoJJ6uOkLmMNutCsW2NMIt
WDGj3pM4Is2G7ZoX++Pgq9sP7G5IPuPZQ+gPNAelugQDLYr2NxFkANGmJogATrQ8
rESc081GXe+vKXvCLKW4jb12GtvX9hqPQExZlpIfC7RcsBhClzBIZJNR132qVETu
XGo6iS/AWTzfJIZ0yEOQ8Zz9oUnIx8fnUjxb9um7t/KplmpXTF/zfdviM79TnScs
zm+PXxOWgHidEeAU+SKWfEp+cGIt2K6wPLD8Dyjos1uccSCvkwtTO5uMpEywUU3P
GsvdxGrmxWIDV53hlm27+yMO+1vAyMZW13E0QxKWDdXoj0WAg2+Eyt4n64Bstt2d
xLqRLSJ3oSgXU9D8YCT/Jk2Qce7yqM3MM8yTsRm0DUBPejZLRsDK6BwHbFgMMMTE
Taq4lefbzr8YckJUhGXhAmHOKBo3F7B8fVkLhp8dB2hM07FdeEFVnhpnnsODFys8
BSMg/76atw9LyXffGUhLqGU4UsoljG4myVI81SYEIP8ZC4Ge5lMmld3mtbqy610j
F0uQD4zF3IIxpqHrtpsrFloCTZhNoVMf2Ict5godEmbg9BVIDe2q7TBp23a7niJs
CRFtsPSaI8sShvZLV6OwRQI930qj6Cy8Uin7lBhFni6Ha9xxqfPvgvlhcD5FECMx
/+HbJINvUYxTlDmLvW2EzoH0Ys6igYkeNMc9I6KnzZlk/gLOGprrpHZWQx8EWtrn
pAVO1zbu0VYW6CPBeXiMnKPOR2iGxK16OmxzWLpdFZ/El/UfvSdMFywdq0EpIaKB
x3+SDF88LEaX+iBCyRY4wyO5GjgmCZLiF4zlc3xNDNJS5O2jB2k6WiHbSwtydnTY
eAdjAoY4/jkKQUKXbk8JUbNy4yhACSBiVs4Jugo2H0K958wl5Bb7Mm9YkRubZ7/C
uLvU18A1255dC69zYPhD62Q8l7eOnE7J567krdwRU/8mWAUi94EVcJw4lPL6o1D/
UpVeRcpSRpIOkUyiaOxIGI88RiOd3bKn9cMsxWNqft7rMn4DUDg9dpg0oGGoMqRn
zkgf4X86IsnGOlwsEwUyxt+/26a+OZKpQXfG6hMoaKuCAHN9cImIYAAWIvp9m1If
Ry1Yaq8OkK2egqlAOTZfpZhGRfkQw6EIVB/EzZaCPAYKCTrwxO6JW/b3OS8tGokc
Q92Nr2mq2PTRNTjUOAike56fjy4vB2KfArSerYtSjp3Apjm6Y3bpeBsKFE0ESTrm
7pN5O5JChFSPN7DZTBCldQE7X5CLqqAKV3OVYdhCC782Ls2gF0/kjwOgw/VAvGdo
nf7qNX/d9pkS5g6X2jXcw1MjPO6iQkl5PE0rQVR/q/SDo/WZMy49jIWOAjRgQ75b
I7VhRwvNQra7ntndjbKZfDsaiW+W34CuulAjaej7zFpvH31V+pJL2wERtjSUgNYV
L2sJGGbh9/LbGreqSOxMvp4gCimg/qm8uv3uulvXUXsmdZHSG6czqEsUcxpVtql3
36ew3P5YbmD4VaGfvsobg23QMZYnBURZhhaL2FeFKOXHhOt1qiFQa9xFoR1iX7wF
gZXXAVjljCkkFq/or2X/QBL/Kl27vpbVHmuBOaL+NU+jv5IBSgf6bSVFabSXNrK+
Toq7+mYGfbMtwu0n6Cu6kv+2k2Km3WbnEfYUYpWiYU54z+CYaUfjGe1p7yC7wG2X
xV24BZb77+tWw/2BecsedI9FCvkYyYwQXeUUtT8yKZ8VIeikkKNuUwpAxO/WbyLR
oQSRCqHqhrJAInPHOWFwO1pmSlipnGOkvn+PlvIsAEBvpiMstWOYmmY9MAK/VN4v
U3FcEaRX6ed99GnxjzVeu4Srzo3Ozb8XDczcE/4omenjD1YyQWbgar9WIMa2WZ5H
kuTnxqoD/kcnSbRrKIUkY5nnISJmDbD3uvCv1OHLojo4D7NvyJXFZZynv8PHDcxF
dCaDEVw45qjMok5gfxAIALctObpnRvCH7VKNvHNQiAQaRMwDxA/TCPPVcuYAEHF2
Hq/B/3PTGITr8Vg8ejULUJl0ZKEYkdZkkbDJ07Z3ozNwesEz3MkF4tUhAuPAkesP
JRtZY9Ac0bgcT5hiPtW0gh+oy2NXyKL4IwnSDbahCy/jqbRv8yrxRH6jmIF7wuhk
5tOh6INHbVWVUa7Sk7ZjkomaTY8RDFYaBqtee/tCUOOOLopAoYWlQ0vyHuaHypUC
KXANpkvGUoHbM4BR0F8Cp/KH1R0GwvLxuTo36Jy4SdAiTv6+kWJp/PIIZbV4EtBm
WTG4WX9yzVvUNTlUoOwRGuWAOnOOA2+67n5TRsS0ivEqqe9V8MSgONPcjtuY9rxV
qkSdzKyqCeHICXMlf7y6wEbSp5T8yj3mIxqEfzY1MPWqurOt1x+wEjyDDc1+ACfD
iJaszR0I3erKxjV5auWLBcLfEpd0bwGGeQt09rwpiryRiG9+9m0KOcGws9ikUwfS
XhYeG1ggMy5uaAzKvn7x6gHQl55ly91NaaKaR8QJaiO8OGy3US82kwe3j3Hyf08C
DYwPdacVYYmRLw/9+39kA6oi2/Ux7IRrDBH9Z/1u5DrKuyC8bSXoKfh+vcYTf5iP
m2jP278qSJBZYK3palmQ1cDwRmvYx7dEhcl1iUFziAqLMDmyxy7YVgZ/W3AP5LsX
jEa5i8InEUElwY5/6ICUnKzDfvp+afPpu1DgXwM+G1z+bN+/PP4KEc3EEj2UUz3h
Ak6iv3Pa6WLo8DJZXerkkRBpCs9PmmJTOlHIV+FO9OsUSOMmAUpRhrMgPMykVKVD
w+I9zHnefIq/eNhXocEP+qnmm0YzqVF12qNhhqNIIl9YsHJL62w9MAD+xQ2JpLcp
iItTBq7pSxFGsOBxgYiJTmDU3IjEG4CpdwOUSqaieYbY1v1Cy7gjLMO/QsXlox/l
/Epm2XgW+8UFB+sh+AkhNPoBV1JdRcoxrPlk2DbritRHViaYhztGOtm+gSKhoty/
UL5m06C0WvPx98KK4XxLbqK6NMj3jL3XltYslLi+rF8sOzu1yAy6oOyVOtGn/SZ0
q2CUBjU/9ErkK6cVi5fONwE30Pno+95r03m9ufEjLN8UL4deZB6TjJlCXJvLzmRc
i6ofx2JHowi6qCoNgKHu/Jsmca1IXnlfBEtJ++upvoMifrnHIHeJuKcGTWRbTzCD
P9v6XfP2tgGAVzfYT2JiQTW9FN3IkFjeYzNdGSKmpW4y2v/o8IkXu0cJ+KVQYy6l
UaAdzVEG3UqMlqVodFHZkEB/Nl09iZGY0NcBpem+FCmhlyzIFmvjkj6AZ7wuL56N
EvvR0Dui/vrAxxAU4BjqUpibjWj4J4q7HJIx8yXzcdAT9300hTuKUJ3qg3uVGFQL
j8Pm3ywWiEMZbE+DXZ5hz9JPnkA9iMK2vGwc9FEEB2H3DIYL+SVdqd/92LuS9cW5
EwdHzUVsH0UjWKxaGpOZOoPtug4eeMsgQ3EdbYBHyg8+xK44Hsm0VYrvKyEvhys1
X1yNVhRM+RlyCAGwL9tVGUNB0naHBYnG6OEq3W7Dq4s8FGlP6A0REPtQ6HofSIRE
SUHzI0LwyDQffmi3nY01yQcg0+SlBsA9seIrIsnfOfd21zq1UajpRAS9oRfXBB5o
Dr3HoRJSjKx9VQng2TxQ8FwphbxULOVNX5DtV5CdMw/+6gCLw5C5p6JSjrS+hOUf
KO5U35WLxOznxiow4MUe9aUpyPVaWR06umGg7v+D8Yh8D+tc+nIP6i/G/7P2pZ5a
T/C39LAA1GnUwpBmjbTnGvX0EU1d9w+aXCEMg7fn4JcwU75Gcjz8SNQ28W6ANQwh
kFZQ6rgD8uXB/9I+tZ5CzgNBxlHI0/+XKVdNThGGItaAdbe4Xq5+Ig1ANEFWH8jM
7D6P31puR19J5/0hlPBF3mo6eoohAgMkC32aelDp2b1qrVzYFWpmy/Imc+/UY9Df
xbYmNJCwwELf69vWwhMaMvdZQEmnCqxTecPI0ljdRh1Ak3EgxP0O9A0F/7i+kyqq
RUyqXxR6EpevBbxZJNWJxPw9FMyOpDes9uh3iLi91ZG9Pj+chDHWlGVoQ6SpyRcR
OedgFY5WxNonFUAl/WY2qgT5Azk+G/PmRYq7d5dPLRs1mpAbz04hbXMWMvCDT3zk
ohfqXhXD55BvjegOjynVFc7mSKxVwbfL1tLvMX9sHEG/eB6l8ekbzP/9/he/nKvv
s8T1Kq0jnRpVNgX8flZPN2Lq/6QY/uGwGJGbTL8EccN6tCKjAkvbjkLH5kY4vUhq
qUrtecoMjHTqXm/rasp1Gko4ybEi3Zn/WZnXiocEzYv6maZD/0jmEALZ6FGxwcZp
tjQ2BOrg8+UVD0OQnPxSw82O3XhWyEKLg+Ots9L8/5ssXi/Le/EAQQF0K4c6FVQf
pGJcCmC8N0Q5DDRZN5+/w2f6G+wl5j3UMVLjz6bIdwrvkeoK3IFX0FGo4Ny53CN7
cdT8c/W3nq731uldTe7ebSRTu6C3/ieBwLLzy4Xr4HGK2MQPsBCIss0+7aXcJKeq
fkk1obicHeYlL+UyIGy9Cf80lD/18tdQPmGjfJN9ZfGoesiwisQmyEU+S1gZBGib
4kXmlr9Ue5zPzglj+bUdGMAFbdLtb/2hHUP44f3rnQIRhUPw1I6wuuXpkBsdG9Mg
8nQGKvsCN90I1w1zgvbnzBbLXLVcfImDhrPAY/qzQSEiva4KsXDOvXYDzBB8BB2m
1seAmXYaSV/0J4LONDjy8Ps0IruJnCPBvAjtNa5gVkdbqwRYYQwqLHpCgBUHEhnf
CbbPydPddKb7Fq9G1IDTp7GRsbEgWXwLf0mpE+RGNanYnYgGR00O6i4wrf5cyX7/
HQXnfBZON6UsCGnpfpgd7clvs7j/9FTOeSBSU27zLdZirSqeiB8yv7nd6sXHv8wC
DiC3XNXbCe2Ek0njz3H8QsZ9L4mo0RT4UdSCtIF78a+gQeF9WGWv/y89eHEIvbfx
l828UIdhRHoBPpYSGid0EruvaY1l27QeFJ0ielgiWYLYM0ehkiZII4zu2tk/mFRg
BnQwh57QHBMn/1KhKRnOHVmQMuPR1DKTLkpcg15E9sqPEofH/hlIUKL4Bgu5O7Um
Q86RsIppcnLQTbMDDWHIlwA9Ps4iLejeIwGs49okB2Q0Qwabr3QiPHpOxPnm6Y3m
AlBxlN8Ml5QPMfiBDayp9wHyhM1Ta4dl2t5q/hywTIhPrxKmA1doX264n6CSCpnw
GCsGJc6qJDcJybfRa6+IGGRznLMzdTocwh0xIXQIXfLsCysUoefTE1Gm5BP7zpbx
rqb7PRPCLpZn2swJtGRyQahLVp9B0Er/CLga+iBHJYf7unDiq3VsmjSCysPkFjwr
pUOlZ3nrTjyCjF6hFFK7fpfvZTOBvlGlINq6OpLL2OI7fRvjFmsdeI4fmu+L1sh5
op0zLnHfyGhwbxN+KSSF23rmjTo6HxgSkxblBdXK7fwY7C6lSpvwXnKz6PbCbV9c
Hn28moDvR9eT5/4ZGMO/mLN4cOCr99kHxgEMWCKjOfmpGp1hAHwivsuIk+0ZK0cc
JpcAunoCLkuC8oA9nNPS+f83Z13taliSi3Budy+gBMi72g4O5OVIoqtjOMT/6NEu
ge6mhK5Tg5dDblGL7t/D2Jb8bV6mRnb7PLeoxNle8PQJbVV2L6H2TexKwGa60lwq
gKt04NiKxc83lqqOP6Rh0gwdPPKTJXKbsHUe4cHchp5X8FQxBgCewsnxOo38rZql
R5BIMRSmtKwKMD9R9T6YXp8U8nq/VM5bAkG/kJSiiozqALoKxGnS4NlaxM7jbunw
JIY5+LBEjEtiUAWH8Gya60lQpOhm9wm8zezqwtITgffNHDFZF8doyHDY6eTWYjIN
Ln/JP+D3cdihmkmUQapS2dfMmBmaE7LEVSzL2DjpEwDKaQK/Lu106cEhbAD0cphn
+Yf4FYOdMkCkCNn3qnwKi3ZIswT0xZcBu9BZ74QQNenS8ZiZxredsexKkyjFlgPz
KEIMlBk7V82BBLyaW1RAWYTdaHwCDDExAIEDQ9ntgZ13jPTSbARy0wmXRAOWMQK2
xamF+vNUDuSc0QcK0wKIs5ayo+XbA/gVdy+iS24tMMF0EqCWVs8ixB+5AUMfuo+2
yrX2c5BiM77pGn8ndV0YMiH36Cr7S3xWSMWfZHO6LVFEvnYNV6rVgLXJ+PnMBDke
6GnPI4Zo4n/HkxTJkLdj5hSqm7252fENsieJxHCfSGIdao4nfGVXZx1noHM6X91q
oe8rlUNVdTOFui8qmWhY3yJYgFuoVUM09dwkbfh86S9kSb24IF9caeIBNX33bMUm
Fzq6v/0YbuKmOeluTkqQMwtH0B67f+/lCAUcY4/JAoZsldVGeUfG0NJLgZ1F3miG
kPoF66/FiH6EcwXiPOrE3n2nRQnSmUFRyIKuYG7RXq/mikJpMIOeTcoWWOvVu2EB
STKm7NvhcUPzqjOZR6FPPeafauO1OzJaYAeBE7QSYIRpmInv46/CI8qQ8Zqo2lLM
v8F/d0bIr/ZZ0e8aXRrhOkS2udG9Tc0Nx4/Ij/NsN8nSvI6Ti+tHwxCH13io0FiV
vIUv6jrnzQIlB4hW2Va/q4ff2oB7a6j9eZFSycAmQGjkPVFuwoMvnFUk6lIA8c+1
bIEfSp2naxT32sMF9Iw3COab5excfGbYFgmDJ1obDo7gTWJ6tAsv4APXvZoVekIb
Mo8vGyrTeC2I0u+DNV/2lq1uKMZPMVIE5QPbDUYUwrkK8yoDFVa4q6kyXV9shHCR
pdkU7IiUGici/MV3Rc0cXhrnsCXW5+tA7bbvmdnY2z5Zcq8rtegJERPk16T/m7RG
vWMVehoeaDllgu2k19R6fWymUvSzyXkyPZY9/JUDHljJMVPf40XzFM5rnQU/NYEb
/C5idPaYvsVqMA/VnjdfkFIJS5WLAqTf12u7zlaW81iwHqwNAtQE+pH1QPrxBO3d
1PajjR7l3b17rSiHWex2kcc9MSQQiEYE3Gt8rD6d9qn8csAvE1Hau20UHXzqtCom
5R/VCKA+ZAONzGZ9g5NpZHv6JPhOTY+BN4bRT4QDyd28q0uhONyzZzSQTIoLToSr
+nON3tmTl6mWeNpGdolzqn7ET8vJ1OCN5yqSZpVd/dQRtBArCT+WU9rQlSmH9i/E
qv9/JU8HErRbnQ3coNAd4tSui0ztxps42h6lbXd+iTFpCvv/qR3nsmfT00Fp7JD2
9qHlV0xRM/RO35Cb4uul0RlAuUeV+ELj4dcFGbccRHMowWJqWB0VjGjY9LqsBrG6
NGQSkdWT1aI02IGouaC/Y/RFSJyNPv6Bxzso7xrZScLXZS4+07IfjPB9QGdKfDsX
WcaGiEh7PDuRDxpju/4jurh5DsdscFSBPZmd7BSw4JTpuMMNWzCTSPawGm3IBdSq
UmAcFfNZEYabnlsEFgnKBvuBD0HN3THWZg90nEIJ83MFbzQUhn+rjfBItomj1KZj
7nyoHeulS+sBJsxPZbCjY6DcQs4aXO7yQt8ONYoUcJCdbOiwXVzT8wZxxXIKvfPp
wsnXVUL3eFAXKVeX44GZQ19ybkuIktnNeZE9zHLxn0gER2ebtZo7Y69qY7XpHP7m
TsST2AURNVFC1aw87W8eJhCmUHqDYxSEvK2s5lwzjrwrek1JsAmyAd+KBjh4/YM3
qHddOvdFnerQdmWdEWTLjnuK5jUgXUaZOwGzM7t2k+o66tg4wPUR+P826Gp7TUc2
sRnD5IXiRQZyWHRGOYjbh+jI8pbHn7/h5QpIKInVdJ4srwU3xg89bY5bxOVEEhzb
OPYvV6IoMdVStpr/815kp0Uq+IbHldwApSHj5M/xqIMog/3WoCu9DpKWaShsKbq1
DFoaDbJiCIhLmDP6mWqT0qnCIGcmtppm54424RhF9MeKfEo1kyXhteqVBIzPYnlD
AR1m0bT2VSo0ya6AIv21vKQmDnrWLbf9/zH4dqQKN0TJD8nc0thidem4v0/6SpFw
m/TCHiQIhMkPgPh7mrgDwuT31RAH7PmxhNTwaRs/uyxkGHi+mp07xhkcrRObdgoJ
Z8wo1eCkbRKO9nsxgmG8sBWgdWNymqasizGVEK1+4AEI0ohL41x6pi06myUoIvds
y0ejiEzbEMpqXIRj9AiRZmhjHXIGxD+PGP5mHhHX7xzL7Mj9Cmm3jSHmnqMCkR64
2mk1r6eD8eFmvlqUbHHQ3RYdQNbYf2kwxbbJEwgMM7zrQhEklYjct+C3FZNZh9xi
UGSGA/WZfn2kDfR5VpCnvATPd1ez1OhEaxvG84OUcBRMD+yBg8IpFaB3qY/ho0l8
I5fB39QpuBxja2K6m0PXYDulaKxEa7s6dTMy2nxdOmW4nM6oCFDG40XCydT9JPvr
gxhw4sYVtcL8IWzrxZ6VMZPBEXNbQoeME/JkkR8PJAjWboDFYwIhtDfU22UIKNZF
qjQiUWvb2tpmYBkZtmg/ciRoOzQrr7NfgR1OvBXhIJ4Aclkm1SLVL1Em/XyH40+g
mwI4QclzrZ36UFl2mz7NrhJU8CS8RKpRIJ5SwMeo0WXaT1H3KpCAPBQz3EDRPiHa
kiYWs8HJOO4hP0svarlO4MNibgJRgHPnQfKMicoOLzTA28Vd2sl5P/JEzIeGqiGt
hdZIqvLdU187bTcFVrjAcHsHTiZFx/SHnagsy3d9mMOmnzLBj/DDxKYg64IeZ9A9
jp1P0E85RPwfxM/qfRckYUpgCan6IbFWYRaqF9LkyXNsnOjiaj7hNyy0wxOJdhwC
OY0jUUBesrFDVZhuLsPUICwA+WrzynaFJh4ovvJosOltYllR190/mTykYzOlIYw0
FxAn7FcG8lJFJ7QyTlIt5sxONpV815gUvy7akcyoX720Phy7lB+Q3zCfc+ewtOGx
tH4LOqqqThFXVpm3KMKM2soT0rP8EFOgQCd+9qJt0UEv8ejiYY1eu1ZqImjbxE+D
8VGW0oGeyF8JISRGGfxdKhed+a2nCB9TDQ1vz2MXnYFV9iyj5BT+v2tzu1KiAIAU
57rYsAC8+odKbYcn50KzOAq/O0qmd1iIguU0EdqNdPXAxd8aJDPTdERmrXNjQSQl
JApZJB7HyX5s2d+BEmpgPjP4xzqhD/Dio9ezY2/yFu3NRLbKcjrHM7DV6Lu45G5o
ATLeJEKeMn++ZqODV7pMruRTXM6U/QlS/Gg4Nx1IZNiaxsr85gNcHyW2EsNOZfRh
6CGqRqA1INbPCUFYSaViE8G5UZbPJ2M+W1h02/xzZcwbYlyLjVuZYmqCOmA1NHKX
cZCDl85zZyCtEZ1n498AuHAD9sMk1jkBb6Wp0V+3ES2VcTBGOlG6sHv8+8F+rfii
dmWAKOWa9WFCUr28TPlOoURxmPTKjlK7D7yv9CqNYycyislAmnm4molt0+VTTxPB
wjqpysoJWFGSqzMyJHyUZ21VuGdYQCwrrkzx5inoGqeo2egL7csuYlgh41r8MqcM
LsAChs919V9PTYUcKWfCQmGXTpSAPmc+FfS8m3kqYDwMcmQSdoGXPklPl8r5Wtgl
SmhkjNzmEYhLyueluaK38n8XRjmvdfrHMyiPH8eilhCyUD6inKbaqWT827gK9ePL
0kITkgo2JZY8b9GUj+n5+PDFFg8p+Z3BCJhSYuoE3OE5tcQGRemLh70mUnbFMuyp
m9jtS5W7JotV0ZPxVppZ8JcFPWObPwipAq1hi5r/D4VMy4RNZnX7ZXBZ5Eu4Mvwp
NXU/KAoYBX39M51Tws2qRAEOeAcrKXcm1azehY+CMdEqJLsnAz0P89sonv7tdLua
+v06oD4hlaK8nSuZ7i++oPjDiIN02o5FBQVpo7xzweywQNDuAegvyc7G1PnLr9Ek
xABtxH2u8f2z++SIEnC4XW3kzMqbb3iuW4Qe1M1YMFPZAQYjvF8r+ika+dvzUeg/
PZ76YIDw3eMF9FRQmluxoju+S4nX2u+jcLojoEazWWtJ9Wrm7hs02LdpGBYFNZ8b
Etnb2nnx7K0vX9QXhBlJshxM4rKLMqDXn8B2QImSZytMEp7MlVh/Je0PnhEo43KG
E63w9SCH3vpSBKpKVqsokoqNFxCTDKvBr5kcQypqnFrY069k0DDTdPQtZKQJGnCS
+PHIVhHTdArdczQsIZC8D0eei9UPj7QR4VuKTBha16BPlKSC8gLe8M3sYVrdcSgC
Zou6/Yb/n2rAXwRH/birP+N7fjV6BStISxkaFVwRMnu/efkRhKiMBqMd5BNU4c9J
EU2uVkenL/W2yWBCWHhPmxucLEovVFIxgg5aSDtfcVq6XogVZlu7cfAhkMNK6ugv
hYFaMfW5jnB0KCbAMEVOGXCs1U9re1aF3yw9xkJFPkq6P7VBKS4Pe6EzFyauQmel
j+ZogsvBX0iuiGs0u9JtAx05DYYj2ZoT1LBAkTDjukqjAjAQuoxYra+HfBMVM6wo
JDKhFNAfv/Tg8dwBqJM/fpA4LEnXk9ob1tDmYs1KUsKHM0KA8J4+E/L8fybhqnzt
Lemu2FpX9lJf/qIYOOrYN88VhMMN1Tt2LqLEO6ZmISk40MP/9obt+AlpD7NttDKM
Stio65+N2JpuZhjQrxOIwZNIRfL3KRkkCgf3kCsTTX4rQHnnSeoxr/TwJ6Unag9t
XjmG5tRQG7638rw3+Ey9vQPzuh8qXEtK2hCFbujAStwbd6izt4xXRslV1bGkdbug
UP9QrV5i4kad1Jf9hHjiZHaQ8jB8cX0G66o1jbhsmJJEkWE7XaFmdTU+MzjwAbar
xBWJQEjfNCjq3LfvrEsTpvyFUfNY4+nkp/soQ1ezDAi0uGzMdwIOjLXTb2/+iI+A
4RBGgCkehgD64AbHCL3K6NyT87gaRYsA4DZ9kBfkY1w9MxKyO9buF7J/yHu3Vpx2
5ZeOcrdRaOFbAf3/p5+WJBjFZTMiY7Q6tR85XXLUeSTCPQLzd/bMGq/A0BjxdYBs
ooRXD57n4ohF0MG15OhsmxAMswj+3J8BKHWuJi0pjHSKPN8PfgOZnd0Lpv9rZA+6
l0F3LEmw/baQJpzcclgCQBRPSJypM5MuvT91aGHgWCLgGs7CMPYLI/CULnyT5ReJ
6t3ZRIEDz/g7DRcQx51SALMfRtO1h0dulxdyiI9AF8N05gMJAkhNJmI93PAVllSS
kzsahV4MYF+xPmiMU242gCFw1J/mBWOmeRsDuYKjELgWMIyWnxTooseLzQh/MKtV
uM6oJYDcIraRnYomrIr7EFUKwEohz0WsbgTDEQjLIJyReYaSOFt2/a0i+1Jvd00o
MvA9cEdeBhRBAHwJhvAPsWXU0xT2HRsVPmR/WHo2uXcriZMI2gc4Rr9pLReQCzKz
1cOVwj/CD6RWp8XACbb25mU2lX8i7xqhy6JJzbs9Jf+mME95qjdsSFIud1NKnC+H
2ewZHl3RjukLM/NCWyVvAO7k3fxLFzuMNQj7Au6PlPZVYX1ic6gUsAtHJlHB2HcZ
VHS/WHD7d1Rl8I3zrYiYOuhtmnSoZop58o1ZYQyZJZCht3IEg/3mCIqFHsTuc8C+
SE97kLT3xXUpuP4ckWCoqHCHfhyMDrXjEwBOQFd26ttwlK92IvasGiZJlwO4oxhS
I7AFtOpap5oUDLHCAXwB1t262Y+H39NEWtb72l7J1iq71zedMc4LWioRv8C3fjSW
/1cOOUfibuopdLlGpgcwWHDhLZRQ+5TBUzMzHOLK2Tc5XgZ3/nKiX4yx9lvachXz
fGPwLq7Mcj0HkxcfgRlXZ9cYAtN4flH4hXcmD8CbjaCco7VSIP0wy566rd7tflLC
YKrJ55Y+S70y4D3qb/sDp/EGvbVLOOEdOWIc3Gcj4gJlGEM5aYcDvVLhz6f5+kwY
YsZV3TBrYLDdKxGiSXx5lUP+vcWOawM8sAYtUpz1ZHn2A7ETtvn3vmvXz8lFuXyc
c356bDo7OkqD19ajHpH6K1WwtumsrxxGStAZ3svLycrZOW7TJ3IMbTWBlpJv2+pd
QWdxCrwyjx32STKM9vO9jpdRCHf4WWAsINLaQn7jQEvjiCRmw7PueZmxKgf2sUHV
5J1S1eE8dSVayXwQh9FqPvMw1AobKdizGDgeOX/emK4DNWDc6l+04UwjJL4lxv/s
i7Ait4TfRA20/76+rw+Zs3QQPqs+VSWX0GU63G5RNDylwJtRGfcHQzvlFf2JYH8q
SXYLpoyKszGUXcqcISUbJztEc1bZJshuJgc7Mgb1c/BgBZa5VrBCGXR8ejqK9R4e
CrG25Q214BOB6KGZaSL4Yzqk6b7FRW/STgNjUc3H/6Gj99PGG9KJF8GnsPTp3LAQ
APMJHnWMwiruzwEPFu2zd1BaEo4qgd+RzEQ5wQmzo1LLEyH14BIiZmCbSMx/TqGh
cZGZu0LxGaUCiRQdU4zZv7drHQ1rqZOIEMhUz8ze4DIFKMS7sF7zC/sHbV8Ng1qu
iTzV10pnIvr4pDrJsHz5V9ORAWHZ8mNUCXtaDLY6goIwnnlSQ4IJg+G5YvXjafgT
c8fyGZ4zFq3pK0evdWUb+9q8KShYGsOehie/16ewY8lV6E1Cr04oTgkk+Zwxu335
oi8IkHldk4DdsjoxkcySA8dZ/01sqcGb3k3NvncA0q0QgrHoj4IKA7VVeDk3Uj3g
8TWDTFAa4O2Vt1ykW8et+mCUA+A2hP56RIAGylJ0u/ykAzdnYe/dyBVlcStCigVo
Hwe/HOi6dzfGuwOUShKTD3EhtSCA6lHAUuYpWgqjzOzSUNYd4PA6ViV5igG5Skum
9DMMRY/TtPA2Gzxox05OwiPuUo2hJadvqgjAqEXsy8D8NqLWh4d5kIPRd7QPo0tj
Lp7YEPOXMMg8WImsCwMIu6LdNxdWzexLmvjdF5JlJ4AplNCvnk7zMEav+wuYhGSa
O8cDXIO/rWkO2rkC2t8g7t6+2Jv70n5mD5u3KqK7sUXXZiD8PpRZJvCqv+ulx2TY
BgVMvau/RZGu0pttuJtTd30nt6QioNh4GnrT9vQFfe0t7qbsYPeVacbaW6nQcXXa
B4B2/2MT8X65blaiyfopVaCEDNICAbytismbYIS/uZg0Qzn4Y6KlGY4iN6/VOTwG
nyLc+o17gmpebtUPN2aWRBesqPIo0rMZ3ifWxLqEep0x6289g5xnQ64ofDOhxSuu
WaEqirVpdnzZbgSqej1WCUxq3DG1Yw6jKmsiMxhJcIJxJCpN5xB3wPSUtbwlJ4FX
ML6k9TQRpVmHLWiIWPt4cf/fY4GKynUL1gYpVeLLmqy2YsJVL3oIwIsUmD+QJSU8
OYzDRqp5OzrOAc++pXJqkIVASuCquSm8GafS9lVQb1wb5+uUtFZ27bmvt8RFbmkr
tjIRd2lHo49T8artQQUmk1f/OXv7HNK3l2A94PsPUnYsUA5/itl4cuMOoL7g3EsL
1g844hTs8doKcMCCxoETzWOv4d5+9jP7bbSoN75wkpnF9/Gpy5QP2/QB6vBDcjon
UyD+PVhPSX3WsK2WrSa97vt1rRSRsfP0Xx02ttqnAAcwCEQTlPNUnwZOydxPYvQS
bm+75n429XbGezDKiosGDEn5sl5S8oxtfwuuWS9wzoT7yRhPdo6kzeFsY6WnNpYq
zjYG9O8xP9+HSG6vd4k7BjWDjae//E+1FT9HGhx2aq1yLwIBhKH1L1fOOfFh50kr
jPwYdtw419uWTl2Bt1VdAzYBZL6Ga3KsGK95z4PlOK1CVx6qz5VQ54yZug9Mv5Mv
SfWNj++OgrnPb1R4zTUxU1+ysKUXMGUAKplmuwR4poeYC548V9jiklC83Xamkuup
rVak+DTmQ6w/7SvVa1nEYCT+5BxsvXex1U5BjCoC4PBSHmn7C2OLkvIAixaDbBB6
8/PXe8iOB10AzMo5Z8z7Rz5YNtlsGoGfSTJDIQXoEMj5r8ic8+/7PnjAkcAWn8AN
AAuM660IdNgD+Z+AkOKuL2FMH+U37vUdEiozTs+/6aujkEOUg3+fRoP9Sm/Tyi3x
4IPLGG45tal5LbkRzLmTH1wo7QasD+QZ7Tz8uZ9IYkbLAfiX9/CrO04lvIFokB3P
66pactbjN7m+yNjfgALtXlvSVsoajEn+IPz34SEXNLTd4+CxI66wFKAw/eMDT0tS
N0vKNQt2myD4k6DlqBZma2GOtICQVruFzAqUbu0l5zn8WG9B5P1sEfWeXfmGcKAg
J5fNeGl5HmRCnzzAOPaUyzQ+pVIjjt3YgM2lIrSPVFzf4OOK9+wAjZ/PNTuiw6KJ
Qw4DQt0e7e2m70vx+Ha4Hvea3OCIub2KRWN8K/dugikoBtrfLzXjlSwPiphTbq7W
i8Zux+U9G2QwjFanuF6TAseQ5HYBjOnFQ1yQxXAX9CXVpXfhrCWeMl4lbG9/Xqrq
HR5R1TYn6yFp/MnQJdC6leboxtAwXsAQ3sOpmMURQFb8GD8vllkr3ZORLyCeMJHD
vilYk2n1pD1Vb1dwS/4mCFE08mOKzu3O0mWcRlR/Ym324LeMnou6P8cDOsJ14MgA
7TFxF3rywPHAhavB3CyMpC87om8aiPsEX3q+zbW3TXirYRTr0HzxoZKxuMS1nGU0
DH1gbiHTe4mxRnV0Mes6q0CPUEmQh2ccYdYzW7mwbYo5p13VbLjHy0EzmFgEUppy
qXh8CoNfXvphA3DO2/K3J+ExyHUcLszyvkjW12nNMz8uySLh7Gb5llEZJz7ytmdd
KHr61TB+EeoTWccOd8U8wzD/ykFL6ztlKD+y+5ZVz/zjb2ErJiljDxVr/AEKhXOv
usO3iyAwpBS04SuRJ0QK+TZnpAax8vchTq/N/ZokeO4krJ975StlfjpujF/IvE2L
AM46kC9skAAkn0Cj2ys1LDPQk3YAGFDBcvkEk4bJPqogMpz9oZJz9hnBFVoGBREz
VBO01cIKVk2tvQ0ZWE4A4DOtIfjj7n6HlPZY39vY6RPPryCnKbG9pHkfSBwm3LFA
BYJolgNIwhljKMuAavFVL4ognhkd8cPzZG67XJnvyfdoaib+iqCTz4tmKLLQRleY
ol8XbJfJgAYDH7EE1bIoHOB4U/3LQQ/K0e0Oni/7x2m/X6Wz97Ss/MrOOHaKNTLR
VUmQI0Y81QXABfkKF0fvqry50uxA/KGlMbEpc3/w2g8vi3M4eazVlY03unyhXOPt
V3qtn1QFdEhKFquIolASjCKceLjnmM0OhSBWsQMCTdCycMemJ8ASXD/Yip/JT80o
Hrcwf3aZ9s/JVpx4VOiVlbeC5KIybk73vnAPlE23JytY2xMgzESlzQCzhI+v31cy
OpBSOT7RX3HT+vkueyZlsodcIel6Jz52TGC2qV5uYc6m/RXydNbFzAhcrkXNh5Hf
oV+8XHK+Z/LggD+NaOGs8gNJJsvODyMIqi6i6VViDFgtC5/Cv7y/0HaYPw6LAuiI
fprIVd6h7mQuM/ez8q5UbfzLS8Ik6VNg4Hq5eOioZBo6HpetS+zQGqS07iqfoVry
aZYnX+iGsRuB9dyw6kNMM8or5i0/fAS2mz8Lt3IHiXMaG5L9r6xrbTn2x0ls9PzY
a/8ZNi04Sshcce+2JwjxRYIACS4EfjHP00J+kHVbjF5AMIOpeahYRamiWLYMNN8a
ecq4T63JLzZ+GDB+H/+acg==
`protect end_protected