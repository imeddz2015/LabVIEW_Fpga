`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 4496 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/59UwEX+aE7FohaWu0/8IpTj7mav863zUNIsgIH2BWb
Abd9opeuBjbGF/waQMI2vMJTwD1ie1YueHc3nSNpEh4OXp8P5ybZFY89uyGz3ztU
W1EsuUnchJoQgbHZ/sLbgtGRgsrAFn+ZoIeGN1d6RAF2wAESJmYP8zw+p00RvjZ5
pBGEHX7wooDexzkaqKS5G4ICQhHwxvtVBamvrp11Os/SmotUQf7w51JZyhlaN22p
DrMUbjMAHX7xEIXjFdrlfywX2EvxRlvou4kiOBFf7GPcWuZRGmque3SI0WKJkgQV
MzrSLqKs/bXofSC3kn+XAaHQAjqXNOxqYA4U9y7xTDYSaaltW7EcRTUOdcl77G/H
7y6dFh5Fr+p4e1/Co/DlXiOgBVZvu0XkM71OJLdLrJt1cLq0W/dKKFyEvJK8nkcE
x579XrxqbZDpESEPVTBcTOrwk1elf090JEwHHE/MET0ECylgBxOGEvSOxTgeUJzt
3XbS71+PAoamVJvM0gziS6ui0rb94cahqoK/9EyaVDBx7hwkZyxQkjV7PX4hb86A
WUmak65vRKA2qS7vCVmKrPY34alrcgsnZAi51FrdhOl95QjuATxGmfcB49ssX71Y
n2N/NujBYMyFlCZQh1rjCxskeifnW6tKVpZ90dfTrasVKuLhc9/m6gydZgJVJc15
AZ8EzrQbMbOFSpnQQLK84GqnObnLTj8gDCAjWC7bZTGRCEHT6JgR3CiUSTINYqjL
BVKlvukyM6aAwUR/4dcNUjfy+AKvZLF809zwji/XOHoMOZAoLQewrFsCcjHE+nq8
7vbKct8zHalGxZe6tp55Lo4o5pbNeiai850y0BGA1pshUBFkLWIuM+neSpzlAwOA
8ObVJpSJCPzEEhLUDEEvCBzhVfcKnWIPm3LAjccDwcE+aWxbS0m7cDjzpjLuQ0VM
Efcafuuzg4WmZ6iS2bJQFCcaq0kW45P9rkivzWP3boXqRDldR0ylq7iq/Jb1pEzc
Q8I1o8s2i9eSgL0q/xJ4tQpHenlS1p8f10JWzqJxsCyOGgxzTFETDshQJZzDVj6z
gpyTKrM+WCOUPu3bgJwzxQSxHb/2N9toU9ZEK464JQeyGd1fnVcSQ+PcVu5NkgNh
hfDq5hoFB60pnzze6Uk+dNLEE+BVlhBVyBSYm5D2dwxb1gsfF8WPWm6QkpA7BZs+
JUNrFxC3nSh4TDTN2ygmr+JN4i9HQxF34nRhr2Z6pOt+HarlXwjYn2hARKzxmnZK
rSex0A3Nc6Sg9nKjIOUJpD9G1gPzn5YBTQwlFMG5tq124mx+Ba+mUH5VmRQqb8N/
heXt4TZQQHtD3Aut02dv3dpnyUDfWpuqMiqaULgaOicuwIaApArb+pO+ocwpy3oN
3h0zOm+4sZSIhX0Uasrjh0DK1xbOB+/GVb+5k01dXwqp9aTe5LBSPf0ywr50pj2Q
TKxhilxrAKvwBRzmUV2wq5GFavLMwnyiWk70+F0Vmd7Lk7RBjPYXGDeh60K9awJp
nV0qpYhFUjwEOuSe+dT86Gt2WJfUry2Gxxj9+YiRCgICCVjTtjZzyI6ON5QRHfnF
N5PtrsHLkvyxBFrQLPNPhOszhQP6BUtts9UDuDbCYdcY3Ces2UX53SsHGHR03P/A
WQ55BR9PAEuCZJBs7NmyonaZ4p55uqwJkJ6OQQs5YcGmtdXb4U6e2uDrptSkVF3K
1p+rXXJ1x6NQDu6ekVbpsV7V39X76yHY/F9f+F3LQbkg493O17WA3IN1EdSGtRDK
I4mnC9ZZ+eR2a/6ePsAMSDUliJ+gLCsUNEUwlUPfnOM7krHbRZnpyMIgxKLUE91A
oOcmsm6PkrQZoMk4cF54FtHfBG5wxaZs0UWpPPRPrjUxzIpceI3LedsLBA1LFaN0
IZQohF+90FQrPZNVu7rjAp8cqThMjexQVWE9YeAHkUJP2qzHFdq5++j8x5JCTO56
oKoUTHf2QU5y3faf6EPUnkhyjo9jKCRIbFHbKZbAe4hJEVsacyMXuCBN9uGqlmYV
MOSD6Y92sDvleabGE8dDeJ6IVcpuIDquQ7A6HBDSlbWrCKeN2kFfDNdbitspIq+k
IjDwsF2Ka5EFGbz9ypRaFThUHhgC/d5/scx7IibnB9ztlaVzu+SqLh8xEC5Sd8J0
LELGwmKkDy2I8KbSpUUTK86PX6o6ctg5rvy2h2gf0ZbtgbeQ93ZbMIAHkOwk2J83
IpeXdlNOMT13y+WKJVlIZBvR4TV3LpIp1DnZmS/j2YQnrKGNuNdwEAz/zodxgzJ5
xDhb8ps7moSNtKiFPuxIx4emLLCM8j2Iolr+s+h3iE0OpsoOolSiEEb3m7Wvgyea
+bpvkUi+b3ujsqrkvX7UsESI8BzSgh9u63LYwGzCfDfvdwazVA5k6icRNXwPE4Xl
f93QZJSSdrvlzHoRt+OyfKyCdhRPbs9H102UpYRsl5K8gLiSSwfPs47hS7eRkINq
tB4pheFoCc4e2pbnFv3acId4fupb2c1ysajADBpJLUl3Scfm7d3c+UFYeIR51yhn
h5n3GdtisTi3D0snOha/lo7s9TGXDibRdnI1vo+k0INZ7iquLtGVOSVuT3a1uD6C
+snWe1Kmo8ex1iRWrJaaV3NipaHJJgAZy0Szkzt73IUEWHJt+PDfejSvZn4ZQXqa
UgdX6RVQJ4F6S+qd9BoP548Gy3eXNozHjVEmuuHMyTLZfZlVDwHlL+LiGClTzg2L
lqIKddVwJtaUlNy+Ew+xfhBoayWtDxKYF1i9m0sA2SbKk32G/YDCrqmIRuFox/AK
GxABVR/g6KY74auFDNjVMSMwz++66k3b/h4HaoXdpTcJdMkU9Mww1lk8GmgG6vLc
+QebSqwHMI5uzxAQFjGZWvgWehTAfrJxOD5CyvsaJ1r0vTZTX4zDoUeX3K/eb8hv
1N2kamra1J65cUdBPnxvS+KB5sc1m5WQ0pMXE8kncNb4bjVVnc6byh0uoAgkQBk8
208x7oKqL0TZEWb7afPfeIZihTEFW178W5sqsfPli57a1LmLcY4secNDp2FX6L3R
6F5byG3bPpQ1eVtRpgt7ylTnKHpWcMdxXIozRvxTLPy/SiqfzDhnVPqss20eGFfS
YFCB9M63vGfc7chyNl0TF3GXd6sKv8tW2Ht//6E2NYDh/dEjUxexD7z5/41hmvmk
C2KWV9lV2XIZPbRV91q/Nv2H1c6uwsWfR6wL08qzM1N4bEyyQryVb1AeJaEw1DKE
Xp9Cd8+Gae+DVh3SeqR01CFAH1sxUwL3saMLb4X4O5kniRPpyh9EjVK3yR1scJSp
zPDDbamaRRsa4ItZzNpFT0rF+yoL+SVEFS83MQgVWw1QhEU+VEvYDvgmapwvpUkH
yMVh23VAvwNTJThzOXTWI6YiZ2Nj45f5yFM0NbcQW0mMWm0GOkhi6RYbBcK4+o0P
sYFytgNtsnGkl62Y/6pR/yiRFfns0GEkCxJjuYAi0fkc73Jd1hjwJgFOLQAyELxx
OZ/3y4z6jUtUdzxeR2FsmsXZTYrD8my5PTKsW0MKADBNsFHvwrhd2/5XyowMwX80
OtIHCM/RUmZiDL49Y8HH+Q8r/9fgGWHoVA+WWcgDcPN4Lp5umXq4fnBtZ5AODRwF
YGx8928uyeB7T4+MbqJrrKPZvREG6NHvhqiGHaUE6UDPp/de/vm/0/GliRZlrx3S
2woplFT3Jup1z25Few4kMF4vGSfb17JYf3teGcFn0FOQgKOsP4S1AevBIQ+GepZi
XTezvj4HPfJ0WucHcSiQDohDezfv9T5KjQGrHFZiIBq+A80BJpnV1GpJvRIVjEKq
A4ZC6IwFey+PHgyVhbyfysJgPpgdjv0T0oWKzAOoEL9xWc461b4wEr7xur/w+Xus
ILWIFz3nJUuLPhY5crVIvzitM2F/TCq/Fq0zKfdj91NBL/p3tsO1GVrxIf+wYpfb
FzaBlVPmwgMn1Kbsm4Fyzrr1x/6rm+YWaFiwCqLiKWDbvpBi6AHzBC/d+fzPNU1Y
zj7Y7ShHvFiqB59j73YptE3rjDdK7rhpsG9tl6Wh6FK6cIqYjXlJv/mgLtctEWBf
yxspH6nvfQ8suUy82VY376f3gC8LC1lSisNORw5mq+Fz/xueyF6HtM2RpwFbjZKo
Q/gxnEaqMRBvaISyPkOVwbq+ZiGT5RhdkEyZ2R2kegOZWowPaNZPJzx+3+QfK5FZ
uviO0DdTkHT9CKSyRFJg+qx5tYYpqG7qOTghlE2oH5Ame28VorEH5+wlOeuT2Ai7
tBcQJmINrxbqkN3jDyKY1sHsTTZ6znJZ0CKdrzE6NCwxCq2Jyybgz8U3YLZJN2j/
prtzFhqxRdt+E4ao84+y2jSbY5+cZiCw6qcYXATsQ4Z85hvgdSdPvw7HLFkHV4py
Y+kR2ogOrN4hdE9PgeJsZnX0wX1LYaPhYK01mz8flYtqckU/OnrniP6rmK0/V5nW
BbmPlNaf7cbfTLhOLGG7DXrItie2gIFhLUu/v5N77CMUKNUggDv8fBV9fgbgiUyj
dWEb7r0aUpYWj6mBkqu6PhtWajP0aNh0u6uQ6H1OfzM5V23E80SRtT84gXdo3hqm
EBPGOeoQZLR1LTxYaBzsuyO4PYHZWhJhLG1VB09K1AV36DWj12TFd53+34xwsLys
7Ohbxm1OIX5bdgljCbA5nqxDFlF4DNz5aXjkyZWPJwhc+lJiTaPZK5SSlhw1WkzY
9WAaBXBABWFAjX4fQAYg5xAU26PyGoQvXkCOTG+fHIrYv82tm8NXbNbbLEfMwPTD
ZZHHbzUltXaHirScPGFIqF+G2bT7oOSkubGOcXPiIJ+YrBXGxQL9DG3jFJTheA97
8BUGc8c3k1fV+8XD2kBTxCJSMhnv3pnPpZtI9sNBQb4XXCLHWTQFR9dx6X3GwqWK
QPLAbyqf4K5isJAIkGK4+wujoapq3Y/L+A7xZVhg6ZXih/Dg8U1MMyVs7Y82Mcz2
/g2mOUpgs3hnGsQwkQ1Hj1zgiDj7HRSiC2L0hVepkQ006/uTDX/afPJY9KGZ+Caw
Zr9Q+8jQGj3QzcI4GpU5dldq345qD2a6H7KRlRxbBnUuTYcvruZtpOZGuEzUpoCI
+vmS0hErScKIxEX9e7ys8krPP2m/hw16D0aVT1Ty/QRuwPp5F4O3z/dSDNcyKUpD
q9jGHRpIcX0chHv8fR0rrjkIh8/R8KLoSQBHTUkdXUaQEjNBMJ/X7V9hExrgWq4V
ZopegZjbT2JqrVQTDMtxI/OhuR/Hm4FXcrhuwCnsqHpItZywUEMTpjEkPkxpjrJg
HCxe3d30ZI15VYGW5CogIlQZ/gi+w2XbvN7no5WN1jNJF2R+NZszwiJqgVUbYty0
ktVOd5rGp2zzZhQxFNERLevnNRXUnoy1Ju+MB6VIpIdjl9arKIvVBMAAHwv1Qw9E
DvuoWynNfOtyMLlkpw46MUvKmj6H/CMTWJaRIe5VSOUxeC21cDvX3kVf/RovOP0s
8jyd9K2RQUnZMiVLNhn3Gn8ir5Qe7wGmK/gWV37v8ARoBqb6CeduDbcCKKT9xvos
vE9tVBzqc/vaYB13WV2Y3sNidsI74ELRnW48XDqcHEeIs4+RYCtjR1JiysumEgbf
okgxpNHnxRCdcKaexV65VJP9ghGwDLuGWPzu8YiYOWluNJve7CT4F6mFlZCMqD7x
no2t0kpN/wi2fLsrRiX18n2wfoTfEFvQHRjZgLCQSrPd8bGbUB9FD7xwQoY2lAWP
nmcmDUwDzO4VX6NBa1JjL6ag7kUN67pNdMUVKdHwy1ogxZxkNqEUqeWjhLR5VJJv
Q7bRfanx4aPKzIJ535hRjs217HwbV65lUWjtYffwiT8icUvR4c2ypT/ynQtTIUfW
eO1VyoWExDnTRdEJk3BnJbuuJSHtXMci4jIqNyc4ipqK/GK9FE3cBxMyWY5YMY3C
QSaGXuHpmGhlOBLpp44uF1s826ughRGa5LuON84Y7Oc=
`protect end_protected