`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 10720 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/59UwEX+aE7FohaWu0/8IpTj7mav863zUNIsgIH2BWb
Abd9opeuBjbGF/waQMI2vMJTwD1ie1YueHc3nSNpEh4OXp8P5ybZFY89uyGz3ztU
W1EsuUnchJoQgbHZ/sLbgtGRgsrAFn+ZoIeGN1d6RAF2wAESJmYP8zw+p00RvjZ5
pBGEHX7wooDexzkaqKS5G/Abg1I9DB+g7tix9utv583O92s5ej51plXD4AgkAJ11
VDv55rTojmZmOEJXmkY9ioP9L/kH+LEf6pwYjSgOa2f4xoLxK+xHQ8L1Jzh250Rq
TGxLo0W++rp+DuqkEJwsBtWwr/t4nKkhxBmmtqr//+Nh6jv8mwSSEvUkToZ7pRgO
z4EVfV5sS+F7uF31j7h81Z1HfJ00pf8TtwxrfXuggnffScdNrTIDej+bhv1faB/F
16IRuqxLK2OZVV4LqtEiahvQ7p2byFEfH/2ZcL3BJzIqAvdCZIyaAFKfCGIYgvUg
9r6GWtRGne21zFExcB3V57sn6hEofBjCMRoaTZSH0nDW9GHWaXkA7a39piXF5d6m
hNwpG/ji4EHDRFYTNb2uJgh0V9rJABRzupBreI39vgy8VgWbb+CpZ/H0FQiP/4Q7
41NikqAwqB8CCeuOJXlGqoqRom5KxD+us3pXMB18JyibesKMYoU0ZkoNlK20F7Dx
YhLcHfy8t3kBExkqpYBWqKNB+pCFYp9bVmO/3jwh5xd0zIk5lROg8GHGmnN0lW8X
8rqQQh2XqAwKo2euPWbDKFQNQbKFn9x2SykI0TLewC5uzMtvW2yfRAUAZ72WpT30
5QIi7oNIY3qddIKjdWh5m3HHJZ+iNvn36dMZMTLW4nKPpObzl6pbVU+RNqQ9SfQo
V52OKTLzqE4zMSAsk8A2pzsorVgXdtA3afmLniMCCwKcQFYvn+9CCZk/25+xJJ7R
PdfZE0qeTXfWEJkBBR4lqimP05f5oQnf4vInkhll9tKXzfNly/N8cZ00fqJB8wCw
p155XzmzwgyZo6nxSyImxVr0a+6lix6JUPW/CKVzgH2HZVX4duhQG/XNh5gVhuX7
IWqgwX8ptGMU52Mh7RchzA0VX4gOBB1yqV1RQggad78IaGass4Aiuk4X18OXpg0X
DG1sGF4C8Z7ks5qaby6Zgx+QP0dBngnSfc+npDuthc1zBkU4HxLCVWYpphAHTmkQ
fp2oefQPfIIHw3OMm2smVG2JVaKIdJmQyFSNJdTO/Yx+Ju3wFxX7LMKvSHasOnbW
c4ucPbiq2W/Snv1cLfEuYDu8g4sLLp/4uURhEw6r/TtoNmaS8Em/e4js1mO5xa3s
W7CZ60GAS9qZB6mhYIUWKPwch0eJgruxXE+TxPV36GWJRXKkbyXMNIa6sGAZl9WE
YMbyJJSRJkXNqpbLZy76C5sgMWxzNdyKapOj7dDxwE00hCv5c5939QMpFhQtNNHF
78jWZindkDODXNhxxgcCLlozVRbCNa2E3SAZbnYhAdTWXi1Op8OYFC78UK067afG
cDa00V+ZWNB35suvtQ/Im9h0y96OYb7mokHQUmb8FsIrCruAik5RpsgnfeoBJWDG
YfGHnOxBNVI2m6E7cp2B0pgzKKt2LtRCgEhEAiEiu/q3XzhO6Mlh5s8hqXEG9zZI
ULc7a6txUVL/LzIVG1KRT6DWm0eY/pQgyAhCCL7x0nTEGSla8kzoaXgQzY2dUEpG
UppWF1K4qdS7A3yDK2xcjf+WztuQ83n21uMNSMo+IXJRjrrZfMzumBCPMmP2XSAm
Brf1KonN7Zt/hJpWaRF2K97/qUigz/coTupHQRan8BK8ex60PYdQgZB2JKSecUzu
AhIv/QTLyBVhc2wg80UYXdfd63szW9vny3Dk9nmxqxATgGHesvzOA4C94ENy+ALf
RUKfRd9jUuGArJvmZCPKcCuz/nFud/KN6vx1EfhiH47akOdYUuGX0t+DgOMXeLVx
M7MpBo7pYLCPv4TLVMgdJL+SjSY/q3goJm879SzUQ0RcjvA142e5EleBUtiBB96E
4HNlVcvznDa2o0Wjuzpu3QBpbofWv7dE4l1baw7mb0gp5IfRk5wL+umQqgpZeGpY
PmvXEDDPDv88WKQrWh9X+uWqgcdUS9zhTzmGKRGdXC0ioR/0Z+Wkw0sh6kHzSbqI
7VNc+TSf0H56jtBJAQAYZLZ8/kecQGWiiGK8nAwVFG7AqCiY7BPsDln8IW+Pokz5
NR3nKej2/rfG+Wjg1Z42H7Owx+GVD0jN+CCV4BniipX9L91v0vufvhewbPivCKaN
yr4CNpqaCqEVhM82VuL/OrEGsPEYVxGpE4ygd9Uuo0GGkbQiOhqVAT9+pFrhdM+t
tQWOaVw7HtZvH2Ev6xNOq0Vhwq52LNnxlcZ993mw7tK3PBk7jW7JZQPJS8A4P0K8
30BHT+aCApn5UPzdOe8p3JgvoGn/FWL/asPt3xmA/vHvDcentkewtXx4rNaI5UTY
ubBYsr49fhhSIY5vkkDHWHMc985nDrjwqcMPqBGdRUqDPvsLkI+YqyYYcokpQw5X
gj8dnaZgGsbWKO3+CLDDPfiOwMBIBLr2sUL7AeezL7yH7tH82w409t8VHW4Jzgkh
OlFsqEJvhNRbecVkNbCoKVjWpObGD0wh7bDXsyMfJa1cA+EvSypapB3kfL9xvc/A
xYuOfTPIff7fZ5w/Oj293oYDlvN93sslrqdbf0CQ0cRZCK5UDKxkRzQe/0QeqRDs
ggH3W1Bx6holWjAOHsVT0gkvhhbj4XjjEBEEuHypdFxVQYtoFgh74Fk6OCDEmxYq
ok2+meMOQaaH2usBGzYcS9fucMQ29qpkgluW9lUKLvKIgwqsTzB5Yv7thVi5pLo3
OdJLU7XQlu9kjvyjerkA7Bk+5zwBDIMRDzH9zDFuXPUA9QH+MSGjBGZSIXUXyKbG
+Ra7xFhuyU3vTh5M9tcXhKJxayLkdMA04VJbpAnJoQf/yO+BmVGm1njjS0NZQ9pP
NiSB427a54Pt2KgN9RNm5Cz1Lzoeh1OS24QwyrhS51oh4dJBNiCvkBn4iIL6njG4
euC5xh/OAhmkEF5Z5GS7k2DBG8+Nb2+OIuPdlzONxwmUi3e0C1A/h3c0d8LzY9MX
lAiCbTdzMFTBboyXPC1ZmIFE4CkFAjfZXQ7IqK4hrqW0L9+MNIlNkXkMEvP1Fhxi
buuLb1s9B9uym1p+d3VSJm9LLE4aPIRAxJ1H8ATYYiwGkFuX4icSWz/NpNhylqeq
lH3V5CRT4myBJR6VYzqg/eNdVt6Oe0qSl8k9GSnBwGtkUBz9CqsB9XS1U3TszWJY
B4cNZVQ4/KVvfuo/PyVu92jyuKWT4CGrU2bUYuuYsXxfliQU/7ffNfBF0X/9b0PH
yjiZWpP0y91vo7ipvgT53f4mpwBM/v8AyGLLfyJpYPm4pLE/9gzY+bfcgnwZFlrD
TozZ3UcmAfO8AvxNYpEdvNbPkOCf4ZHB/BpPnIY81yD7vWbDgETNwI7Gg+ukIgr5
Y0h4s8FO4xtIA7WarwOp4+7hn/Z/rZe0+Es95QNvdRPXZEavlPuA/+7TMpg7MjIx
gd2SWH5APDgYF79ePM4IfpG4l0z7ioAxx+wmbMSM+wRYpK08mnLAGI4fu9ZOZART
/p/VVHYfq2rBsy7h8t+LD9VGYlildMXGzspuvGM9YAs4DWSDmZ7bLNnWnd40UfQG
NCFseIu44Kw+BLrEPPIn4lfsTN0OFWYsocLh2JhwJU80p34Z6Wivyjd7BXD5WyN7
B9amS1mlrnTGG1LEjLo83d5ybLaqiTJeVjo3eepA7e9GVIHSD25JBBcb672G8xsx
chwdULNK9zh2M60U2+6Da1uqqOU6DE8qnLCQwlgmvyxpgXmqFuS+IteQMmp1chtE
kyXxIhDdf+LjPDfQMuwwHyfmp4Sx3p2LAZ5opE8p8+zm1S68d3usPL5a3MeOLtoi
b2G4vuRqCuH8eUnmqSq2tN+11nkdWmhi7XTvXe1eLQT6ifzL6AR9C0qfc+I9p/nV
mmM4Xhvuy6jaH5bqCsS++9GmT4eD7h9CGm4dPq7x+0l0iSya5V6RpB/tEgo/i41E
NSfSMKL3aXeJnH34Z/auaZrDJ5Higsvudwa2LMN0VDOMAwzhVtgwDncM3yJu2N5+
kb/U1NM7UekvmlJQDdfcf0OsaLlpTsIVg07RT5Z5eALe3Gd/5rcu8Pz3tlwEnLKO
WWUV6P9SWLWikwDxzmd2hURjjc3VofZUD+hS8iKKZrer5qT8gjVQI9WKYJbM5aL3
mvcg1EiCKyo62F04dp/pvwQcIneDgUTKiJJ/YpSXwOUgqG9rOje9z5qP8vISOaK6
L+AYLtq5eZ8UwFiZJlDGAF92BuYobgWxSe9ivajY5Fl5TQ+slKFcFKIUf/uJsBIl
ChwrsoLERmUaU1ppxDhktnyt1oI2BizqGR6f6pllmOsvBYYTZraAlO29g3qj/NBS
zpRwWxejzoM2U/M9Mai77GmtPYzD1VPlemu/Jjekvzfwc8uM+oAJI5m2tbVYjltz
sye5xcmvC2fJix2VqSC/GE/KHX4cXOtYQm5S/bZbiMnCMLYqKiwprboogd5ipVcZ
L4yE7WMj6cyht+PPpmv4b4fTHwW9idmn+fi9e58dm8vfCVXbVXmuOtSJgN6BHrY/
J+rM/kkcVspIShRpR9SsQ6wkL1hdA9IG7SMXB+f7cLXoXNKnbRRsxpTxZJz1Pn0e
K0D3mb1iG1dtIH/0TFFZXKeZsTV1/gb1Go+lzTpqFIV9F7xAs8xgPEx7mIA97f78
Dt+xI0C1xuA1VBghLSF5KMvvtGw8u+XIRHT+8gKbqVwWmu5+u/AosTN1d+z4W9ci
owvHJuDyzjhP+NnYagDCAWOld9D/GO0U+JLpCmQtxliU0ODLKE7aYTj2AWj3DRMo
OoeXdFlILHk7Ru+gFAiVPFUxBadzl5cjjoeVPIZqfivI1HCOuGDLlOf2B2VYpo+u
hlybvhi+Djzi3eyICE4rt+6Ef8elzGTpS+E+7IWwWZP/HSxsK2OfRZLmqv9huL5R
lzw4v1FyXyLZK6Suqrq85+sYTIUGfb3V0CXHG9IzBvuwnmLRpftCRvpsEh5A0OBs
TbFWO2UOfRrstz6xTpmmKsXAXTqbw3GYKn5IiadP8WR/cTpW7aP1p54q8AnA4caO
AkjDN8uNTZL0XUIeSiApsqz3rbQHF/DUmMFPTjIqRPbFELVtlFvQNIDMMXTx9OXj
Ehq1zfn5prrAi3447Ld2+rDVcXQa3XjHQb/EB6PLtQt2OKjXMp9ewoOWvSRvTf6P
2am+gHaxB962AE7b5G37s0DJqLtCRwBSv08twQmAfmSNg0hk4511nnYQXwcK2MQM
/rYmHCz9PmsQz3VsxB2lD6kb4E7E/gUhdigazj0wN5XA61xgDukLoGpvzXefIVFF
BeL8ml2+ziFQP7EjSetRQpQq0R1vscndO/zOEmN0Owic4uEuU8iLPXvjxvHbEXFm
zq49p93ytLJMEZU423NPS7wGydpQ4xzh4SHMGgo6nCtxaTOkXDnkSkXTUc771/6G
n77p9EfvsDzcthXc36rx+jv8d9SKGDejozB1nvmS++DekqtKH8RUT22RCj++JfA+
gYqa/0lZZ17P7xwxIv07280TYbAl5zVzmdK9u60ROULAEGsQml27hZ39YgQmSY1s
EpNhbWr+5Huk/F1m8SYQ/Wc654jqrJFMT5pTu0mmewvpVELfhiXMMzJH3DB6PRIV
dxyMNSc43NrJhVBXixPOe1vPim+Z1pJidvJb5QCK+1tTxhXHfPp3WhOHdoHHoKgm
y+vOjnZMEJY/kSXL2kUnJNfx6nW06ZUHS1vhtq0GOhw2Y+gEZCwOlfm/0Gc+ChvS
r9Q3jQfr7HRSz0SVvLLFuncPWIbi+nFaRNwWQKwk7YGdb5rZLqBstgczlzx0pX+J
Fr2EkLEMwLBwg5blVVZfof4gmx9l9SNd/LedjsAu8MTbPP9rOHjohwPrQ8KnjpBC
W55HaPmvZT3sL5cSnYnmxC0cb7NZzEbxvfhYhMrmsNI0d9thMi3PjbMHM+iesE8Z
XejLYfC3aMpnLPgQM4NJ7X8FQ0EyX+uRjxjO9p6lcg7h9NfF7XMrQY8AWUzI+4uu
ebMfgugs52OVucII9kaofeqYDcloglGORMB0TqtJinlJT/KHSK+cIAqk2ZEHk1rq
JHHaaAHmySUFlWxJ+ewLCYtqO/tV5ibXXElGWkQBOe2V8Ay55JR4mmSO7SoJ0XNF
9HxoEFSJm8UDZ167CrUZbu1Vijqcw1fYmLjZV7N6gK9PIhE8/54WEPqQYXl326I+
9GnRxLkrRP0VRPquOUdh10cYAPIP6X5+UZI5CXjBZv+7irv//DhftKsIdbhlEgJG
ML1BtammADSQ/DAncAiq0mNi2MFT4XDJjFBshpMfWoPefU6wO3KFyRK8ApdyRh/I
nS1K+mLn77NuCoaY5WcFb+Aqn9FTNsGoh59Zlfrh2h/f7CA/mq0TsTh3GwugwOPI
lMlTr2XrVB3d2S4InQthHfuQqtjw7CPAldAzXcqb3u82bHyhA4aoxorAKShH2DVe
6Gp2ILs7MRkl6hn/H0q71E0LNxa7GmbfofTCiGRI4O6suAmFcRO4GnWSq8yTrPxC
jRK5eMpWGcyAECIRTbG2oBsM7DfSbEjkQolRrGMVTpJzo89evoaJFF//MJ0Q/6iP
cuuQa1qfid8v10aWWLTxovK2NK5rOcd8ksBkCd5mA/jd7CZWg8GCpV2Zz2nyf8Vx
c8af5GPjyTU9muGUkIczHGyxCXsb+uAtxOhMzIIuoD1TMO9YCYdMTE/PDxWhKpqw
aY5zy4Vv2vFAdT8F4vRaXR4h4t5gEk7NtL/wtj57XQQebCzNUjY6mKgQADQIxy3M
F3VLDp3OZrduLIithZyRyAS2H7jeR8GWwUjVb2hjuFu1rW4TLn3ZLr//k3IiaGBW
gYkIvHK20YRe0VGc24jpa1bon5tdEpl1Sqhzql+g7Uigfz35AU5FylrQKCurc0A5
p8hiWQ6ruEq7GzXx8C9U2Jd28qQe9v5WrlhYu7U6fIs1GDuhQESMavTlYaCMvmfF
vBBt620boOIt52Sng9hq7LTgPq8iUUrEpe2GzSj/rqgASmlWfZjYGKGaWKAJsPPP
9KvMvGfe3dgAwB/yC9gesVS8ugRaPxGl/1Lx95TSYSlUMMMjjL8Jw6OqtL04N3X1
XMO139d658lFs6e6mxXH3EN7ZnzHl8zlre0gr0DXT8h7HZYVCKrYOz2x+5/rXuTb
Oj1Qm5jtmVMUAt6qPS/eYfheSfiKKye//q4J653Mv9Uk12xzpESCWazbIFJnrplZ
ilKMujzYifSICQ8HxmH/5bi0ghuwpnH/PTDjQxBE9wHFr79qgVrrEsUVDj+LMoqG
GJEUkruS/jI9zn3uDdYR1uaYX+Fr2AIQ509MtrJzRTWdZEv1ODWoEdFYTtNIHQKd
sBEgKqdvW4YbUhTeRL0VhFIV+1HMoYpTUZpa6ODkJiPbiK3+CFxSyEH7XY+VLkkZ
cZQfHFXLIvYVrJlqY0dpT5y9jtLZE8v8GVy84drfuKkmaDYpTzNaQHHL6Kn/W1se
+LyFLqoTFaa2sYTZ+7fiiJZxOtgVXiQhNNo6y8Is0Swh0XLTNP37Reyv48868D/f
211NEFan+8VE+OQ7jpmgla8p3xtmotxAvE58kPiVEp7uHmN65ziZOSw6E7cKW5p3
K1FDu2RxuS0X/bZ8YVNPfwW4+JNvNmUHiAA5H80et3PQH77HVBJQoOgzusqDHw7I
zQb1l8RYlTKkR89KxTmMHnNjBr0YyblzFOx0izKSHcGu/JObV+4BJgBYDUqybbD2
sq6VUQqxDvMkSCOk4u2jtc55tNAXclAdNMNEcmvioRAHKq5Rkg7HLLF4nzT9aQgu
Vqo1CT3o2rGgdNsoPKODpzm737I+HbGEvw9CEpIjNzoJA5r8GDTJ7NVw/kVfCxSV
ZsqybGt87K2VIcBArpDfxdmiyaNcg/JcPTMXg0fSeIaUYlm8tDdmcjNLofh4YdVo
4BPQQJWY4OLq7g9TDpqQd1I4Un3+xfrl0PUJhypGg/R1ySKpzS1aMXOcvT+Jx1ae
k3ZVyIyZquLtqWAhbt01jxpapvJU+Syyxt/MdCmnrUFdQ4uqfD/4/VSaRlExsB4u
CsKKNmJdstCjIeaIpuLWI7HOnztaLg3UI60NnxJgE4RNHXYKJatSKRhDRHWq3kVn
9P5PZTCFrqg8gt64J0yox0LKfCQt+KuCrKmGLxIzPXbPJwDI6+1Hjz88XK1wv4nW
yzAQOKO3ZckBGgCoh1cz8ov0v2XR/H2O/vSqD1qH0vsCTXJmhC2uLFszuv0bw4Pp
uMAr1crm2XfCo467n8C8g3PW+gaHdMhyfczfhfsFqMcuZwQUruEma2GXCDynijg3
C8KrvakE15SaYwyiHraC0G3wiiBYbWjQ9JljiKA+Hfu4nBDtpIm1hr4yHl7SOlqh
KQztSKljE6ith+of6cX+JQQ6XL1EAdBi2r8P3MHbAyn+07TTF7rOIoXkgE+aRWHq
JGDTGWfZt8XKgE0ndg81NWb0YucbPthqWyFUtUoEWlNdh6jpsq7HTb0IR2VyPUGg
m8f1384nptBVL9hW7C6htljcuSymmJNMvq7xckTehancWe86pQ3XiFSboCk5xKW8
r/l07KITWjR3EL57lXlprcr99nrgAkltmCI5MQ4MOUR4r2fBMA/iqK4DRO4oBy0E
hQGU1dzTGE1b7IOXgm04xFUVmBtWcZuvXFgv6AGf/CJ1xr45wofVXsDtUR7NssLy
uHqoI0sMORm72ALHwEC/toexigqXIpunGt050/uSv9qSl6PcGAYKS8VxWn8PUs3z
G4xr2tzF7srDMMJx5++/mhNO/s6LRSpzYUpubl/RrW4xWW7E+wZj4WiRPfCuoN8E
yLHdekZSeBTW3+Vo5cW/Xp/wbX1is7gPch5VxVo/4BeKzMdSpMkuxILht/f2jKvl
5o3GGgMg2p6pCD0PxHHX7FsN0kIb7h0731PkHf0GspkpkiUUTXfEXrDlKjCRfFX7
gsovMVSAJa04rmD2TmRDUTt5nu1VAEuSf+cWcyBLFnrYNFRNCWctiqMic8xOfrAV
lYHzYiOqbO734FDhLWW0SzbMIBzgXE/YaVvGQgsTRx7Ard8hjDzvO8eyK6cDeiJR
kzBpjGEH8AzNHMexokMHM7JRKvvewCVHcfZ0Am6TlrGqsQlaM7Nmm2RXAo/0UK9H
uvtIAqrL8VwGTW0qm+bEAL9U1Jo9RwvqRk82z+eaoiur/O0Zl9zq12Q4o/7LSY0m
CqIoPBrODqyR+fSUkEchV3+J+GUDe6++PYeUTdSonvxJnla2KOpLTN40EUwbD/aE
sVTKdmaPWL+Wh2Z28R6L5aTeETAQ1Y9j6YQTCmiD0798fAI0Oiz+b0NuLH0NF8qN
QcYM1hAmvsKrErzIHSyvHimmrCZlxG9UNk+L3yaF9R4Zv/4cyzcalbaZVvzCO+y6
Ka1TeOEXvV+TatnWc0UighnVHVKDrmlxuUMIzjUgvD8HxkbJ18ULZYht6kSMFUbM
wujlpPNWv9Ns6N8BJtO6B/7ldZeYhdirE+h2j2nik9ol6b4Di8e3dLJUiQ/8YkP7
9aueEd07BV4sA7YsVEEINLtDsFtY+YmmJgAUoHaYjD6Psq8/UmUPVHPus/5C9+vd
687+S12PJ43EgxuuXADKhjFrdP4Rw/4dUuITX5ru1hU0T7XussngeHx0hvaW+6F0
YkffSav+Uzmv+2Bk1sWNoNeYWNrw8KLTf9kDQjg82eL8rGw7n1IOv/rl0w8ivdQ0
QnRsvy6v2GUawwmN2/n/3MCCoCU8lOoWPikZQVU35MBDSWlnIkOlxTJ9rwCHV3iv
xFA1S5JokiN8bVV7Xz/oOp/BOdjG4KwroFU4chD7WKxuTKbWYMWequUaHWz6v68c
3AGOtK7+M7uvLb4T84jWUJimrE0bXaKl6hMzl+3OJeegox4wRGL4mMMByjFg3wD6
lg+RkPZH76pODl5LZpRitdi9d0wmbM0hA+HsWzELT6rW2YeuZZpZz5PiCOqUxrHU
ONQULAsGt9uhIHplF7a2YHA9Kl36LKcB6BEmqPf1F3kNU0tymKWHcDoFKRfnCxQ+
fC/0DPpHfe6h9iAE35JH3tfkp8FNLi01GGuIfCXm3P1aj5tiPkfhuKskUmDcORuV
t+NS4Wb0s4e8wyInd5ieEPndC+yTr+warYaiYl64W93xFe9NbYjgi40IA1YRloqV
Xi9PPKNdEYZASxJ20Ax6wvB/dSBHtz20adi/m4Ilgl6sncqvO44BUsohTR96XVWz
/ICmPGA2jhzfJr3HauY2HEWjiv6+ij4kbmBfo04I54TB/1lOTXP0nfqOJGp0xgZD
WFoGt+vbCaH6i3biGjQ7oFLJkyI8K/YRsxjfj8/w6TI0BkuC/P+DLeF66j2v6v/A
tae29FOzKJkYN0mUN3iMX8rj0QtKRd9a0xIdE4bfDK6rl3rVVDp+lgOKDD9Xlxb/
anoPdn/+6bOXvE0EH2xfEYCSGT5aTmP6ouFPJzpENc9yC1cz+LoSdOdNbjbeR7QW
xl8jOlNsG6khZGt5F260cAQ2xdbJ9o9LWCmcm0aS1jbH7m1xI+LvqLFuI6dHMnYl
77oZ4ctMS2BWtWO1b7JC5R1CH9zbqzCGTbqtGLffrBANgRZz7KrCZGUxUND8kOvv
ay6eZWTBpa4xMCnAF9sAbGzeCcVpWqnYMPUSAsMJ76bW8mKzc5s3tHv4AI7g8A1P
S3pTF52Q4BD1KUbV+ZOaY3fFxBkiIj520coQMJXeUnGU2oqYjqPayn4+KMdhV9xT
2Bf6+f/jdrSTgtW2DchOIrwF3ECLKElWxtzwIqVkW00NqwNlzSQj3zpZ8blhHcqS
Qc+My3FyR2Sm6GUwOBYrz80aGjTopE6mSKt5fXy6bHTTzNvPBQXpDA23zskXugTC
WgcpJk6NfDS6xvUa0d5S9lYRd4QdAVXC5HduGHXQsgPLpN+WNfbVksRV19aa4Sgx
3kLVndtgbNT74aNtTIjgaD9YFLDTaUxXUozam7hCLzI/5uo+CKcgGYBYfM57jJre
y4smWqcWPESg1lDmpUGdBRfxP6b3PhH6nHYjWb4BGrIggp8yE52olZfl5RBpkPQo
QKrxZM4HgWe5z/lL782CBJE7yRPMWF/FgOX8Kprpg/6RoFfjVYCV4bqa9WswaZkL
HAZrNaDlitEI94E9QBq0AyLJ3Cig+H38Rs8SDLSwU9TZQGBNPyDXcV9cq12FzHzt
ysCAH++WnjcVMguE7nXqRQv2sEys73Z/7w94ARVm5+PYHHYB5PE9ONeKHNStxcsV
KBXPfS4yFy0OkyZIfjubf/qm6sK7wxRgMJ9F0RYKIyWFYO3iVkxwZWqMmtmUYSQe
pre1pUCVYv1D6Vunfo1ghNuFQuvlxIpsS42JWWFgRzJ+/ydOtbaxLzUC8MRS9Pkl
HTjHaOs3DO89yQ0lGhqnF22Sb1OKEWrakMdJj1dwXSjZoSMc1n4b9SKxWg7674O1
+wrgzEKKDC+6M75be0kYJn7s91OCjAvGLqihTJz7gb59XjqebkYvBLXBMmjhvmVE
B9ZBTR0D6s/4oYxKNpXd4GUMXCsIQlRcw5yqhCN1pGFeI8oFE+4luBXEKBU7OTWP
SixfJ6ha7bsw1j+0sMdgYppDZ5SxdbAL0etHy2/ni6V9XT0uOzyv43a33NQYIewP
uMy5t9b6lQDDJz0DDpoGuLiIdpH/+swhPNFn9XcnskBV9iOhnYfRB+J/Hp34ZNwO
4BkrUgSF/zYxBUMni33xO0akFTHcwxTgUAya5ap5tZfWR3sfRe/DltzX9wOJZ6UU
Tg6GhOR5ZF+y+lV4lNRrAF05kRkjXcRgHIAQvDCDTQLxLI5S8gtLPno+18X7xzXF
7/ySMuwkQ1ZT86mPQzpFCU0Ikxyi16ZWqb1XIKmPcVm7rPkGiYi0XZqdlKDZk79C
bDv433kTrl0gJm24t8lfIaCVHBe0LHUlJjwl34STW/0VLZf0kd8YH5sVCGDgJkof
QM5jnT7IfKyzmpDr+ZsV/bnQ6VmxZT7ztx8TL0YC9d7vrrWgEt65FBbp4qtxVfLY
jO1Tax5f+w1muCc+suJLIuLM17bFCZNpDtpNXjW4NKUZaRbWqs76vmNC5gPQ+pv4
2hVrOHVg70oDhLaP2TN7PzrF+lJzRltzqV4i3xbGo1anXZPzMTvMQfrEmRmqMES8
XM7mETTi3EYTdV8A9MH1HVgap5tYovGgoM7f8imJqagqLWx/NIWOz4CFtGRoqjBm
/TrKgwyZD2lG3NSl4X0/IYdEby+h6mnwTYXW6o54dcIy58PoSslwLwB8E4Xh+P+f
BrlfnEjjpukiZdtioXrVFd3tC48uQ2XYOHFWrGRfYtT5XSAxpkPziNFN4NAw8p0W
b7A+kkTerCLdMvryTpmBlnQkJNWcQbt74bLo50PyETuA+z3aKb4yxgOOJ5B+9pSI
fbyl9wfP3K9bHDsthwvO1pcsb/TzzTWJL/nkxroTRHK87yySp5g3PU2EyjwJ4HUO
0pe22gjl0rU3nfNBTjfAcH3ohX3FiwnjPWvF+XqZqp86Wx65PrMW1mAj422+B3rr
vM0wB9nW18C7kkMnqcdMT0pUoW2WURBKGkEHrYxmUjF86ARXV0PayrudmwkOQnvx
i0cJ2MucqSPx60AxM4cKTX/fJJfk9Ey1a2gDXHL5zZ1xmwIXA5UTWA5//L9R0o0Q
A38kEGPAzvWWSAzCGn+tprPLS2oRhcnyJtJ2Zdfs4OFcTP7Bb1J3imkP3EtoYsT2
qNDvmc7blUk+UJ39K/QEx7471je+/rRKq/EApl5eDt/1n3LWv87gRTGdlfkg9ibz
q6lBXYNaEoG1a7A52hwMZRhRPB80X+fZW8gcRWsCi6Sdr7DStilcqYroqdj7Aji+
1gFtDDvxOKStvFxTwLC746HOfSgeB8997k1ba2htMmOmMoNJpJ43MA2n8TGvgMTG
TBllyJPAXcp8LvQPDGw675wwFu9zZOQfVg0QIrZhFeJOk3AqqBcRMpYru1wdfwxe
yd4GVbozVeYOdpaUOkt1ka77+Wvpgm6YRKyCi8rGr8QL9PozFaCUZfxn620rxfdT
4WibmfaTZKTyMv8NZICOBhRUm15v9tY1v92Ii5kh41kBhvPrNzdnwpv+lapVGvJz
SKv9kMQPrndmutMDziF7Zu3QBssVndHutMTApXsr/aIctPIsHJcXnxvW9+Ua3sfQ
ZlmLIjgecyBushcxHjVuB1ztsbFNVWvOPhfhRL1jqBOxq66jk1sYwPwkIfEtzT2y
aK5BJuFoqd1zEV6Fgf7h9BzD5DaXSPO/qcFxiODiqeK60xkj1h7XDt0SkT+ZsQKY
zeMkUM32rXmFFwBl2dH5jWGStP5LS1BZFSG7GDHvklQuJc/L0ulKXEfZbE1bAMoo
5x/0G0bCW0+8pVGM7DqEw0DW4NQiH2g4m16aWa5zgWZSXCaaoZe4/iajDwp5vS1p
ZipCmm8EbEX5yHFKbTqvpQSSMTu3JrqeGH7Xpl8sxPmv92OxU4wZUvtuwWqqMCNs
GmXgIs0w6F7XTkzPzktCk8GSuh2LJndmv5YMpHvVX9ulNqxI4PqAaeZjRubthksZ
KxyjtFgvwZIoWiAAmSdI/65t36Mahj6Dc80CTXIuj8GYzY5IXaG10XjGEgoJhL8j
QFlPihvheW7GxsPK0NE1SUAMJixaYFXY0h/NagQ0WMt8c3arU2X2DenvWeap+lxz
kCxVrzHJFe0tRVdtvVvvtGy6v61D72Nkxkr4PBqG6R/rvo0eUnIEBox19DLEMXEQ
qr2NmHAXzmRXE0zdcwmdRPlWEEPScPNbxO0lps1QLaPRNHn0M42KumlXp7Aa8TVg
TOUJHToHiBexQKJlq8Ku61xmAHB8EqdDf9EZvfd5weaLi3w2I2ZKaPPYUAaBw11Z
XwYTF/S+vhhX5RTaT2c12kMTFCjX5MYoLFe6PKow7IxMUWzid7yqzNVm4HUSl8oN
QZVUqwGpuUGClalobergEH8igP1uufB+4PQZ0SdChgSf0w7ePn2qc5cjE3G8A26r
K4g4CBs07UR46woEi4IRFJyFfPChK8elwVcksgj2gtXzThvFHozCwbk0WwEkqPOA
iLeVksrL+HCbqXXHT4kBnGR3SaYqPXgXCL0o7dR2tWV8HlgpuOTbtAvrIhhWZa6S
o5Hx7Fcj18Rf1JaXwngFsw==
`protect end_protected