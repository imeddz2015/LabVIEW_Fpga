`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 30592 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/59UwEX+aE7FohaWu0/8IpTj7mav863zUNIsgIH2BWb
Abd9opeuBjbGF/waQMI2vMJTwD1ie1YueHc3nSNpEh4OXp8P5ybZFY89uyGz3ztU
W1EsuUnchJoQgbHZ/sLbgtGRgsrAFn+ZoIeGN1d6RAF2wAESJmYP8zw+p00RvjZ5
pBGEHX7wooDexzkaqKS5G89Hdhj/xm4TeM0cDQKacmOyDw34+N1xDhaU71Et4Yl0
rR7rBN6gpMtsySm1WWrvlC3tiqGZodWo7aN6jPWJNa2TXKUM2cyjKRxpzAA79tS1
DMwPr8XhR/CpJgM/FD2GBTUf+NJFMVRF0Ll44k4A/f1x14mR7TrzuQ6KDQbvHQl+
hbw42OsRMFd18X293eAigAWnnlXhsyHiBUgCYWtbvMRe+hGxlWcLGyA9Nx+4hfN3
h1yn2p73DCBK/Zb4davtRUHDa2Jkja5LZj4ullFRnQCvsFz9VQbrXya6vq41wtI7
Z5YRcco4/enME8+CGdfA/g331pFFuzTbsDGAZtGRsRHTon9uJ6L0+TIc5JVXgs+I
wBKXtkKR2cG3fASyFhCjXNT3IJD4L6udzR0ngna64skKNNl6OtfQMd8LEIzTE5LS
K19W40V04kz08vSY9t4JX88/12d2fJucyHqjlMXz1T5tKwg9z8U6HwN6ibL1JFdn
D3Hpxo2Nkn8bBSrdtphbQlDMfzd8bF14l3o2Tc2isn6rGbOUvmst3q9Hd+4/Zmiq
uPumaw5RgnE4YalQXwdHxwJwTbuWV3zfwAVes5aY4AWiF0o34JOdYu0+rSmPiX4M
Jl1xK3Ym5cdsCYGKb+i93LzIizad46XimbXvxUXHSKShyMYiAf+31XqSLP6MWuNn
QZ777Bi60pw2utJh3UW8OPM1hrD8tYMzKtqCCSBwDlDRFxC/zW9fVbnLne/uKl/O
kcL/IvCMCnZfcglPh2U3eB0EWZ3Mcv24h7851eSAmclsCm1/vs4li9HX8SKNCv7a
7Hqi/SHTqjv0/oadOgI6U4ozmEu9QVsXP4UGxJb4ZJOXk3RLdRWdLoTUB0STKfft
HHc4Aa3cuhRs9YGOQdzPGx7WN1cBUdMzLzYteq52cUIR19WiMVsslYJaluO/eGV1
4c/SCfn1FpyP6nwy0g4BdE4S6egeHHf7EUFdYDDEQ3DxgClPsHFVtNKsahoiGSfL
5hejIUjDgfiRXVOXhBsM5fpgxeXoZEom89OdAE8j0CwGcUi9iNIh9INSEXfh4XMX
fw4+0LIh4NgdrGVvRKugmv/B7MUfU4nRcsAtbDlQYgYY9sFpDHyOGib87p8W7vJJ
5jmLvTOUORDQ8txUvYfT2qykbjX9na00xi1HUQpAZD4kcrXy5ym7WcFFQSIgMXx2
t1yuBtFuIW+rpkxP7W4G0BzWla/BPWYNRZ5YoivWRPcv1kriRzrtKMH8g4QTPUqM
HkkkEHIl4BV9GaXxNJPbNbsIqpN6jb5yOu0ZmPPkFLG/lqyGK33pwEHWlPx1SYVM
zLndc31L70wKGYqDTAdWInZbGRgOYx79JKkUWOgEQGK9Q9Y72x0bpIbQ6aEB+8R0
gt/f6A4fgKLDNsqE4i8ohE0T4VMXwCLjqnXWTRdsKxM0Dd4EzIUvva8/ZpElH8oH
SphgFoX1ixEmgY/a7ptKubZMXGDKhENfc+rDl6EG+n//DTusNVszxMrBWG9G8Xja
pxIBoR1d2rdXJz0kGmORGANPUoKwP87Hf4Rou0phQ9lJsmnTV7o0ycKNevRfMpEV
v1u4epjedfYaAWPBdeDGOSdRVbiGc1Or+r1PIjnMqauHm8IQeI1XSofDjpwcsS4H
v6kLD59QwjR5Ad12xT6WsisLgZLDXF+pLecg4o9gKwHG0MK1GYLOoMN9ekhiyCIM
hP/L3VcElgfnBtmBMm/POTzoNiQWGIFuheAbpIEYMgwRlu8Uw71RlDUmYc4MynDG
r303/+YHNLiF5jhKbuEIVr8zCami9lGNVo+oRiZJs3+VHjuFqDE1/9ksz0qTYU4O
P/zHqSJJAWlfjHh3GT5v5P4a0KIcOLFZxJ+65WvjzTGe0NaG9WmqkTJOwQD1BvZV
55XuBkq8kwGVqXlbvrivv7kQIvlbw+RS2X6+P4R3O0HQQjcRYvtnGz2W8hn/OkIO
EBi3GnHn5gXtSZ9rdaNZLDBGau7Ip8gYwmupY+MaVhUXHUjQy89AJnkeekuYqluG
6m0GluPs59Te/roXRCCccVeijez4cON+j5sua0wTW3Yy5KHPIv+kaGK75UwcXc3n
85AmwOchw8C7RcXv2Zmwcxc5AgvLSG4i/zz94EIti7tkCrYPnwLmwdpQccmmDdp0
DfXqzlFZyJQGOkxjCLlMsB3oOan0YkpfLcckKUBX3LrF0+3ooBR3LVTiL7ZNxtjA
NWdDrJSeRf+xMqGy5jQFOjDFC4n5KHCJMSKfrmIf/7rkaT50LRoNCM5XeEl3Vcq9
GQf0HwYpe6BrcWvsBv01JgleQeDxzTyRGbNqPloZ9z7w7qvJPtHEsSrRA6UXmygV
pETJCQmEIBXaJhS5O4XE+K7wMCJ3DHhjnzGl2FqfaGRLIHFJCDMK1pkJx6MKrNM/
Pru0UEoVrG3KSA8yxl/nKu4EX+BSraysTYZuBv4ULgQyXWukTtqqQOsR4/7jMMQ7
0DAvmcLDZQWOgs3TWBl5c3lxvHC3D3JjdqHW8IC2HIl2PIsvxm2tHM93g0joZWrM
guvDUb4rv7EgWUUSQymi7xTa1GYZANv5Cd5T/XBTXpFNcSJJl7c3KY2ioq8zXiba
tNJ7RSnGs++wPmE+9z17WnSvQPibBoy2tllVmYlwzDgLhH7uQYSR1ZH7vTYkgunM
HAtQ24l1WZnGvJ1q+sekJ02+L5PK5kqtnK/J+P6STq5AC0MjUOXIeoD0rcqJCCvJ
+h/KTuKA98BjWGSig7t2Sj0bhzJ3AcKyDhlYChICpbioJHHEoUTcvQH5so+3HCCv
OV4O8XY12R2b2HYiA/6/gtNohJxhz4DO2cvIipmqdqmANo59j7q4LAuta8OJDGmy
SND9803iTm1HbYKwOJg1/lr6LWJL4jcZTphCKh3wBG6YoaGVXPrbdavgyRNfJTg5
uWQrRQy9YqjGJ8oTdqN1SgMH02cS8b1nLbgA66NQdbjdqNW+UaI4HSQh9tqrv1Jt
DkaL0lDP72reyBJhad9G+4tTkozTdExYQ3gfNRbYaVBLoA/uwb1l14lavpksoHMr
SJlE8o0/uqnEBAtZcKKFaAedJfSu+XU2IWAGiAABylxmVdaySbGokVK9TbG0UYiE
uF9RFV5NizgAIBmMx2ju+hSppRrBtU0PFigBdNPoV1d4CeUvtYCWT6xaXF12GC4Q
PsmqnDHWi5ezAwPUHYzRQSqfcjBJLf4eAkgLJulcpNxEuu+1Z+mWrWkPuFbyK7pm
AjoMuzO8irNTNsY41fBm57izHn7vvmqBz/4Wd63cpiU2dchw+t9ikEiA17JTF63+
g1N8moYICpya/VL6P94nlimGOU4g1OG54HaF/KeWKOvaAMfg1e97Yns7owvmPpO8
XmkiUEZzsrgx9PgZyPbsnKTjY0lh/PmSoxyNVLDNNCG97tIXTzdeTQW7r2ufygCU
B0Fa1wDJULT/dxaM49rcAPnM301q081jWW0C7JuO3cpuz663Z0TdP1TVZgkbAmxt
dKM/n3oOWRKRuyE319Jg0gw0kd9kgqLDdD8w0QrxuV2eR7ksCFL5tqNDnqxlzU4h
2dkF7LJV+b5K2VgljTVnjpOEpCySH9WvcBaBtxP/UKjKJhp8wUYprYy76iZ/jDU6
7IgUrEMycNzSIpUO9AKoUOPC5+LyGoAQuk/Ba7gJ2a8ocXxozEEwd+Imdiu/rHk3
2FPsh5VZVtNIaesf9P54WFpUULdE5aic0Pdtd0lcdwwlkdxSAeFHTqDX+N7fF82M
Z+9De15tJ0sTaDGalDzSnQb9w7iIAfxecNOcrGvG5VtY/Yuhrc7klcM4NGlDSw5e
O4cDUpEHHm6W4omooCsSL4isgceFSU3Dv5fPkJYzaRW0Oxr0ZLSimXQ6v8TiyKpv
C9++Fm2UtpCP6sRPpeWDZGY97K5J57sWvY9ppyBGz7NFYE6LXNN5k7rxK8OrEky8
9oD4bEgfK4FoN4cCsm8Bh/akQ7TaOGzeEG8O/kPjvWart0eJC9vvh6I6QwmxUf/x
7FsHO5VlNMWsy8OIbpUG1GtVQGo+nm7XTZcQWYF5Mm0cUNvf99RFv+vM5KtnegAO
WTkqCY9pFMYPH96Z66k4lsyDlnZ4coTTvPUpYXhlN1TKPfFBHYJevpFYNVzXHTuR
LEUgr4NvLtbBphA5sDOZeRQIV212JPTMKxLjqwIOhxOzGDfs3V2b9haQnaeP19aW
vI2cbnv5NmwfAc8/rVk/QbQ2Zx/Dw0YMQIJGD7YZG2m+Hcnbo18PURjcmpYEqQza
KbD9Au50HdWAaFiqpql9bmwcPv9ql+44f1HAx7fRu96gUHvo/qv9ptkJZdCN/5VU
sdm63P6NFFPlLUFQ/k5PoU+eiHOj72mUEMfxqdv107dFbLwHCVY8PE0wLvk+2/t4
tnEYSu9zzJgPis+haBxmZAVpVq4WND0VjSLrlz4RFrp5CeTZzn6Qt3NkjjijsSWz
SM027rTNqH8ZV+YTjTZCl9LcHgnxIcI1dLuMgZidSHLPlkP/5TOOLg7wqAOdvH9O
nwsoOuxccHnc8hbf4rComkkJZ76IFol/IpYNfw/mVQNp4DJWSmEoSOjk4YmvTRze
c5Y29CwFsn91Rf458CLHzDTgeYXT7p9Ivhgx1iTn4ert/V4VNF3fN3dgVvE66laK
GivjhvGc9HsHQAPGDeFpfIN7fHM5X+vHnOxR0od8RbPD/yNzreTdoBrynQ9EcSGY
5/o9FBq5PEpSITBjAMAh/KNzrgSWaAq2qVTKMosPoIGPB1eQQRHfHzo9FeNLdSg8
rB7xj7c0unoimivMIEsYi2iyPj/SD7u/nM8N7uLHaImFhaEPOTipoeIx9jynshE+
R0TBoxtritiuhKbAKEo9SeT2jt7J8/HHMG2sCpNut4RSBEQtstpMXAkJv9fJfm7b
1vaF0PW9k/nTZgdcNomeQswEZQqXnSHKL83SpL5HSc4YIPX6DJ7UI3skoN/IXexq
GbhUIHhkGGAC43b8LigSPhdCvzuDKQuDUaUs2Qq8Hf6kt9xozcAAYLrpXcUpsqQ9
qS3zZwf2hqmCCV5sThO2iK6VAE9MNu67EvC1uvV8Qipw8xY4H7jP2dmX1sXqY335
IJNEu1o8akYEVud56X4KwM9FKyRFvfHb26To2MXf32L2mpan8fBhTBYYse49gWVv
Ncb3YcGW9j0ehpK78QUVanRfhjw1ENdr82hMeG6HONkXhtxCGJl1KEbJgIEEsDiy
z6fIQIYHHoTVk1C6kC/nRv1LOZHMmlXWZKWxlNJd6If/NfE1mqifquzWF5UCP2sA
wVvSAUtNoeJnUdb9T/CzrmUcnFwfSovDreci5+0HMcQaFwmCOb4tgq+yBaDvAYbs
fNesZ4FKBbfR7+qo4ixPN4faNPpd0tSTeXNZPEE/Qm0xpA5sbp27zqPW709T41XD
yPOr0deKlZcOGw1brPkJ/xaRKuB4cKZiw1aSJa+n3w1jclgayJIg22YMdP2OErU7
N8frHb68LS31ckOIAOesKkCz767cnrQqnrMVGMyr5zPStgZkOo7ipkoXCMfgAhrI
x8Bx0dhsuth/4obfVga6bi2OJUye+q2WtCKrqaPs0M5C3bz6L1zTsXqSxuA9TYDK
spZzjCPMED3nv09jXXdDQ5F2XTT3fin6ZLZbScOnAvuc0gtC5fNgqiKeyPlLsdAu
+/y7Wj6yb/+uJixGCQTjjkVmYTGB7O524wlNXxPw0cxErpmhG5DrMR81PMpKeO+5
kRLpAUFTkdSb++FtfpT4w6pDQjJFpP5eKf1qXmf7woHH/fxA1PDpqu4QxbUxWOHO
10Fp+QaNnyQ1qu15pQ9lnfn3c9jaKbjjuOS0rJUsU3gwI1U4kASoDQ9ihnojIgnz
gn9cxGmhONTLUKsFTwO1PKupo2Y2a9zdiOLSofpxV3IiEPQuwwJzKDFmON2zIp1G
Yul3mulSG7qNqxDimapWn/5IVq6MJeo9AWtImIhO9YeVL7Pw4zD27byNcX3JSeW2
NP+AEbouqnIJ4w5WvcdSRLQf0EdrEtMyhNG+MblqOkMGCUJmVmxZtcsATPg97duP
wFtM0sgB2xgWYyg6mehEaXHQB1dM/e9DuWSBTKw3oPwFfh4HzT6TRcL3OxXEUfD0
RN9p5hoYJQeRmVI24aR/Dx2y+n0vBI3el5PNuaDHta6L0htaBF/HqPTw6EK5eydw
2IlZ9aTahudn8kz//7+D6Gcf+bB533UEm1QfvHCnM7vgjZYohXm5dRRDHsYIu8b2
NbYHoeGcQeraXfDoUu5h6CGyrftMvJ1PHba5laYhuIYMQPdvBvJamkqikzgrqqM7
jsLxHQ1LhAQ3brjqIWEBV4huPuX8tfiAfN5+mwPs4ojLclW87fDqJ//+kPfWLQOs
uJ5hE3rvo1GupVMuiSpT8NfQFGz/21XS0K+nFpLKLTcFeqissovUE4yY7QqkU8/m
39HbMBzGkxBttockjHyu931X9vS6ziiO4RYrheYd/MA7A6OoYaQhJsdb65KW42PG
5SJ1bPyT3bjwahyiKBEUBO8u+JPsdCRUxjP0D1TTwj7Zl4HwnuOmBz1tfl+XXhqX
axs91JNiCrV+D7dsU1w0/i4+eEgAsKB7sUCFRsvMXfJt3q5ibUZSQUKFXgB7Gy4M
ow1K2nwr2fODhDxJfUbA/Akdn7ipZUKkmLsBaVrTc2gbuEOBJCUuOxkdKlVJjzaZ
eeJy2pDjyT3CR+7XlKRJ1XXFHoZ6FgWU9Ocxhs1r+7YSQlK00E75gArXA11Sw7Rs
Fh+o6j6d8WJHClFfFYXB27z198KDsKqk+NtBqcQUytOl4h00uopCCvWrdVhUi1m0
CutLur7aPPwoWiIw+Mdq1y+F0Zc7fMS+fjM/X3v+2F21eGjF2Bt2ENTJtdp8tMvi
Nq1+/ohT6RuMhvDUYJh1RWdDKI4sN7kVsyqz3DEQ8swA3be/HuQb6hHtgPTmzyTF
elYYKwcuNE6IfZhhgRUHB/6vVaMXKmLikdagYxGWNVohK1pwUuV5BPrLoUDb2Zzw
HYzaGUStyUicjJwwQO86d0qbsyN0wbHAG5woraD8I9hYzlwN75DC7JgneMi6y3gw
2u/FujwAKu2+UxQj/hiMUWpCyKCKV7i682uGbutzF8c9RVavUVKdKeTFb9pGayka
oBoHBUWMk4vpcuszqOZZSkW+lKEZQJ1kK7q9dYq3WV/+au3d7LvkLGKC452e3bQn
DcCzttKiFV9djJf1z8cj0SjWihUwVRDLzM9p+WDk4OipjKhlBXHskfR4i775qywC
CtrdamnO7yDrMIsCGQNrKNbDq6pZ5wB69GdKlHMXMeJNc3ax9sxLFlWlziyKBpxK
MLBOTZcXHooqc7aLiogvyCMg5tB+XxIHDBX8gGT60+mt5szVos2cX6YHUV38QAik
PyU1PCEVuFcNw+TqSTazhCcbn/Ysxtxmdn5bQP8nNb8z6lAfpQEyg/O3oAh9xMix
QrjsNpjFdwVJQgOkoIjmjeTaVLYz2MVogoLbdul47HIhaFCiJyog+mjLnb3OudDA
oJYv0xM/W2w4i4/5Pfl5pFDfbQGT5Vpl6rwzo7TqbplsfrmF9L4zNlvD3+2AzOcV
yoCNqJhechUVYjgkEVVgYmq62Cv4W+egBgqvJ4nkbU0mC4JO4CcXstt5uci2lYXN
Tj26FUwVicEyc3t8GGeT6JDbxnygFtkxoULBFVKqSJ61vMiRfgusKGYrBG+lQSXR
WNfphIlYzUJ1p7is4UIW/23l8Zd6WnaFq9+nhdHfbrMKajn3iDfR1+SZrSOf7Htv
viTYIgPDP4zrVuEJh2JwDBz4IC/I5KhaHerDJTGkPXuu/WtTXt4srE1rcseAFmGg
rwQY6Y0OM32ItjDmQ4xmgJ59k3qRxUGQUNkfZWpV/6cypxteDIt916UmJ52qkkpr
cCY3+5Yka1ZBpJWgapNuv3bgQxVQm5msZ6qYfsW7ezO+J7J4DpPwA4VRmyGORVie
fT7y+5yKX6/EHh4vLL759ZvHc4Pq13mVsDmm5IJAVwwJ7PM2MFyfh1o8hk3/2Jbv
eCh0ZO8hQgyKGPpW+u6OVrHjJq/4+XLONN24Pb3JQ1aOQEoy9ZN7Uj2dDlzCYSxv
9jIwOgIbe1s2kPCiE2TbgX5uRuPLFXstYqhXgC/jmRSGXI1WM0kl9bns/zHkDw0O
tjbIZzZdCDsJb6oUHGdqtVKBIGN7HBN+yJcor2JuDz9ylrPYowlreGLBa3rShsfu
HUdoml/7o1BDjHqxVAEkiSZ+rml+35CfN6yKRL2dBSJx9v2ijbmibjEvyQD0w8Xj
twPEk6u3/IEYjmeWCqbEWUjiB2RUBt9tTOMkCTDFLTte4ot58D2hbwGnitH2+UBR
P7KhyVSPuL+G1KrV+ZeIjEWlcURJig8AqbJ5DGyc7JQ3cKTSIe6n1GHAckzj4KcR
PZbJ1V6OldKS0Gob5CKOFmBrnmB37n7uJnWiJCCzpvnVvszGyEp0+M0YVc35cDlk
DHVWKgCUxFbEYuvRVWIaAbRyP6jWPabB1SYcbzaumKsTfKCjFCbS0rQCaDoZ6mNB
+WKgotGqY8IJRhY++RFYJxYT0xE8qVzbTHbk+bG84lKIoPUbH3ud2LRJlhnHMN4r
4N5WienNI6yY3XHyiUA5Dovrdb13c2ljQ+RQX9u6uaN5p/PYRwY8D5F3fOB6wb39
h2uffN4hDXlQeH05TRHA+ujQIHJ777Zpjh+ss3lh3RilwO+cy+YT1uvEirUoaKfv
P7TR4qoAHT//ELQdM4JxkRrRke1RJIgXRwKMagXfCyxAX17n58ClznZypFOueT3N
PjTTaT3d7epNuKK4P2AzL2ZhAwAKVORAYhGP22ktKap0uLycUbTswx5NopxpUnuB
mgiE62rpmpTj5/E5mmwZKxEKns95UNS66yBJlXwW9plhkL/giFay7iLQfydtA/yy
ZaHSu8jnDliJCsX93t8n89IXT2E5Lg+2PKpeVSwPCTJKr/TxUokH7xfwMu+dS42D
dgjT8OxpRmr+jq8DkSwIMqTufV4bROcyynbYE8FkCHxLRAr5iMZVavh2PKtOkp/J
k60UyqzIE5e6ONRu6lwijFTEOQM7orDttpHUAEBA7d+tk2gkJHbORAjsTKakw48D
J3K4dxYWykqKPaBpFne5BRpDHIUWtiyw/N3mpGDNo9VGkJMut8kmwqytWSCy3tIp
ZoxXddGaYk4SvYcXCceaAZJMrAHXLA0j4wb4CHyYD+xv5Ov0dNbdmJPfkga82JTA
6c8qTvm8dTLNURnOfjFVG0XdFgnY+WsQxW/fXp0AZXUGt6IZr2JfubQ1rhvsPx8t
UO+Cnlq8JqiDzXNZSL6qixQRArCsgF5R3X++osNAb61A5sn/JXAIoQqgj1sFk20y
lnxh5QMd0kC7Xhi9wIXtOwx0EV2pMW4iehx1MY/Utr/s+M7pXNZOMK4MJQYp01s9
gyVKIjutTmh+vzg6cs1YpUWhuTy5hcCd1sSCjAvssP5N9p19bbkjXEjlFowyh+vk
nze9opRQ9tsZwp5XktCw/GMvMwEQOaPf+VkM5Im7b+3qhijh3LpZ3hMjIYmpQq7h
X9a+5zSEHkKGpK0T+LAF5jr8OORi01hk677oBQR6KziyhnVZ97bgPrgxiMXKDmod
g/QynsAAnSZ5Ed1kkzOaYnRiPgEV1EyFYMJXvygl5NYM8SnS2hGJuWMzPAwXOpc6
QsfZRBRREyPXA2w6HcSzB2DTRwnsF1QQJ27/MgDIegTRJOEVkYgsIZyDU6wOJ9Nk
82T3/mh28zGa+1d8fMNYkafJbN3FDpr/c18cD3FT2WR2OK6/6VNkz7/+FNCJkTcv
PEAdyJexFZILJa858qDQZPSu5xHU6CrmCGL+l+/wsBvXFpY2kdQN8q4r75VbQO50
DAY7uFss4a5jlhlDl51Nac4lK4td8UfS+1UPvT3mCv8Z+udGhhA8aSo5cpdrLp/D
4MaKSR0//dBI1yiGk0/6Lqj7a+Q9N6WkzAOUORy1b/XrVMmKWiVxJQDb80O2DeNb
8RcnfS/AqeTpBOU7jKsHP+2kGwvC6qExGEofo5OZKLQM3h+DCz0jdmOYPtC98F9l
gwpxglpJA3bzaYVJDoD+06/+4iuROhsZY3kaaYoIg6BnGTZlHXZcat9tLZ/RoZ8Z
JKRzbfu3XnkqHU5sheYHzcBLvbeFxB9rR99tE5DbqYz3VxD/rHWE4Wen3gnxjAqy
C5qeFM9tBKLj2vH6v92ttKgHlMj6NfLaaUfgV5t9FOSRYPMBqMk4quUeXAR9BsdI
jTg973uSyeHDRm5hcb3+g/l0JL7IGGzKecD6OGmM6qV5mx9BrQ3CkX0oiLVs1u3n
sXE7rlO20ygiDMlg0X9BIanK9lvjaZYL9CE/6oEma+/fn473220FO1dwuBsAi3lw
qTylev1131IuekDXRBZkWspWwjW+f1hZHFcplZwNOta2k+me3sGINXIPlWJJ75yC
MHfYMPeDEP5JEQV7W8h1moKpYdouUMpClzr4sWmrn8qcE/lLpRT211oKf3RdUBmY
vGObZqvfjREm0BHTcQrUdM1ex8JExaHUb9xBqw5Ie1r5Go+7xazXDA1aVh0XiKEw
WKbLCni6hpwXQ1+w7Qff8EODXjKqXUPMIpwto4FniehoWEOYUyL9WMnwcGglrI6F
aJdwGcNyF23C7IN6u28NTaUtqArq6iygoWZ+WmM2c6SFmhcUIBo77yeabup/ULis
UgGR1NqpvoV2WtfEJ16Cw9/AwRZ7rtShXZhKILLXhZH1vBNBZi99kTk5WL+OqLLh
1+cVFp3WgTmIQGAVfmP16n1yoJP8YPK6B4ARvp+te+4z/g+HmNJ56Yg3NmyZbu8X
FD0Ny/p18wCmRSr9xZXAPSYsg3QTuN8EHyJUqW5+7T977OEAahR7mcilQYRpONMZ
smmUmvPsMsp+IfQkAr61nslSvyN3fZnEMzeC2qhf7m9s64EaHA1ho+8htZWqHGvz
HA6masHvV5awqgJe98SRFLJjHm05t/x8q032t1ntxy8gv7wC9MF8nBUSMKP5XDf2
TqkWFA+efuDe58IK6PibkkV91HIwHsBUEjh+cmRyuKvN9XukbSiit+f0JkSnxlOg
TXXw2N/sTA0eQEuKUBZPriurnvE60fh0NjfNeVNvd62zD8g21awIxgSY+JlG58X+
DYWeyCjWDCF2KuOt5u2iTfp0Z56rl6kGya49IgKBADbNEfYeZ5JoWg0n/HRKXIN6
nCT69F26fG0l/TfWBoAbF6I4GZh8mxdmWX07Esp3BE6fX9DUbVAHmQRA+uqIlyEb
Xjwr/GbWkefi0HFygRRkBMecKRvdG+Bq21Mg+/DatpjuUd/oPIkT1A785DMJ6I7Y
sq55ynG5/wMF2B5IE1SnlttYXBPpj0kjmq79Z34hJoABXo0Pft3JAcngzhJtaPvQ
MZ0mHlnC29/ksrLFfLRVm7Lk5J8Jeqs81vKXggqYa7TMPqHOVgeMLy2fF8uOfMJs
jEPld2HtGrSx9YRRlJf6mDy9bw95t8OWHGq29T4zNyxUBzvBcvOzMVqu2c8WKQkj
2O/7iZji3Ihm8us2gK1Ij9T0LPLuLZ2rGMOAbVN2Z7X0CCVDX/dyJ4Qa84W92+Aj
3IlKZitPg+728OIciwm+kVXAe05/50vnkIt1hL01n7mSW0bN26GXCM3m1X2ohlFy
Ufg4axW5vj2CCdTJOcHdpRE4tWaTg0W8K2AJPP20pWNtrnRjL68/ZHg6oBjSMRS6
6AVq4qNkvn/bxWBMuBoBZ9ZsYGEFZhzFSHg+Gxx79lfhRlefggOexP1TOuNjP/G5
/7llkpIWxXxc/EeG6p0lherDiG6lTIimsxWRcxmD+si7mrlUhA0XC0Yy0A2Ed+b9
H7rqalC27CHu/3z+h+jVjDuLbuYFYq1vMAHZHdXVRT9yQUVBBy6eIevDoOhk//hI
NeX4aqfCA4JF1sEDouenWT0U5ggZ6AmDNzwXlE/oyRuC5O0b+2eBJB7JLY0m0bw/
WT5lPRYvgTZutPhRtjHvUcpFTyli81gQLtsBreEYp1hxsOSe7uLBnpWfVeGcAD5L
3AbNwz3Sod36oi+hfaBpIjVPkjXppalsf8cS9VInxjPBWmo4MfHQP12137gTgCFa
G8M8h5ixDNyYPrPARgnEP9SLNJEM7WrO9w5h9CBX8bBH/HpyUCml+YeyJbYPS2j9
iLy6UPuYzMZjsSBuxSF/LkZgmUfdzq/cGb0aA3FzzVbTiKrcb6Mq1qPzX0A0W+8g
5C6va487jazTEQbtfV8yr2+tPZnMyIjom0HYj68PNs9zEJgvNENQ2BaOekyvcjJS
CAe8IPTqBXmVSMLVBdOY1lpwyrvEwZKUCVlcrgVJk1cMwLWS/10XQZFYk6CyjzzJ
Obp7dHVMZmV2OyxUtVumhZIWqyqP89t0h0hT6PjUpRn+liFpe1hUD0+f4ozF+WBH
sB06EnPUBWD/rbJMyUMEIBgRztmCdZdM3T3vue73Fdl9BDRRp6d37ahvCPt3bVdU
DnhQcfflBJxfHFkwsd7Q6ASIzGbT2xM84RbHrD5rmoCSdjQ2GLvNAEucaa2JdoW9
rEamY7JrEGi/v8qWpaUgWywZXU+KUOzrhOHP+5iaAukA/7YegCLFDS8JuYmo8Wtp
kXOFRCiBkSvokJaV3LGy7ENSZJ3ZjHDDQCtt2Mv12YbSJghDndl/mJ7gsamhsFpg
CkLhMtCBHskSH4IA9HCqJSFiVsHfCci1JDWtX1gwAiAio9ZAVC/oVlPc3rvsDh5I
aWHVwqkWdUWtPNguRlvTUcdcNBuDTEzPjjTvI5OLZ36SnKAy8du8cofwGzXFVROY
9LC+Qb9PeWeoyjnwljvsoR9mkuH9jPRGAmeAkHQgbXJU6YV4U2e4XXndzJsk/8Xc
SE8h35gY1cJf5Yb6K9J93HWTNOzBrLsV2pKorG7KEfuO0NJMWWIqfc+Gm9z1FvUA
igD3/tXbRGsWYonYtmtPRZz5TPWpzUHkCSUNSa90dsy3UhWZyYDLKHVkoM3618p6
urw38fqEcf+ONsggejh93LDasViPuquBu+ah3DOiediZ4gaNu+IxTtnGNbPCyw1K
GkCN314ABr/0aGPi5NqeUzO43rd6kr9L0JRnULd9TzeoLYQlPGPeXcwMAV3Q+qFu
HtctByR6x0BZw/UjBwPCX+nFs+cYKAG/xcZS78Di5xrhU5FuEqZfc0PMeG84TOzl
hYs7Sbp3HRTIA6oz19bZzpI5p4QYiPI+qE1b9r790ssFFXeHSRqK9oQenAuMJhN+
JmaJfyleiM/CuBp502KQ95HCwZDZTg0bGHlsigv4mWnugdAEbRHNT82pqtqk0+lQ
NNi5eE5bw/cWe7QxLTez1d4HsYgmuDeqrOOV842mmbr4Vb7v8hQv9BA+B7FGTA7H
akce0t35s2wMqrhsVTRBuqv5VAdkLw7jsys8xr6lwSeTK7gdw71tFyIzS8rOrx8y
9/VKMLfzMK+WD+GiJoxx3YCrQNGtO8SaVfIcYz9W0cEV9pZ001X2DiwzMpzSxhk3
WU3LyvXKsag+0HHjzPfhwESKMOuknrgsY781habloq/CAfBpSy/4dkPrCtntYDZ+
G8NihRn17TcJKlSQqgu1bP4mEQ5MwEWA0q0OacKFFLreGkRQfhgsapz0ebZM+SCp
mBpCSJcCLImio5oZIfwdi4TcezAT4c1k8UnBI2vI9bh3Xhupfkq6kF7WU6teOh1L
GBqknmhIgMbOPR3HFCLsx4/Km3mB+O9IxCsCzr2AGCN0CnyEkgXdzsP6ulfq4L99
ZJmSGTLvFumDCfO2EfozB1PL+1S7ndIkx8Q9e8AXE61yN6lFVKn3L8TXchR+9Dl3
W7FVH7YzkSOM9Wk+GmrU4BmIIDKnE5+/HSzKXojjtNKRGR9iBJbkdUQWo3WUEjgg
eeLgNCIW+qpLImW0ivTpVvZGnGjzpGE1sG0qpNT61PVH1/8bygTvzhMYJ6+k+cTS
PEuiesl1FMProaQnC0QoHVmYH8tDPujuaHCCcDZrwoUzmNreLLbDjcflCPY9OcEN
lY07P9qo3aX0bD+bV2pjS/I24sG8d8myxn8mxwDH7OVmU5XbG3PbXk6EHjog/ENi
Oo1GW2Wdvl0HfzTIUMmy/RCuuRz9fVqLIvrAZZUqp5/D2yymzmvp6rJ+rEjjWQ93
tZi4TAQd1nJXaAfNMljyCYnufX8qXxCdZkgl3KvAusuWoYsxnxJ+XhPlEv/8FMXC
6Fi9aDvgz1qz18+jyAYeg731Dt98hsBOVe/qeRs0mvvt5aVkInSSC8HxUha3xvnu
mY1fYzkrfyBIUiszaCtQCpUeG8AoXLsuBhl/YExOqhC5pNBiQRRkRhA+iK6lomff
9YTl2zR2gUSjmXpD74hqqMHhdpK/Dqd70NYPevYH1pizBXAt7zXKdL0WcISkLSmK
I0PDPKq/w3kPxFC/Z5NqRtnHr3ITFLgQWyWJMRVmRpbaJXco7dZDPca999s9gWlJ
G2oouRumB+pDxkfZX7Vzm7/69chEHbgW+2oA1hdiccNr+cLPIG9ms44kJR6eFYk+
cXMVuDKFm6dp6DhsY50mu/gE9R0YrqPK7c6ufNdotnuS4q+2/KaYh3773PaF6ECd
/6lIXvbEwZJmYMp7cvkNl5Ff1daxYP26ZLGaJwXvu+KFMApXC4HgSldBdiVWpdEH
fXZkslDoNJ0PaXR93tsaQRGO9kaezB+ViAG14wu1mOXW08NS3ba/fGxN4VnWs8GM
7Ouwoll/YxEdDMAAYw8kutEcwbAHKPpO1SQerhmBZRiP2r+py+TAJCZjIyrMc2+M
kIBaVgpZ+aPX77wo5Uq9H+xyqtu5kq32v/d4zTapH8HpVZk8YbCG5NG+8hoX3Ft5
dTvdELohdgj0A7AeWhfMZ/esI80ND6MpgOfphAZ5gTxjpgEg00CmF157ux2pfB0Q
YtpRGVg1jLxDnJWISBaXPL3zaDo5UcgvOSSqd2/zpNn/Uu54eU9kdJrSE2+Erlal
iJ4wfmzEQ/6D1pIA0SSDWOIl0y/JK4UaTwoANF3vp4qlAn9cxBuhj+wpdq3uj0SW
DvuROS/XeQq+koRJC3dPXok8ot65ptZbTbbXteeYkxe0DOyjFU377cAWfNz6n1vu
0bKbqdEM9mO4ANt4vizxNj2sdWb8boG3aZDTWBisIsEmwlYITrCtmX3cFtV7HOaO
M/V1COP8szb0xCFAacWgWhgnNJ6/hNyfPrEPHCZGaBa8ZHBevJLSRu45dDcus/c5
fljmNzi9y0phK83qN+T+QQQNBjBribNVjZEc+C8UASYSuKhNTSmeRSm+tV7k1tJh
aDIQpjocC1Z+IFJLmiSYNhDrG1uqgV8TehNv8Zk6GGUc5KVOdsItumE1ZLuyRiYs
KXADGd+PRRRrqyKP8BBsKV1v4CmDfWymAiqfuq8wFwQaHWqZn6i5gkEfXaN+usor
qN9bmLYGvIp5+X+adPdb/6MIiAwwCR+EO4oXdLsWGe3CJRIjhnjgmvkBSj31CL38
VE+A0wx9CrvBQwkS/XOIu9n7+58TBx83JTObsRYnhhzLxXRj11HPwBCFQHRtges2
uIpDDBSFe0+bVFJNkUovbPzNsWBTyNKGjLNtg7X2aELajUfPZiMj3HzYlIl8Aqes
Rkud8Rl+FaL7ydLSvhTbF0u//6KI9w7RzcWLXlCleJgA7g10d5TpKsS9suL7xc9b
tZE90SB0oa/cMYqKMm2N/hJOv622UX7ltGxKuBzEPOgOg27vUkKes/u/DMi/i9b7
V1tMxmTsW4Z4sDEgbmWv/7hHsx+S9KgEry4kOXWuc7suGnVnjAjvIJUyNYWWqCYi
solq4z1SrTWyQ/oaHK1JAlWVlRIrtAdvWttX/t10dZW3q2Bj0uItrOsK5xz0hdhp
XqcOLinHXOuSXq5Vhx5nGCiL+XZtIom8zsm1jJDX8iYYSzkROPsa9Iynl51XjF+j
bzmc37gIdHh3Z18WDRydzuIbSPMMANEUWrkW9+szWtdHK3jwzfcem7uELBSGMsAz
9Ly11sXd1abzq9ZA0gAIo20oX1mGDW2OnsnYOigCyv+lKQqYNBSRWiZQ11vnOfD1
PpGCmmy/r2guYplwQLOhUpVk/k7UMJRZqTfFcJftv6qqb3OdBHiekXV3qvTrjrfy
vBww3sz53RLWou3tQ+beB4W2Cizx+h7hBpplqH6mWGStTbX7gMaWC0O9LnUiEHqF
NS6+rmc7E023WnzRqRG3A30P1o3ayb0/Nho/E+BgATSxrkPw1VGXgaO06JK+6/ae
nOBhfGHs3/6CyJE3nxlnrP1cHBRRCvMzyJlS6Glu2jqa8fE8RLwf3wpNpN0R6RBB
v5e6sjMUhlngjLgoQk+hytBDmmYtVWm2oihzcvcTH0Fo9BNb7IDPnPs6Kk4avwEf
ovtKpf2PAIKLtbIv581A7h82AQoKyVIfKqx2iopmyHf8iFplABK+IWEk5grg9/jA
faJQGAnIvokRnIG/gDzlAmud7z5Vy5yf0lT0o2YT03jY+ZUK57RUfN1p6ySgWmi1
Nk0Hkzu9iRYSktMgXq1yoGyo8+po32uyEjIRvt7KpIEOVLlXRiAT0IVimbOCqbjL
fRPYoGVQUnU22/8VUc2LDmBl4uEqkrtAc7rKGbFxHXZO1CUUD8afT9UmrOPCV8bb
0HIqCXAYZOd65pfFoy40WrwZKjkNJ/BoNOpY6enCR2oMwns23lE2LhLJyjclUzUE
Cz8i6VyaI51P94tekB+BtU4K4MHjgqKGXYViznb2bdi1G8k4yGMfnI5F78NdhxK8
AMQSEF57MjLEfzkzrqJIcHu1UilF0RUffqUob3HRb0l5jqEdZlJCEv9uT3oV0IKK
//DkvC7LrX8XclSzY5REANyjNoN8HWAcsDsSVmf319dXhIeSp+LRn72f5Ipn0kyl
pb4wPuJrR14zluOjrcNwJdn+7oL1e2n2vszfWuYz55JnglhhFiPAeo/+GWrjDf8I
fnCr51IV/jcFFAf4GKgRBlKaWgeZwbXdSu2m0zntesF7bhgTWNWsr7Zs+XMaK0/E
vkaA4qqFBLE/atA+sBzufFENfMTyt9ehLXhKjSXKSVUaKMIYqH9kWGRa3cy84X64
q82ZhXsQaqhXWewUskUoGY/4pHxSTT5jkm6arztIZ84C3h1nsMcSHvmF6ODfWQtS
ziERToB3Si72dTYB7FZY5sItcU0e0UWqiN/dyCURITRK9RJgmSZ4PSsKIkPCu+MB
imbo4wtUJ5n1/1EMGwANZfndEZ2/HnUiSf+J3Ouc7gRkel4EOR9MR/yyPdMs4kca
sTXQjHNrhtbgMg7AYkmUZntZ9nU70puyQY9CytBgjd10Wpz4XVgF0LIhsmiJNPqe
liIngCVyHeqdPyx+tsvj94o/Scrf7EYr1CaT+9mvrLnsK1cMEWxZ9tMkHEXco/PE
ISs7TnuFzm1gYSURGSpNeLuf/r+L5dhNZQiVwaNBGl2eD/yKcUGTrE5YlGCOxZUv
6yoh+sr9BMHH7L5lpLj+pgYv8j4ifJ1Q2tezRnYSvJx8xsbgOuwhvikD69xhsPPZ
Cd4YjjuH3y3ymBKdEJ0TXKhUrWKgRy+pFgyHp3/fQIV0GH/t31aMsO/6enZvbFiE
l/CyAZ4+b3E2DBc51dJNbvILTye3iSleBySGAP62ZimoyTGijPoed4wxY7QoDnTs
S8sbhu8naArahlpozf5xZXE8pW3EoO2vdmOrAzitMe4mlzh/5eoJWbGAfvkELaKi
RgbBG749DDsauiMNWTLW0xSzTB49XVoC6gjpGOHJHWwkEj5ZBUSJj+si8Xleb7Ow
fKM0YcwYcj7qVNPo1+nk3kgND+3+/YE7IooN8c92PQEOIGlZ2QGXAO8zneeDFE8b
xfj2KydwuENMaNEAeyO9NihKOkeBF1Ck/50EJjxFQZ/hzsj9+mQ1vZ2TUNtRNJTN
ZDnph4su59kxcyAWKnkiJr16UVKxK6SsjTEU14xMl/x4h3ITIF9ukO7rDWEFerse
yEu0HhbVHcmQF21kMGeXf7N7PDC3z35eamJkQSz5kJD/+CU9fPgfTwJAv1TNfTDn
Baer4bM2IRasO/CiXxQ+mDFM+ue6Cf2bE5QoukNJITJD32MVooY/ZBHcl88HN0Wh
osfnmbWYw4wGXs8cfh4H9AcfmT5MNp6rYm7RjIweXslDtBLG/WL4NfTzOMdzgzla
4lT7nXaRrgi+x7uA0PbmKCeU7i6d7dRDdeumXnvdpE8so/1h9MuCyT+sPr9XkiAy
tGt9O2yBRqIJykV8CUTg3hQvAUIM/JgxqWemKK9+cFDkOHqbp6BGzzs4/o7YnCdY
mNlq7pLKMeqvspBA3nWdikSFYVBxK+WFg9RFjn3bKRGhQoFhgMpcYvKUCpRPa4I1
yjxo1VSv++gNKDH+JNYpaf45NyN0EhSsZ8tLyVhslNM9M5neAmiDygam74UwciM+
fPwruZMexLZlQZvoPlJ85YNuHRHENTHKuoRdFfS/XYRw4dEY/fD4tnwvN5nHoQoX
cZOBckhGqavnQ34lPFB4pdocSoB25XqAc2Zg5ATgluZzHGu0lKEPjfVgO3HxwXhu
liiQYTrM/S49juMOpUA2Jtypf3YgYeoCPudpSeFGclgtUu3/AuPpmrXIbEiIjQs+
DM1WHNytTIBgYLf9WViU65hdrpAc4VmeurX05U5wJS8fTn+qucfJCoDtvn7P5NtG
J+5MxQZjLtZ2cMP3Gd9dxG717rv9zKcW8MWKFHNgQAQScZ19mciqOSiA8Z+4P/+0
DDdLl7zhn9K7vhXCR6FR4UBObHo4+9xxS5wAi93uZFkEFZRNwzwvhclpN5J8zK+F
hqCaDckWezf//L3cXeOvssf56Y4vQ7s9eS9FveXUtOod8QTCgMifJRVSizu3TC29
iskcOvTjGytMfSKCXzrmwiz8EUaGeKkxqbpDTF9GCbOdO2cUR0Efz2zPz0DJz6It
zCqyRCdeaNdh65rfPw9drfLgakQhgMR0kmIWc+l5SO8HgB54dJdPQcmtN9TbSTba
j7eXMUcjCCo8yWMel2spGNBiWigbVIgEyVpcE50jZ5JUtMlrE4DzSPIzE5ZCyHYX
QLZOSDAi+rrf/vTGPym2n03g6lQzXv5KbtaPVYfIHDCelEeQwyfHYws0DOUartmr
Hmhgf9A7g909OFULIxYmQs9EBOk+g0jnSw4KtYW508QMf/dBZdn265bOaTNf6wi4
yUTWH2ujiI+lJmqrCM4VmGkBZm/T83la+EGU1siRWF2IgHsVhS2ak/sZhscHr/Hl
BHMK3U3VSZtfbTnfhbp6gMmcRpcTkMTPR6sAMaZ9CDmuZip2bMGpi2p9rEDwWfcY
E28ornYcYyzZvaqGHPMSphXGFvk45PKZA5NUivjuNdke7pZynLfXCNhAeZDYikdg
j+u6UfNgETOm1nl7eiINidb07sP8kzv/1LPpOswPvq4Qe7CwIaXO/CKXODRb+nZJ
vg3XD60yIFNsvzh78MyFXXpiWUv82H6oFkCubFWi4ZH3M7PFqu4iYzDg39JSfAMY
UON5jm8sXdUz9Wg0i//mQM6WuFPvcE3vPEUWf2PrwiawgbSdAt8pGC5DoBAnW+0j
/9259G4rrgGhE9H3q4y699tX0FfHBcQIIpjyQp/98eI2X89oo7yPOlAlW4MtoiJu
nlobb14sA5jFTnPTVSmuVepT950N2TGDjamZLTf+I88TIMIIPpRpRuQFtM+urkkS
Pu4lrvx35xY2gtBEDLZOrMX2kbURBp9QFrm081syQ/cShTEj/0RsWGgMMYYmnylp
IUubbl59+vXHp9Tpn2rPwfIHcxnSlLR1kSyo3K1PhHe5dM/A4xmL6hctqbnnYbdo
aVdKkvQLfzPVCLszRkgaIVnJf+AoCHGvSj6YyWKs0aZzimsKilOwvgluL769/ig9
kjMyg9wY5Gr5sA8LqZxOqVgdmyTySrMsWTJu9dRTo8w41p+ew1FgKWv1mhHBFP7Z
c8v1LodFGphzx2czUlFbEJfakDRw/KckkmrO3ndkdgEV2iQLbiq91UC7zxEgdMTI
IKMUdyUScGOT4SbIAfDySCK8QoBsfqrWrkgqddBLXuMOZ78i6t3Pudw91tJz6/wR
p4u5vCa/LOrh+ajQXCwfug9e766BCIg8mLTMCxRn72RcVzJc1+hreM+BJIQpkT2p
RE2qmnQLxqZFG5BhxQVixg3QY3DE5ZHIE/sk8gZeHT9rU5/nMH5bemBsnAh/w6it
JKJlCOo8TB1tOW3YaxJqqiUI/H8gWxmNfQ/Qu4ubPfZwdOENVEF3xrKCjgja9xEp
H6mBjGEO/WXWI4Zm1RmJR0rl9lMQcQpWxXBTeoqfCCNHlO3PnxgpElKy/wPpX89g
1V4bUfOgr0PwquyBVEcDM5O/jaTRL+ko70doRy+wxiWqBT6PyoiEuMcKXH1sd5Lx
aUNVsyM3Wpt9jhqoz1/MAw3k4miO0x13Luy4b7kbgELsZUrOLSn+IzRG7cVHPtDu
eNFiUMjp3jgktz5j0R5VeQy9LvUIPzAN2txnkpO7M+tdEzVPSL1ZZylK2C5o67FL
2xK0eUNk0/7cn0mCOyGIBPAsZdVTeqG/3I/3zrVu4KVRw8Rodkp1wkXRDIULvxMo
uaUVGq5015UODEwLRDpFieoaBQ/Sq6e4uKEoAV/wZi/7B0D3D1FwwHw0CuV1aPH8
fWlUvBpMOBk2bO50H15n9KSvIkfLp1PRcHR0dSRnpwNGs+3sIzf6Ht+YNvrstpy0
YQkcZ4cD6tteTMkJYCIgm5AvT2LFvJMFFm2G0JDeiXTlYiJRzoIoTpmlTceMRFiG
6YOgqtisIvxi2VGVVF80krG8grsib8oKzjOZByX6EdIXR5Mtle+DiBKH1r+kKBv8
SU+VEmAJ9wZySAW9mrQjnTeDy632ISHVNE6nperWvmF1z7ostbHn8DQTmhPA7+wv
phDzHn7LIF2/p6x8VKCWjB/uvKeAlldibaUmIq/MmIIEIeaJ7FC92O6LtbDO+pqt
o/hQM9YDWK4h05HW79XCcMXXHvKHuWosDCM0gjfMQlDUOT0MZoxfBYNThd/+OlYA
t/YINytve4dkAqGnQDfMY0CFc3lAFugWBX9ye/ZoZ4cMzCesaegFmzwJYd2qN7YK
rpH8dRNSQxk6u0qWqBfEV8Ni0fXS+Le9w9kS3Z99LdIsiuzb0dT6eQ5RfEnWUbAU
ZTzuh7qqJ90L57elzeJyalcnUm9gCR1av3M19O9pPqUN1L3TpIJHUdspAF5o22zD
PwHxuB2G9jNFw9KFvY4huMXQf8bd7K4AaptAO3vRDB6g43uCE4WVPHDeXPJDPMxR
UhbylqpT52LqITSetlF/aOlp7OCbslUERlToSQIrSBoPuQBlp5TRRyOOcKP/+Xsb
qH5Qv9deT+/qF4V8tDszvHnlgqnPiKnwmR5QF02neSZY6E+FWeVknKxDl5rQjMFw
gF2ccpnfCKqX48uNRfOO9luZJaTFNau7umtxk2l2vdbHsGSnlsFu6VlTZHgjeaEj
p6o/Z7hBS99qabPPLnVbMrLsTMs4LHOi8GFSi+llfdJAseitTCx/ES59fNjKq3FR
OFN66kI2qPkE3teJ8e1h2AQSfwXc9NN5Ynxkf9vNrdMg+z/Dd7AmRpAHtxKvqWmx
VaFL0jokfAKOXscP/S1ZtzrtrFmnr0snrBvT9JWCtLQ11f2DOkeDeu/jXw09Lvhf
frdz6CXtX13xxWl2mzpt35PqawUMdPsCjkKrF+Jz10wX44f4WnsLmdRXBN4rKA/y
1U+48aVho9O80vPzHl3aJSoMAIL07E9ebO/I10bOF39fxz+C7Frlw2/GB+WhGAYx
+SnNCAewPZxtsokvbITtXj1qbcERUn5zPO+bDOrWWr2PtOkzGzJqtBuJgZizx4MD
mLA4BBIbCLXMnli3Jdy3RIZ4POKEMJ1QLzPqZVjA3bu4bWmPIC3zd1JaQON3fLfI
LF/XgHOM9AbMXOjC1UM6IXuKL6ptvARH6fyFNfHRC26qJ1/l1RKEwjtcLctXdB2i
RflZWSRv0CXZj5IgNvi74cfcA9HZDkSXSSnJcEG9+aDGg+RKcbN3BYhYbyP2iNfn
Il+7M/stn7ow1ZVa0cthRSf1bM4fsNkFmvDV0yHyc2E5GQX35f+0qcgF4GkmseXc
G1qWO3WpY4WSjLDANSmoEe8tUGjuyKW81YQDlOqizT6vpqQjfgnVR6M9QsaklR56
r1NuMpzI1lGE8JVOX/RRSwXkQ8fC+YzYWkqAowgHF9/BvH+XRbEi/yTTajIe/s3P
KJE3QzEOUpyYtZk/8gA3e/txU3yia7OqfO8Q3cc5ltQ2frDv7J9//6vdAbvBIpmo
39ZaUpLoER/tU6gnMEGwE9/PHfPSHKaYP+Dzk2bxmU+A1QefnBi0IWSqWDHkjZn+
tfTz3CtOjc8Q6KS/dCCfyBPbEzeB4qCe6tETj8sR5FoCuL1ShIYv/vTi7jw5wsYP
6aZ+V2fGG+Ti836t8HEd53KMXbOb8JBtJUCiVdRqxQ0m2Tt9gLZbyIa2ylaAyOJw
/lmGCjw+Co54CoJe/oo7o8KLp/t750cRKDstCD0wtrLy5RhEBdEcwOQF+Cij9M+s
AwbTw+PAh+cEyaHExCCqYqbF0gMApFKz560c25tOMO98eJnBcQW2lxkfFH6Y21k2
Bjg6pn3FHRqj2HeB8XCcCdfFouZUPlR/8tC5T5LyoteNduLVEuu3rcqsiNPDajAb
S25PEik319l83i+BnrZqdeta/EUFNn4VIbR86jxjf0aKsm4ZoJwtXDkatI7wZI7r
7gls4qP81bv4k6kUgn8DDqtqRp0S1cbcD7mxy2qOhf3Ifzxwg0jxQV8Nbsxfsqnx
jt1Dsuaanlesf8KqIrAaJsTT9zTMhmGJAxaAScQiwIEXvxhZwjZe71FJ/8Bm6s3F
2PNIoiEOQ3KdXVjbhjOWBFWDVHazW0gQHCbuBJKWJenNCF7x3divKbCltsavV4Po
1bcUKz4sEvMpXClJKiWYswcT/7G0bECzTkvJ8lhaoxXJdfhdZBoJAc8twme5i0nM
bBEbmSGOsByihdL9ZcMajOXub7FcCDnfzSnaLA7pF/Zf9ovfL+qD7IUt0t6npIzX
k4rjyoHIXSKNi7TeJl2nPzrHihJ6v6/5iO+AUrPG4CU8Cial+shKMRYT3q5+9c7A
Ve3UWMFjTY33xbqAMEo0XBQjMlMnXES0OdPo+386kBK8YtpL89kQsonvzkGo9ded
pm/KV1sQGc7QtBSR043eCzOPbruOP4m3Iuf0y6PZZFiNwkm8zBwls7D98w5ih6dy
+Z52OrWIEZJKGyb4YNt3XMDV42IY6YXBrW4fNL4Wgzc4/WHHbfAdewnQEv0VNFh6
bKj1ZrvXnR/eDJkYECU2jsD+HlAMBYfyurZnacnT+6rQGNTQdFg/bVp2nXrbUXcy
rA6VU9lxPif+Yv8NU1p6t+zxrcaZneZfoRwXZiv6q3DvOQANcjmNXbvSXm0F6DSD
FzE2JA7IUPZnwKwCim9oYTx9KQtGKBiZpKm6dtPsQYb8mVPKuhQD/DnEWkJnytW6
EbT32gXkOheAZIs7Xlk3Cet2++Qcr4zrnv8DT81tBH6Tq0XOrQR2qrVpo0b/CG43
42IkJm1pvURZijZH7lRM6AuvrkFAcFpIOx5MZTYgrrpw124tDXpakg6Xwuvb/Db1
UEsOP7vwYoILALWE9h9XdoAHwFeVsck6Ha9PiCWur7udRLhDmOuFhHSb3UjsGRFO
yanN9mnAAjzk/AwcoRDFUHy8VrFpZ57le20PYx597R56Jcr2xX29Ofim/sb3pybl
J40m41egygC6XB3h/EFG3Tc5vrJ9/h+u0POCfqqwO8k5x5PzzhRun+mNX9LHwPO0
DCC69RiPi8giFGadGYDUAinkHTZ39rImVx290vjO6x1FO3lbdZ8auZV8pog2j0iX
z9xq2oU4aIhJpl7V6ZdsegKfXajLjjFhkfizW/M27i/inqeIWIpFxeG40dSAq4n8
ngh9xat/apd2KIsyMJr9O/GG4Xze0evJPNObXD+GLuBcudvgiYdGXxwTmJ5noTQZ
Q5GQpQlPuvOJ/3QUAdLEij0K34wZAGzsn3j7alGqOmIB7FpDRhAoOB0FKqKVTrMn
F6BuofMy3/+AANUZ3yVQhB0WYZpmDBCzJL8NZ1UIJx2t2mytM3mRfJwoiUTvtKQj
7StZzeNcE2TZG6WSwp5ZuJDt5AvwrKLIhmY35rnfsuUBs5ZZLkAkEmgwpCLDyM3R
ro7NurOJ6X5Ib4Mak85odGFFFsyG2cw1GdHRN1KdB1qaNqIqJ6UPT4PZ3hQ0p08O
uGTPIgeECuw+dPEcqLPmm36/ozMtpjdCvm8En57G4vkGxpezJxCQhb6crl0/xO0K
CAd+0o9YPLhwAy4Z67dWCKvMWSfuveXNnPh1OrB1jtOXN3dy9FAi8MQ65JeyrGUf
vZVMTT9Vv3JEONQJjFIFsbBHGBfIwac5EvSRKq/mhgyzTXzu7wXtyY9aciBYbuUa
XHl60Xsu9a7l9yMEc/EQLWEp+Tcf81GGXXUd1T85zd+7rTCVhDzBrbaODVMdAbBl
sIc2YCxZxYk7K6zKywLdIRvWbA+sfePTo7Z2ViTkN4dF8rHRh8tmnN9bh7FoY5AB
eS7RyQlffo6pz8u6J3d7LnXD9d58W37UeaPpO+RZqaXGK4zCfxwpCtOpTQZifkEH
dpwf3CjpErG2QHanFsyJlL0Nz0bwqZ9WZMN2vULIwc/fHj378XkfrS5xxpdRHUKX
7UoJKAIgmHDKPF48uBKSKQyavFfPFPXjEViSC3xo4JhCvIirLGhLk9aZUxyrQIJW
yvdgsw5nOU8mOhj4Seult7cBgIpkL4dy38eh5ZydV90QJFDSU+Ln80wZxoILqEUf
J6yuE5PMHJ0TWjLtss4OyuY9xbie2b1mjcOFcREj3xCFpnq50ZyGzDf5QfAKCN10
lEmn1USjj2Arm2KuHQF3g2Bw6JAoEV4lfZzVkxhZPA7YHraKuxj9JaIUMGmVHZY2
BOZk5lGPHuEp8tK5YIVdwmBc6JSgUjOn92NtsBW4hFx3ZMKTaQMLTD6FORWyGlnk
UHt0cWS3C4/fx8RdPCy/WZL1iUzBMJHNBL+XjasP1VEFt+5F/usQuWgOV0tqm0uL
G1eJhBQGHbckWa7GwlLBiDSEdgxsdz9ifdsL5mVTDLp9zJUm9FiS9MsLQ14zaXvn
u3XBJBlXDP0tZwe+r7eQD8YEBuO5Vs1E3CEmIGWlB3Mvzlh+TAAeDkchBROz61/J
Ry/QOIAt3r0i1afPVJNJdZDdj6pmcOo97bZ8Lu9gCiFvhaIKcHi7oflzw1Uvrh3a
ddpVSZxg9fZgNGK5vu84TdlIGcirWcYGGb55UoP5YPsRmxWhKuHIJeu6H39ST9fr
rl6neoq8ujH3fDRz3DMLuZhaF9Vhkdr7rt50sSvt18/5rUVadl6/UMOAS0by60aS
pFA3mTLQ+AAmi33yRFJq1g6x7EmuOQLtmaq1cgv1gL7WPxL5OaQxDIZTB4XlA2XA
Bum4iykwOPg0Fk5Tunp+JSzT9peZEC1ZkQrH0X+oZ1pZwzWxytwuUvU4M76WIFMF
j/SjuH6Ksw9QBq+7uPfrfSy9CXqh7DhAW3Uy/Kwuwrun9NffcnkexldbOMFb0Cx9
2+tWVM+RYyp2KRIOFI1tZUBYjF/BcwrpFsRVq8n98QhGT3gYUYfmgjw8q/qV39dn
MOk5WIX+8qa1IGF8YM94QI2cVavBUb2IVie0eZdeaGLr96eJV05rcs4HADwqf16B
6VcAcFfx20RU6oC+C9EJ0ir8D1EElIDRd7oo2d5aEg/Lj5LXdao3M2HQdM1UEQt9
yF5S/yvfeiqD9Fdv+CP/eVZmkowCQp+F8zPb025gH9f2fN2uJa9OHJYndJNtsrgW
2r8IE6IrtrXe15clrD3nhxoyvRaaG3eJw5JwoGEeHhFkji0vHmjWNYHax+re/43h
7SraMS+L651+mwSp1PQIWKQfR7JkAWfi9PV1oeNQew9+wUEe2Q1eCYvFt0S8ROHI
3COb5tAgjXmd3hiX9LIp0kSZJrncdOQBfLxfLXRuquwyyd5oB2plLxowaPtF8jD9
HoYlh5JDwYGzmFva/TUJbCnOiK1qbFoSzkMc0sXu1tlzO9kph1JKDZgKOcYQ79nr
sKCH0QojLOiJuPhGIJWeXVYlBiyBLLc9V7GYw6eDvUPSAqncWKGbNdNDYjh/glDl
VKW5OyPBv73FBnsVjXVZ0nznF6H9aXYGBFcKtd/TGJbaXb1rULJh3Cbcm/NVhDfH
LReaSxYv/+4DhfvkXneGCCBeLsqpUmKbHZYSOdsITG4KaVKK8cx3elYcTfmShZWG
S5USrXDXBZWRCp3pa3WsxcPAiNKm1x5jSLe+VX+Xf6K3A3BUlRLMbNn6PvkzkA6g
V6P4jElG3zqoMiF0C7XG0B0sPI+XjNn75KSG6ccPUOI+3N2OhT/qQHlM42cx8LuC
59mLdUehirf92DeUW2o/Gi9W4DBuBFmwM22as6zap2UMm8LyHCwzMoI6mkBlWB0V
pwKlNVEiC1UfPHVU74MCkMqFrR73sRlmvVin6bGhwlh8t/9AKfS4FUlUEMBJjRGV
7K/M+1NwyHPbOtRKkUSpHJqJWvIN2H3ZsFqCfbalq/pczaEgXFtHX30/4J+5TamG
M5zHGfbWt9F4IznPm3Ez+Z+wj03eQrzWQAEAvdHFIU/FKzEjaIScziEPWn1jN5zt
VFaN9NBs2/ss3w3qRIS24OJK3zbA2iHKx2nKeXF8vndN4j4vjS0tcoZeRZ/v7+GZ
WdxMbLrupVYnaZiy9/aIczwbBnCK844hnvpJMRhwP92WCRGH6zUkCPmfCbkPXHsX
g+Nq2rTGlfxDTaEVGZfmzZyITme625HNSHcOultCuEfz2Q35dEOpUUCQ3xcyJApa
wJTxRCo86Vk2efTm0hNRCHG91eB9yhgujGpEx7kb0bRpEKBQdZwW8Lnbnqz9Dfiz
zNVBzhQzeCMFAngxJiB3RDdW8uJH8vZAHd4jaNBsbv7joOItisPv0uVPY9I8ljQG
nLW4TTP73Dfvwj42aB1JcF6SR7F0Zk8PqpyRO37M08p3etJ61LSeKbayIIyIbYId
wWfDiz55ERV8usJXP769icqRYedEMObSFpqf/kmDQr2M9SyY54Koq6NWeZADsl6U
sfurtrLD4iPEKFko1A0iM/aYj6WvBJmg3A1Xye2+jO+4qqcLEvF2X/WVM8SwxjfC
hbM4PEwTyRoMMU+nwNZqhNQgbxdUktxtCGLfdDisSoM6F9AGVC3Q2ajmTGpVEJh7
QJ0tTATHnD3oxM5aUWKtCYgVy8XH+8Ht0k/+mHpbAi2kdNdzae1qJNNBi9fEBax+
k2fBwgYeUSUnflfAK0BSpIdpOVOtV7BI6GPkjwNj2wkOaAb64wWwrWmslXTpkr8n
QrtjlMWCU+qr65Km64/raN2IGa4sLK238iUox0b++rZQFIvq4jo36fV7RDmnY5Of
76PQEcEOuXLugKF8YFPIswAG/e23woaiNlNxrYCPrdoRiecZMfe6ulI6Fl6ovYSn
P6vnlNc8FR4pMH/+W5Li9qntMrGMM3w4g0GI3Cac7s+9utcVCUXtocpTzO6oI6Aq
xO8gKyv7KXUXyN6f3hIg7cVxQbbMQuZgYMGp3q6y0v/x8/750TImv8YYcQKy/yKr
WhLcyKpcPDUrj4bt4k59KEFFj9VzBgloH9uqALuGSe3Cr6l34Bbw9IieGt7OFjrP
eNIyS27l+zyKAyjEks4+Js6QzHSIKMjY2mMzpWKU8X7tYsz1vy2efLpVaEaxSu7V
aitxyl4oseksWpML6Cvn16lXkpHsULNJ2U+bNETp9Md3JL06EcEMAiswp71JUEUQ
IyxSBQIib3niaqvlDgbEeVObyAL4/Qpw7IcjaDKOiVRu4ytf3gSUwHn5ffCqyOJ9
Wb9b8p0AxJcJatX7gJgok33WY2ZW0HENKi1YQv6avH9THsXZDKmkXh9InYTaeCmR
vQuDnZgMhegvWRvZJz1iBjlgr9tkuy9uZnaqt+WKTQy+uevG0gRw+Fb25mGu9kjS
FwWq2TuIxZ5iQacVSFS8wgvJlprPZuSEB6gMjdHfjjwqlM5+PiOUS7L7siRXghgo
0sg4YZXAR4ABlf1NMldv/gYHF+V0Ear57A3IIOuWNk1V1ujmw9OucFkkA+eE7P1F
aW6RRrafk7kz3JmBfFwNcytWp7hjRI7XWJsSb870yUhd52uSMwocxUWvptRcc2CY
RTVYhIF+gG37LrNppobeIehiyDQm/df2mu/aD3fPdVUIiLTyFMhFZVNoyllj27ih
+aTBviuC2gElJ+zvUkVy8hMYb4r3ha1phqdcJYHEwV6ZVqljFtkU1fuKur7Q9DdC
IEonrPxB5GHRzsB5N0MclN2AbaZx+B6+RJaOVkFLpnF2I0cy28BqDk0/4C/BjhaB
VJA8ohO0RfqL45fD7yWyNWFAVKeMVb/ZAVwdSbu/QO7fyp27Saj3Bk1vYoWZIWBp
Bbb8alpvaudm0TvT1awBqWAYOHuAG/QKovuRe4FNnBTVnK7Fr+e77PI/Qvf7VQgk
neNgHyD6Ne0D1zoT800uYYOHzp75OLVmZkHlHsXvPKlegGQ6S7UFNoudxT+YNToC
8XwS569/x/6gjgwoxaqXAjr34hetegnUuxJNyTMFKMDGR/UEs3kJpHHYR11gr0Tu
cgKoE2HEh1Xsp0Bd4iS2WxqmelichtYcci7ijtdqtllD1HJg59hPr1BYGr24Mv50
j56fzw6269vk1ci6euuMnuXsuZgPivSRITJOE6NmqJVkQxMBIbiL2Xorl8IAH02U
Eo3/5nCorcsB67hJtJt+YE7lKS5NsTnoU7jvTCDzPFyGUAaIL7n59UjrQYiKR2Tk
h+PlDtnSScGm+0LcGcPewYKRA7h7PEPBHaD7QyFHXk/o46cvYFpnG2Yse1Rx6XrR
GKzxT0UKbsH52aeBsqk3Z19Qmrd9dpqefo5TSYUOPCBcMjOMWvEjT/MqLR14Rv0y
6CjPwlc+mcgSeE9TM2tB7vrzVJ76Ddmg6mhHdyzUDKtb0q9t4/7MrwpUKG2LPB9s
PC5N5EFpEYF7ZeTWyim7oF8hME+BhC+CSoPLNCQcmPHXKlGtfoo4xQ7UmdaiYoGY
fGhkSfsev5aloodN3vrW6Tikvy59xogbT4U6UNX4Y9LPojZY+MSgvyyKkk/50R75
qaoRVywVq/pEfx8XS0NTdZEa0wEBu12SKWh1ABru6f9+vj/nxl1lyPkiVwrx3z8Z
W1110b7iQpo5W1MvsRFaGmmYyuf72kW/uH8zUmxe6Tnxg5I4OE0g0PfW2OmL+yMk
alLSCyy0SMb1QbimTL8o+S2f8zRCczN9Ior1/xjb7OURSIrAr2hEKw40HqkmnvPN
B1DbLJJMNdyV2uCuekz6Up4P70I4TzQKzJISrC2VZnI8dbpSZwqdEFJ9epgdjXmD
DVJl+mMNgRAIFjXiNOzYwnL+UQQ66Rur3Ui4qYLl+uGgF6k1keHE6hbYzLNLPMUZ
hM/rbDcHujB7dc+0DcDSKktMOU9fTCNJ8ElfaVLMA4PIY1LMiJsC8+vjRshTv1F9
4aVC8CwUZgoVscyS3+QllkN5dnFm2v/sUswzIJ1hE+YTO13rVFKrNaWD3emSq4+H
vSZaqlazLii/A7y+hzWvVYjslF8DnjTuXIoLaIvwd1e29EP8d5IZCVuxDfbdGaNo
4jOoxqQ7JEHcTbpLzFaPNZWQIjJed+H9zDVnkF66HM8bvma6ahdMelnqbgsGsdrT
aOEybep8a4XA7xt9dI4ng+g/rqdiFu/eomQw3yXj4o+ZgwxGR7YD5ZFRlH5JAo1/
6QXbKng/9gwAXcFEdi6jC2iOfyfKZT4nuv7/ZUGQKBt/3px5Mv5tNxbZs+hoCg++
QcCQqaM78DmLrVZ/IvXzlVcimBDnnw7TsgyubESGSWQGe5Gf5eANocpNdPlgODZ0
PrVtDCuxHtEXMXekMsiEXxXGj7XBwEMs5UJn367wU9KR02jFdu+JQW9yv0jJvjde
CelrfR4y8uds1+ihtq9fiu7zC4pbuxoh6SIN91sHdvofKXLCLxuBDxxft3rTFpBE
kEWfONv9Pm7LbRdXzAZ91zDkplgNLOO/vl0xxkDIZ1lXUyvXt1vjonh4kIDHFi5U
0LyRkhNfKCw+R90JB0H5RtSqEbLniGT36Fvo3oIv13Q9bHGlVS2sz2sbfr6Aqtwg
JJfdkxIm4ynquID5rCk/yp2iCSyc6ejB8XkQQFMbMGTB3a0RhhAND+aRoNOBb9BJ
405Ie059QAdzN9x/khFSpUGfZrffneesNNjnk15uWG5Sk+4cEwt8iGh4Caw9XmZC
vMECvYx9ZP1zoZM8CBlcBoVkrJ2UTWbNqGcMUzHSV7No62xRypK1gHpQjGFOa0re
QgEJv1vIUYupXpQVG5q5mNoJTFr/B8Z3TpQIhn809phZpRXjkTPPTjSMjWYZT0iR
lo+Fi6TogkEXSsIKlH8gYpCFBaIyrQJT/Cu5Y1H40DgkximxNjx8u9yF6eiSdRJW
X+n1FrgMlQtqIAOBbdDDkH4WMIRO6BGL3gorL/3vDGWJ06w1ZwyPMo3ddGPMV/Tp
/SNZTHWEGkGZaD+wOP/kQDTPteP73fVwzd2YvjI3ea/n7LfqDri/1VDn6mzg2K+N
2W4pYX9dJLv+hPPbRFlD9Qqapd2y5F77SZVCsH0A1gIt3e8yEh1F0OqDXt590SQl
qGO5r7zeXvHMkVPhjgKEohJ2kAARQl3TXR2waAFHsA0opGjelOkFOduDd6+p0GXE
zNzyaWUE1/3XeyRQJvc4feaLa0UN9UdlmfyBQjLM91ZpNEoRyuznA46XulrKQxXf
7DV9yZKaTua/0RoGqwBmRswP7kZgJzZCgjYqngJvBH/qWsdIBzO4RouSX/c5zLMG
v5hxSHJ8eWUTtRnv5N7VzitUkxr5JFmNGawyEcj3hJPLVPyJTguFmkniUBQ0/dvR
bRUyn7112Emzzo53dJFMibIARkPea3kuuCyEsNcj3gsfIs96da9LIwd5DcNSgNWN
UDO8BT6W2/bWHdqK1YYMh+7WKSgUqTZn3NLE7i8uNwsITWxfs8wjQlbvrVCMT0p6
fd5lS8uXfPOC0nu/WLvplSt8Derm81+y7bZFvxFzz/slGg4VNBQD5xqKbzgqY2xZ
Ht3TL1eikPQVNdnmq7mCLglrlppV3/c3RSa+RYWzmDMBjDqxD1hk2FLP5WKYnERN
TQ1TsecSH8JWkLin1QRsoGhVlBuHYnWNoDr9UrUMmcoTtUlLQz8rAYfW+Um8afpa
GU2WSUp5du6+pqyobO6KFMS7VxdO0esATgNvQViU/tdwhK77dJxwdJXhvazI4BJp
H8Qbi2XZEsGjMGW99YqjMsJob24XWLteCa1cusR2ASGzQlFA98TyZJatvYiOY02N
muZOS7JyTWwgR/5tNHhtoaTtTrI6I4+R/4wgMxAngdTqj/FchTmesJKY+60PaFpC
kfVl+vm/65B1JV8yrKnaHBkehRjcA56BAVzTvkvsgcLoIDy+Cn9ikxl4Gr71NPvC
yn398Bv4S421sy8Av3qeTO//gz6ER7f/J4fyOV3JYVP6XmZacoSWkYUDwC9FX71d
V70+KapB9hWzmhGRW6/XkvJlKpUmO6h1j4tznGQkP+NufXxtHKg0N+rGArsUgO0B
1AvbHEtUx3qmkfyTHDj04WVPdnSmTRldKqxrXZ8S0x2oHhalaiBdS65yftF5+tz9
wkJ+6Wwb74/Vx6JKCYJqcy5deyb0DL0kJRXy9qURjMNq+e9v2C0XhdQ9fa5E3Fxc
aer02hb65PEfLRSkUwN5qTr+WCje0dARc+eD0tRGM2iKLui7XNor3dolKiAlOah+
VyzJISG5h2uUhWv8qjDAeVf5en9jtxsWWcdCntJI7AiQ3MWZFaDgJMQjQ2j+5vN1
C07iudXWrpI4rS43iT4Bv2Q/lvHKLjmGhKnNsfjnnv8iTgjXweqOoZbC7Z0UiRL8
n8zIjyLMJpJbV0G4EhJNMRrVDmo8rWx9HYfaz8M/P2SC8ZOXPfJrNHeiJj/nG4nH
6IiNuqLga4akI+ow4XWKncduXHYJ9Ktq2iBJy8xOc2CuFz2UQ6GND1P1VV3JpLrn
AHlAvV0lKXziq/8QfdxOjxQ3D/6ko8hkrPF4CipX+r8qY27l9gRNx4tWrGlz2fOE
pnlc7nTC/OG7o/RLMBboAaACOJ5dEGxj2753noqPbZgnAC0PH+vxEzT25w6hoVji
GSTanZYxsa3XifTk6tucNIdY37oR9MiLY2Mhywiwq7RpSW8mrRQIzLF4m1ouR/6v
tC6lQyPqY/8H6GFVo4VW2/kO50JZV5cCGGeJMIY2GVBKIVOdUrGrxPVxMSdSD3ql
oX3ck50nPyT2jTP3wsUBHWSPkQdSkJYTt3d2l6n2l+mDM0C2R2evQhqTPgJKua70
hjRB3IkvmdOfQQvfKNiRcguPY6ZrLO5mKPz7/xhohTpEPZ1FU3Y0s+eJD7VdOEFZ
R42xelG7IvBhMh8LREfaNunHVpMFzRnZ+lhI+LXogFQ6oczjJZfVEYoZ+GQQ+d5c
UM/pa0yvi2z2pnCOE1t2Knya22nDZRAl2kub2FwzTqswf4+7aw/wEVwMETuvoWjB
fVHWrI938osGI8AEPpeXDEp/baFmwQV9aY9AcRCgjOi2g4+93ShYVjj3dj0ZweCR
xCleanPNtQ8rv4PLdaFp9i1l6JPmvtD9rpIi4SaNsE5Aj+J6F6Uimv20y/12uJjv
Xtm0sEZXgRPSdkoinLuaqFe+qbZfBqBysA4k9XsidptJL3ClUMtsTzn7om+O9n05
6vI4x803/mq4Co8QOvEhONMf8NAq+zBVaH7boLE9A+AHC42Roh1cpz/eZ2EkeeTy
R3gfJZw3l/+e1O9jMMwi9jxxwQruIK1hJu3fE5Xlj5CbTitJqu7YbavfU0jYFKZP
r+XNPpFZy6L8l0VzY5Sir2JOTvLimWLS6Qlc3E9dStpfSu+727/wyOOVlWAA5GZ9
2eJr4yPP4rVpqkU4oOAWWdSOYMxJdQX4JKq/GbDeI9RYyGuLSkd1V7/7o0BzvpfV
YII0x4kwETFqcVdaK/d6kxvrZPzjvFbUdEC6dShwUnAblrFkGDRaPk7UofmoOwCo
nU4wTN0bzI/rzO25rbi8pVVi85Ts0BjigdMkT3h0bxAo65xRbkwa1PxBnRb9X/PS
HC9LFuCf5lPDXXByXxr5yQumM8kKFPSSexYIMH7ytoK/YCHn4gfd3LZ1hCFpv2Ki
YCmwTpbNASRWn11IOKVkBpDISiSlaAt2KoyTSmGHmIq64FufZFTvdZBMC6kVHK48
CxBcJP10INgan/mYG4ftolqVbhRIld8rj9zk92rW4C5ieQ/us2RucSvyvj12VSCX
I8P6pQREBSFKXuU3ZiBkesnNaXYjh/DQikKN2x5tajQ3HjJEW99u8qNr1eT+3Y54
1VWJSUCzGHvhlwMloetv+eL7rPoaWU9eCLGCIYYkG7Pm/ijFbLEzZTY9lbEgTYGg
48LkpcllKUi9JGh7n8Ame5pjjuFtpfxaKGmwEm6JFMX5ujExO4D3HGI07jfUNaUp
c7UURUuASMjO9GPQBtCtGf8J44inZBWktiH/0qqaHbZk4U7ot9wR4jaqYUJcMuUG
Pd39e31qTApVzsTgjKQqLXGBQGJ+IZevQYQviXFx2ssnfRq5C7fDEk2/qjWa/Az3
bvXW2UlSCHHFCQ7QpJT/DkVP4iS5tXIBRW3HZ47Jkv7zePq7wKcD2cKXAIhrTUh/
+KN6LD0ynqVT1T8U1uKkM0/YpK00PBhScU22LZSE+4h9ZY+H6B1VDGSvKLl/3kuS
56rO6TtgEOIo+9/kdFHJFOj7l7oturYAibVHPPZa4xrVkiImfVVU8eSJQw3Kzi9k
IhBxAcN6egjYKshtfvRPHP19xfRlcQwEAaG+RDTmNixqoPk0MHB0lkBFqjKfcxUq
UJ9rkFLOTymifqbwG0GeRH4Ikj0xlh2F94QHzZQU11GN917zN/FY+0p5hD5EM3G0
a80pAV3NZ3V14oo/vzI9hpPjmj89b0kXZS6VrS//wKSI4sBB28Anr2XoI/DIOUjk
Tc+56OkKDxZ5sYW+9PzaKVDw+DY3g5oao/jiDtZahhblaNc+XHk/3091HZ9lLJmS
qAUW515v4anvEKTBdqcdgHa+M+NSyNDm2iIioXYLv4ByQOUHaAvfFRbem0XHKb2t
KRA3vgJ4RQtuQaLaursWwo/tqRLdjWucVZNgxUBOYy9Nw1yFuSTEfyEiaEZP/KYp
5gYlyowWycnvO3CSL78xUaORHHQRlWI3wdqIfgpj7AeoaHBf8c9976fSd5VsyQj1
6X1W27W3G2kyifLGrbSPAt5iHgtrYm2/cGq7eGb9fEYOAy3vAiuW60/Usr16jDr+
HHKsFty3RJGeOn9xFJvgtXLJF5GK8hnL7cW7h6bTse2u8bgEfXwVQFy+Gs/Sk1/s
uvKju6wtbAKaZfkwRwr3u9CqzqKW7exvyZw19KcUX44Oa7AcmXfe5yPqz2peHW0q
wFVizx8bCp8p6LyoGTC4zgaTS1J98+ccEWP3TS3/ijODVjBeOd93eNVjPHosd9j5
v5zc7VZfh75H1ibcMjauIOtIgJsPRtS1RkseCKR0apO7aPNzSkNrhF1NPwjJl4Wu
7ExiTKJXOyWiKblmzfsvtdJHhqdCXec1ZPgMfViKT4gidfjw/yffo7YNjSGumY3c
vj/781B/mjOBObj75otmyqZ9gKIa9ZM7L0ycJDdC/ZN+4zd+JRqDXKp79RejwPAk
FCU7LE98TWXhsSSqSM/rA96BlCegl5CJnChB8JO18i2RXW0KVkciw+r6C80Rfyp7
Fp5ztByAJo5VHSQCeU14cJsbpnB2K9CTd0WQKS1736spRoPpeFFjtAZVuq2mvUo9
keEUvKxz9n4BOGqaah8bVEtZPnuo2PS6/kqJpn9ISZZUoPZ96F5ou0vSWMGZdnMp
ktmTEw78hNyh/iUsrlYRlwFaU+mn0KEXYohWDqXlSxpTpUk5IgXiMisksYIQFTz1
DYL1NsNZEy5RjZk2nLqivOey228No/Jq3bjxTp6T4Uy9lO+jgt66D4cazYTh2g8J
RMNoKu4EU0k21ZAt/u5iLP7rhd3h16Y/nfg57HTaYXEbg2LKGObHmwT75sz4p0ca
T5gd4FFdnpU6WkDW9z3w0BNrUoGHC81pUDXI2QF91uLpT5/E1tTct8yXTBg69KUy
Eq+oVbOH/yUnzl3rfPRvR26OQZ6ldK9JyCZc9o28IxG5Sz0WxCyjMJhO+cbssg1m
fj7SjgJ86xxRBhsS5XNNd45jgwGWMoAtHCSE3MzBivwQ+3K2h89fKFX3q0RYJxKv
jV24cbAvvXkxWaCdV1cImLcaxRdSq3gc2iB86n9yEDHB6RcC3xk3gLJWqgi0weMg
HRw99HcIduB7ShwGdIgO4pDSjNRNhy4cYnVFUgEvyAfpKC1hToHZ2nTwlq5NijSp
2mjIkv9zCIhY1GcZ36BaSVyNeb/PV+w5C1ahEJvGX4bp0re9kqNIr6/5sH0ENZ1r
UXSv4jKt5QcltwzcCdIKlmSMzkIzdM48fEqEjEd8xJyiMQ8+hoidTX556swgA7VF
gvxoPPEcT1G3TB2zsLjbFJVAITQekSN2aBGrDBU8PHqG2xBDRGNkct7Yjzyouht6
/hmxeG5t/a0EntJ7EsvRvti56GaEGZuM8YojQsjotzTBXIQw/l0mXhINPmgmqapE
Rr4+KFHrk6YEy+XTnpiyQ970ritveYOCuAe2BBpt+25hr/3pF4wjmPv20idKkfrZ
Q0u2EdQ4VGgPVKpBDS1pWY4aZD4C7FsP7vL6JqD8420PQXyFZaO+jZEKhdNp/qj6
xJP9D7qiNqIuJ0VTe9udCo6CJxbJUYtUMgkGA0dLcO9/BGJ5LtjKxF4Mrq8/8qTs
D49Nl75mQa+wtYllZ4L1+aqteRD9GxijZ/q5B6E8pIKzxYzg/I822NU9n4MrV4xw
rlCh6JpkZH2BMXDBoHPcSiGnrDUgxAgN4Xevv2U++qVRyQAoJ9NlRnBm4wDwH4GT
dlE2pf+2QI354otKAScjuzJwq+FCfwhTSl5TOGfc7eEOgekyXO3YANUvZz85TX7O
jk+2P+2iaY+i3S34xZuUgUvlKwJFssTNEAgtL80uN5mQexloW2mhDsZf/Y7WgscT
/67n4e9xKnYgYVD41hBI1rYUg8YjjYBIAYcJpbkL7TQGYEPHByLa1QaOh+omxMAP
Xhrs4nQOT2y5bCraK3IzuucpGvxrl4rVhMLvOSFyEh/tXNk8JVbc8G0F+JofpqV9
Tqrmvd22HFo0S28p0hvk7UItatpM9ewzkd3OAVtHWs95nG/KGyH5ma+wA78maKT3
p6EXwYOW1ZG6M+puALmZ72WxRFMdIOptSWAL8o7wqoDL/kje4Ez1xosqyO5E7YPa
kmRSx8YPwZWDzL7lcLwPuXhgPuE8zLoejc1QVfplORcz1cGoFtVom8GwEluCQgdm
6qbF8L/E9eYTymVXHpaxbttHM8TtgWj2h3X5rWYjSVwOdVKHAd9ONfhPSrW76ODy
zyMKqk89tsw1bk96rahaR90ic/a2txVRlXSDMlDcNRICZv18qn+SYEY2EzA9tAQR
UBXXD13Fh8pWS01fqwHvRK6V90kXJ+i94m0CuFCcyrTy+PjsTmL5RACg0neqU8zK
lWc0E1mDS9tUdeRmG63SvNvPGD/WWr4YZYrr3wozFuA6rjr+iFTCtB3u3L6gf3xs
TIDocKean+GwmIvp+MpNCyaUc1HidEhB4RJsH5uSMA646K0El5uw+e3Z43lia4Yp
RmSXj4MzUebQxFh1jUvm6Ku43yY86mpXmZfM4GSp+iudOhfBq+fmoOatH3KpKOeV
yel0/7scNqsbMzql52YNyjN166UbjiaGmFSi62jV0Fc7n761XBXlFLWgss5Zw2Sv
Uh2sqS20om8hcZJr2IsGMlv3JTDReNo9I15daBbfueW193byvfXltLOHpTH2mta+
GlBZYgjWJs8/p81Lu3+PiR8eJAieS0x1aNbXqVKp9YSc48r0eNypLgjuFIHiaeTd
j6wbjUQqfouxTCIxzlC6xIZ8FeAGfPbRFcXK2eK8cyzVe/kF00RMo5lmSl4fpT1c
x+lnL2bURgC/NHjMPDjPavpVxg7qfcVw6DlmHcae1TdMlRHspzSoTMS4rXRu3W/W
RkRn4cP+nJAqySPixp3g4NOBCa9tuugtWJMj3ZlhBqlIsQ8rDkzDlQNtlgk1vSgH
ydbUjGFwGzULeWg/B3YPJlfhuGJTCKSae54q9O6HReXF9zf/kwltdn7OLpCCKwDR
EDe4rgEcLgqPliDxwYQx/pgYpGsdFTfSpXR8DHhfTl37OAYf8+TB1n9Xk2MPs0BM
dRlVxIGQj/l0tL5TrLN7u1OzTfIHgcmG5YX8xbY+1mRUejrjWDEE3k++eZd7RzDK
YX0udo8Nw8TVxbHFb/8a30EcyR8TrWv8yOSaUW+mBWMnvHHCCi1FJXok54ZSphjU
PgPFKlvVW3n2OzWgHPLXqPmZjr0fd1D93FBmJMcyMejlXIX5L+RcfHXytYgPHS30
y0oGk1rI45kmZ4YjAvJPBrDShWPggZe1qTnJoi0aQVYtwgJLwsW7ekDaLktJshFz
bvhxLm1hLsOGPDnlPY75Ql7Nvwtw4paJOpWEOJePKe5doNZjad8GAe+NyxceGkhF
uhr6EORuFRTqJ5YOV/C4YPtrG7Zw6HmAqcXE6rBr9k0ObKyig8HeDutzs+ywY8nN
hFVZoegy82vDttK/iXx1hZIKo+wJDgRhtQOiMSwPOHxsKoRpjAtgngFU2tAL0l0W
pzkrupCbCffG5BSZOfqVifk47tHevMGhU2eXRWAiPrXg6px8bWZROX9uitNze7Lt
1v23eO+ru8pj5wTHBr5lIMcdChz6PezYSMld6Zm8aA1MRPwHm2TSiIu3ecJdQEty
KlS+fgzGUHfGN19vgV+a9Cku1groolcJC6PkjjeG8gb6QUES2NXryS4bToSPR1Gs
ALH5hUrg4WNpVuyQPztFPrAH8a0xKsnVECWeofxmGVTOFQ6ftQJqd53rqIpH6y9/
B3IcGCqZ1dHVZqjlPy0RShWwu6Mf2VFZLkHaUCOv4/SU1J3uNuU1ybss3qiOTBMk
cMpJkwyrrpXoqqx23xIOe42IvirzbOFGzLXRY+Y0mlr1Zvwr4paeK0o4eDok1kqK
/AYD4xgcqmk3uF/fEkNVQJLgXoBRL1aQAOYcM+JVazI5wAcu15hv5GGo5BzyYfSK
D+JraLWB+Cpue+TcO6W3GAjA11SxFhdGAFCLBa0+4KytqznUt4+nMcQ1e82S4+9E
H5We4ONReEP48Eu1BqZ69qA7PmgyuNkMql4g8RixwUZ3TmH4xcLPJ8jHZUJEfTet
nY6S0dZdtRUu6kUeM+YoL7LLFtoWayTDT0Pq+3w7YJgspwkEQFHLV2BTrZSQW1Rd
jo//qeny6saLa+KXPEA+Jc/J6W+DpO8IdxjFLZVnhvHJpaZNG3xsB9fw7NNActOP
V3Ff+37GW1EZXNiAacvjfUgz2mnmDe6vyQ+5y8bt424UZLe3HsdhxbprXJBpNCjv
UVrVt8+gWSPrTdFK1eUYm9aIvA2PKgGqzZwLL1CJvP/Ye84FvoyTp3aeFk4KM6hG
rhBXs5gLZ5m5XMRQMxNH/dltiiF9Mfzsx4p51U1JMGqf1iO25qLwux8C07voitx2
nWnEVvhuQKDlru2FaGVuG3e4bvpqixseuajKduCK75BT5c0cMadkcWeeQTa06N2A
GvC8fNYI/xOHB6X0lKumrbqzKrJad1IrtlZbqkIfCWb6UvVG/kBQ86CPivlx5rzH
506H8wG+K+KDzlATfeMJzm/Hd7qECKC1wlKmCybmKfbWT/Euab6DfSoQVjZhS9Rs
1dNaV+XdxGunOe9XgAxhlfUD26DMND0qOgg4M46FEPtejQAbbZ43NPRK5GIcyDaL
+BGkXM0whjyrJgd8QXBRoXBo4QGMplgz9oyUbcpyjCGCjYClOXDejehHiqyZ1E0f
r5yb6C1qkdEt+Hk7lUiyIyKTv9GvtYVTO6G/EtLaakpzcJ8Qqag6y0RHIeF0xH+b
Z86X9mMcy+9ji/ICKPR+AxAiAqxOYTpnxzO2cwg7nh6FTDOvdkoi5Aez7GpYYmpi
h+PtlO3ltpEUxpj2gQ69H1KkJD1FTOQCAAzgNtb6ySObR3Q3hDMfkxbnRXvrW2oH
qOZnTwW+uOR+rjToKNT3RZTXnGlk2PGXnPQWXxKO0F4ZZGf2LRiPKl9YdaxVskNr
vIKSJN1U8qgxBgcVYA+i0XPrSZV337WQDhyFn9WnNMblTOFslAY5h6ZJnFIpIcs0
aU8xrMTC/IZmFEZlVCscpP7R1SdaFEc1wg6RWA9mVjudnlGW8w4rbAtYNAqv1fSv
BXglv1wqdG0Vybu1DsD12CeHGqW9Mjv6GSfxoes3GlJnnBEpLdsXdGGfysMZiy1t
FPNNRW0iIOZjPhBlNWHktAFfzQnVKHkiLTtesQ6GINA2nEJOkWLfPHmuU0kknSzQ
reQFJedFLinO8KXVxI6KOIafuMGPMLDmFhRQuZsD+GHlIBRiyA/tewfvK57KsNNj
V6KPUatnCOAcMHUuP4zGeruO1FfXKOQB9aV6uPeO99Z7AQw33OXQtx28A1KWV0s5
KvJmNQq5jz4xkPhs6hdiZDS2Pdt60NvgTCawDLIqhWy9xXOwYsePdzC4yV/jSBo+
QEkQDVrccRDowkxe8rm1i2IoIMqbdUJw65RRv/l7WAF7Er0+iLSLw5z3Lbtipy8C
Ox/zsjgWF07v3Yy2NyUcQhADehtHOz+z32cDhXGrQw3/MB2uPaEpX2DmdXJsiLfK
Jay1SwBzBeSE7gjaJ2vVTZePxtvGGmOaz0Xy3TMykpoYqLyGKSqdhXMidXAvUa68
AyC+b1unaHd13k+4+Heil3oYxS74Ljj395NwRSo6Bc561NXX2OXOGqPLMmPs+EOt
lfpqNGugNsYxgj0sZksEDaGthvgnHacHLDE4diz5ybRTVYAxB3X08D+HhVlTnBe7
ljrqkz3qiS/odrtJgPqOlWDBPa1gjfqtvLjOiJ1mRckrilSGZHhXRx+L5OwSxkrf
9eSXOMuS2clnfTibF6mz4KXZF8kQ3pliFbsyq6AU5jkrqqEBZvjfY2zcMEvhmN9i
f9ANd1fERCagfqN7YNPC2ZukrPjk2oWfh+V3tI7nphz+09Ur4SZeE9l3DDKkERtF
VjzAq98dVqnxqTZzHKINfAV4JPKq5bZmzXIn1PPxqZmR7iEtRN23IlCRpPNFxlyF
5NKroVzFKYC/iQGer0wDptldSMkeaNQ1V/U/+4fKP50qqmd1WbNzuaQ2ctEcN2Yr
PZDTe3MSLa2TvQZMwXtDjA==
`protect end_protected