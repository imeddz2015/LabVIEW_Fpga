`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 50640 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/9huKRhRMtvnNqb3Z+UU7TahEoHV+T8U3P3ufru7l1O
3DlgtZzb9QxCbOjthp9+wDkjygH0eUfDrEl1ovhZG63BUSRxcTbq2lzntCgYSHtp
dN8E5Pg2oQwSdTrHgXqy4KnUh9myVdj3YljTOX0B99SIPRsYmgQPlFgKvZWrDUAa
iLba1nS57Dc4qhtc4QqbPSaMl4R6PrpnWXkTWFA6dBaHtZwKA2xQscvvPAA9XP4O
r3pLD87X3HDtvzjk7CpLK8J14V+WLQ2fO4KQLpj5c1+CCL/rX4Ihiyp/SgBhMx5r
5f9HptBWeAyWYwyEB3kKgL5MwQo92+CD39oFEmjSMTH0EMsaTkWOO4wY4HTOFhvP
S9oMLZ82R/O7JdSk4Ym0Xe+KUGTB5PUa7WKrA5Y+GefT6t0ILaRQPlRMDwJDl1XF
VUXxeylf+30xcNBKXqGHVFnCTZPins4icUpyY2cPD2VxSqs/9uSDY13zlWKUB6Et
xTTBVr0cBQITZnZ3P+YcYXNJ2CztUngotgkeN7Zjou8Th+Yez4wEubiQX0pSNRo0
BAME/beFWeDzi2qasByIv0loJV4EP2aWTkTy8iiiiiGfvWv32IFCXno+fejdY+W5
7VUuqXFuqWUDdpbWbTg06CuxmfesEj7RJ+qyTebcYHCFQGyupUFbmYrOaA3XO7oZ
FYpx7Az8+Y5KIenSnjQ4Tu0oMpSySg6UaTu+sclq57qYmt41aB7ISC4BpdgzyWGe
W0pXq4Ilxtgy2qIYLAxKbK7wLRZ7OwZZ0CIAE2QgDHSDYR98300XZBGBZMR6vHzI
os0LsUpg/CPPDeNdRiYQMxravHRgyNIWdorRoXVCMapqH9Js7TarddWkBub1TFVf
2oNgcUXE4T3g90ElOZrtEhyMpiXpksdArPPewyU/64CywwPEl75zzygZLeKv/4/n
uaZNIkOQ80SaUy6Yq5RptZr+DVrIkwcQKsT43yzz6Kr7i1zNSApaxdHFv3wIfZT7
8WqkBOQW3fdrWzky9+mCfseHcEMCYCFW74Fd3oX0b9DDQ4abVQiI7yp+6/Zcm/H1
SJ53Qxxllp+nWjpTQh6gkOiowiErcmMOgH5kpXzGvq6yJxVmJW5LBXn0OJ8NfP9c
oz1VE5frRh1btghmfRYfNO7ZDCoorTLyXYNNSXYp0PynUkyUKHvMJ/P3Po10npPZ
YIBiaxFtwEN39ruDyWg05sm3RbeZ0IGKN1JM2D61MGIqvIthi0JsWHa5pCtncomW
Fl/1GLLalepfkd1LpCzTED/2RSkU9dOt7sN6BLm47Ki6+r1oqk8yvWe99aDJTGJ1
dYSttdnFM+Lad5QR3SBKsca+sPPE79oEptOt1bF1KChs6325zK4F6wkNyV9laOqd
qRn4T6RDEslAdSkbzXJMRMV9uW81RpXlQEoq+0+giu/lljU7ugjif5myNkNN7ttJ
pPDnpdpLxzIBx45Foxum/dtJeay6t8ueBV0uRtAEpN5Er5VmXsyWuHHu6x+xNKWX
NaMOwY71zJpGb7VZI6tR+4/dnnVD+3ho4WawxWhiDbH6EeylkpGrhXcLBKq/rkKk
c2sgdSD+oS9+vsP2fGInM6QQw8F283KLL3b0Edn6z9eN9kZXS0CCDP2xMAM0+vi6
eNhfgsWCLQI9nBFUhXM2Tn+k3tQnjbumeYH3FeRVgRPESrM4zclWJgdqjwUvjz16
SQItqcUtZbFfmRUUER7eGrJ6ik9mp5IGvX/Jt6LYX97sne5qU8H1ONA9fgQq71K6
aYd+/cjNL6yY3p5l3lAwvhgLF9EYhvKdFRKqsqWrnujEcFpU/RqHjb3Mg6EbV0/l
C4LJPZe6TXQcmT3ssi8gDqONazM1V/gTBl5J3WOkaGUntSRUJ8+RO4LAu0b/cRll
kJtgDe8Aln3DNAEjh6PbO/x7p/+sYQLYshiB9Y/oUv0Vifl5QCycs68vju4KonxJ
yIGHCxVXeu6NOpizn2HQywp0g9EGqda3ah40NU3ob0MHwyhvM+qzHzrl7Oe5rjLg
KLFLbPkg94/6e68o1LpdGesrSQtXtLzXbPwkkfZSzwZfGvIPE0DotarOCdwzoYNL
BkqsMtL6vKSS0t5OzRDar1BqU6f6jWvSDCZg5DPHTc8HGHaCjm5nSqHqqn2YJCYS
vvS1So/wZpxm9jel2YNCcBSACuc8yOytHtXHzTwD4XmGrakMO7gSfjUq+rRw/sQk
ye4hjtVYFKmUrNS7hcr8qL2Yjb4Y/1hrDhv04Te4bQKBPV8cetC+rQrW2xQeoqWU
d/qqXKaEBm1V3urL+baNtpk9V/1m3fZDBxlTm/Hd8yu9fmhXZz48PS/Xa/fAY0XL
UBRxxlR98SYN6aPVxSXj/4eAVQAiK7YF1yi8IMh9ojZ24Z7hLGHLWjeLBZbcwe9m
Dej2z/ZcUMnwBLeTh6dnw99VeYE8S8uzuQWs54+bmcdLVS44CB6YmRfgUdLK7gdp
E6CfodUr8/TChJn//viYEWd8OPx+fIvjr4H8JHnPf6u4yMupK6uLlKx3TYPABtqO
3wxrd8HtT0TOns/lvR7edTvV10gtPCcgtg5inlHp02XYEahrecqnZk+fUk3H5lrP
NAFIW+6+Bx34ha2EqQrv0tnMJxzG9gXdvPRjc3lIRxroG4Z5V98gtiYvF1G68dmK
lrEx7yT+Ac8kVZW+9Pz4FtQIz/tNxZU7mxAcB8WSg9Zof+j8cf3MxhPeX5X9py8a
hokg9mvBTXFZVQMyA9RKPV5rHc571EtD9RysWuWEDrHU68Twq/g1KT+LDu1S6nX6
nHRKeJP7rDcXIYpkAByMDMkxECF5LQFhIxDuoxo7gDDHk9oofwiypJs6S+IjJpsV
JC2q3r1BHQXDtU3pMYALf8xYBkUDY1GvJYRfRsr5DFKsa2QeAB5yzDE1lvBZOIIL
SYYYakOvQYytcaG2YBtnGtVZGDGe4klx8TRWHizAivLJJm4xnrXWp3nN0GlUun/6
vOpc+YyL/N+TwUq6DsHf7/TRxADjVr1RL/EI55k0TCsf6o0FSvX97tUsLG+6g5hk
q+PTqDP+N5lBAOMGwgrkKfkeiMyC1dAdCTmsXx5HK3HotqhRLV7Bes69P+t05A2u
FnQzNaENraIl25PKIetMjlMZ06/yApF8uzRl3cMeYzT2e5htlUwsCEO71MILUtPa
N9ZO+d1FGnF2cpnfpR7X7i1/wS9f50ryXOJFIIcSS+QSAcsuPX/BoTFNX/FydxBJ
xHv7ZqB+Z3IpVaCr/MqKPa/XhUzzkk12BIOmQLZD2VhypL1D3Zfo3nqTk2ZbU0qN
MMN3ubDVvMdXA0yIxuQFf8nBpGW1FTTF9eMxDRkmWRwJBHvHd7ydZFcEMsF/LPtc
mJXpAMaSkbDmvi9Thyxxc4+FhS10FfPL46ABTz6NVrVLJxTjgh0B4Me10onENNod
HRKXn6dYAD52IQEgqb2Rknm8jSxZMnRKBvH8T2KMEfCMHfRyeN7rFzfdT8ShEP/E
18Y7xvXS834EXpjnOzR6sIWF2kE0hUSBbN/2GjWWztesnM5P7lHSbCKZUTvMvTpp
A3c9/eRFtB7NF6y1gFLEhx/ZV4wOi/2lnpPddLsdpWF3vnwrvJiRNGmyLfDtioc/
MVcWFXGRh4fkW7fhcLoP1MoZ/ygWrad4rmf6vxQLK7dT1UWVHtmdQW2mPPWh9YBT
psJ0vNKOq4uCPqRp9NEoLC7vXHSyWURhIH6IxmlXVJaxHbuKVRihCkCEmfwnLRt/
ZDTWbU18BHw6JUr0E4LHYz1Ewi4xk++BRHZmJOhpFwXxXibHdXxy5I2Az3MTj15b
72ZPMAkpozR72/Wr84klDxyUGc/G00O13zFIRZ8Z/YPRO51OH7TYCh4KO+auFqOZ
QSnJaP1NRiRYm3Hkbl88TYOa/PQFs4ndm7Brmu8stbPELSF15+nRKsqY5bJ3Ibyb
00swI/GSUk37qy/kekUKDR8pYzOSZC3LEYDAK7kDLe8ljGEhbuc8mWIp7XffyzSI
Kq7q3ZVGSCW54cmNlLyk9o2w0JLidt08MI0yrYVcCpwU10uQGjBUhRe//UqHDoFK
JmMqJgUbD+3z17xfVQThnbLvefgJStP2yjP9zm/X2Wx94dkQinOXs2CNyUZ877zt
YTIF9ChYK6h3+frAF/ZsJ96sDb7qWe/tBbtY9KqlY80bxkM/nIr4Wbaviry83BcS
7wAejkoVOhEy9zzjjspSwkW771O2QEGEMS17opeIrPUMzOw+FwWWjjs55Mx5YJsT
K/lraD/W+yJAFTFTuT7Q29tpeV/d56XHX522xKZSX+JBxkCRMtp5arOFYlJEqyJO
imWzJ8WdgHFRKEb4drykctSZz7HGyJS39ZKXyYsClpkSk39DL9wvc53orz5eKp41
u0dB4JnOwW9Z+4YsY/xoh3AcQDeAw5R+eRvOZseqB5i+3tPCbkzsj2F/Am8jd/7D
s15r8mRjkDJC3fsO03L0N6hNl3h8MImGJoedUeFHzKrRYGX4bng8ZkDfUDWt25x8
UaB5mRNALVBCWTeImMcmS+znvBhBd9GXQdODSevY8axocqyHlthKIDFv7EYQGYyT
dyIqrfe1zUMRQ4a4Ozyu6B7o1FZAdFj36y4+kKVZPlNligKocQcX/YGuLnfDeZmZ
P2v1EFMQz1Vj+2wNF/hp80Ewlcmnf0Bb6cTfFBivVlCq1ApG5/i9CI6YWUlnaP8j
KnKNdEll+ieZ4RVpL0lhOIq9Tg9JclbNUIdlxZvyijBfWlAhPhjXgbnaLA8Onmr8
ZdNzHsM8R6XgkphVh7hNNwYZLEihQNvOVh3Azz+pkrHQ4GyuRXgG90CMMHHSReiK
zgJZHtHBxIUFyqPYKNPSImj135ABzYQ3vDtdeb4CH/Ku9gcztvlPvvHs6+SB0SpD
s058T+7wdSPp286k6oWdhPGVC92P3pPFpWLHEujliMHr3XUYRx2dSs7/Hycu2Yku
Cd0cnpe1Ol/52g0702zr1Qk6Yl9dpRV4/Wf3vjjAadkQgSFudRLa9rkK6q7gIfJD
W1MKc6KdXzxlltdlkWzDmasaFFlEPRE0rZu6NSrCrbm8v+Gk35f2IIuqsEwdbxWp
edyJBMH611mlGjHyw4tiOnaGydM5bRfZ76MPCd98IwwFjtGrfYeYgBvthtMKQ2Ne
ZJhcRLldUXgrJCwm3OrFkCcdURNjqUm3TKka/aeYSgIMlXl9A9zaE/IXbGCLAdkb
qoGCVI1CoMqhftf3QPGs8PkA/OGVp9eXlPdjzg6BnndXoVH/7rq1Qu1CPvkGIxmw
wSMuOkyv3vB6mOovlgN4BNT7tZnZmjuInHtyGfDvvG07Hwb3CQJSo0XXYPKw47Qj
sOSyEVlpdBgzuTYn270LeguzDnK7rtd28t8W41/0qnmo3L+sej1CmoPRUu+AkD51
L9vQItqtCeyZfh/VPsxMQcx0eubsAWcHGdCkU2ElGkqZAVKzI05Cs0IEL8gZ1xM9
HzbDR2YBbdNwfVLjXK9W2nrfltjJpjFYjvhShq8+crsplBPEu+hd2EkquguZN35s
cERj5ciFctFDhh4R1VZPL9MIWY3UwTuqOCj/qDXwpK9fop9VMVRFNzqPbxOZALFe
vIJ8LURTApndY3rk3ePRUvtgxLayPBMMbDcTPLuzOO/swckgqTHK043O+qoMLS5Q
iyzmyxOwJspOeJGehjzyD1xxGTmNmCwsIxBRQtw+9OzUGXO2etgju8kL4cikWbnQ
kgn1iEmZ1XULBvAqeaADJ5jw7qbqR2+9gs7+34dZhO5ryOA4nKDWbz7nOOVTH8Ok
X/4+pDJmrzlcUk+gVGVQX5Pj+cplWW8FrDGdUKXcTpCQfIIoQPDbKNFIu7QDrmFI
nCEFY3m9MLUs9JvvDDG+HToMzG7lYl0zBQXzunS9YAW4EC9MwzSixbR6yPMLxjv2
gOU1Mo0pCoN0pG/46n+oYcIttpXh7Ople0Faf2MO1KwsjyIgst/4/Xucv69XXskx
ztvXgUMNWvxBRXckbqGMTQEKdg2+U8kFz7WWjXg7nntSZSXAzFctE+O/qN33Hn0r
Ykdt7QqOys8uUSqANL1VRBmvho2cizXPL0/vKDpufBylSMHN95t2e6HCk8ZG8AiU
DHPeeOqerX9WH5xoZw+KaVgDlm8PDuve1H2paqO9e3627qJsbqPLZsCkGLyccLFF
O1frbnu8SpXHLXmIh+teGoYW6eLpUX+4u28IAwsoktrG0kg194qx8PgfJWyttTsn
w6vJYHyr9GfPKahfNnqH8YhwKfI0YNpHw9D/xqVCzL2h1qpRVieAGTJ61Ymp3De1
5gXXeLwMTKnAr/OUTPXwM+2l40P/OERQXxtyewQ/uxS2A9tYcGhk1AfJxSnplTq5
Xl3N+GD7zBFxW246Pqq0NnreuiDmCZxqJEgo/CV1vWvg8O/eNz2F1oLIzNE1MTLR
iLb05AL8VE3qtut2qGbMhLrW5GTEZmF3IDUADRCgI35UxqdK/jmuHvT481ZtzVHD
drZYTLtPC391sev3dZd9Tf1HL6SgXVpfJHEt7FZxAQNPEzs9QzG2KiWbiv6BqukY
9e57vhWToPyFP1RRQbvUbkKc+voUbBvBDIB6t/eoEHsAwsPg+OiZvmeP2PipKa3P
d9drAoyj6RzpofrJGa0uKL2u0mE6bNNDJpd7jH6aF98hpfxKalaCMglqmmaAgu1m
pkK7jTx+hZhVDRaat3jeLkzdRfXlhYiAxBHjz1M7xgW//9a6Mftdh6xcSj02JloT
t1E95LT6Clezfg7UxKChcN9yHRq+FVJ5RwSJY5hbyg803acwBowQRT0PnXHVNbF/
IAJa4hI2JAs0K4gX0MOKzJkykLIpGQ9hNNzny4F1eSxaf5bMk+D466dvjBpOMXke
FC4P+5kcvUbjzEm2mHgdSy62Wkb9qzXhZhIHCuYa3cbbTKJBuD+aR7wHayIDuDfd
+uOhUdHasgMCUTmY/GyU2gNTm4fNeFKidvfCUSLx/7hUKkAliC5M8Gsxo1+3r/mm
+OX2wbVGp/sZl/b+dFcwGsSf+MD0T7GGpvJE11PfIrxJyZq2cMveZRzR4lBhCgCj
oEB9UIBznBxjJszFBsFjFkI0K6XEdgZ7cWZgtqDO54lJiPNYHxMEmP72uQEvKGHa
hJayY6Ztm/lD0u0Cpq9dLR6fQpTkmmt8Y1XI9APPmU4KmXgX0zqAX1KLRaxdYeu8
pklm9lYxalhk9KFJQgR95rrpEFK2xN1Z+4FxzMOQqbCJByKpuCKgbO9NspVG9DsB
K6HD9GDagQpEiIKUYZJDiiSVYpxwImeuRStlDrGucqqmZ7QP5ycAGWvMjaBNioNh
0JG8dzKuCwlkmD0A4S2DxtAQjyy/UHoAq3Rbaffi+0hY39MuH/GxGCQFVX582HwU
YGuFTVdR367qC4CHy8KZ23yMVcb41FN8cYCdaYe9qlvyqIAPN3kkuDJoYs6bxDfm
q1IMQH6SJsB7CMTRRjAyYDR1aAO7vcpweHj5+LTM7EeNL11nZUCmsKsAVXcvj4lw
/tcXXmKRMn0rKGihDorwM1XavkbWsspTGaVLjn+a6Rttr2uZX+7PQpE0+VNztaPx
lhsalKWSU6U/9Z2I2NV0YJFpRvcKxOIynNps8Z+/14QIWbWi9c2k4Cqtr1nqvIN6
aaOp12X4ZfjFndXOLIuv2XuZ/f+hWELTtB23oWMAFb6ifF6+ZeHltONr522h55A7
7ZeeihmATxiQFj0DfEDu7GAdohIeAT/44X/HlYwDfqd3NmjHn16cxa6pWYHsmy9S
a3hCNge5JsiXVZ5Xks23RNitgbD3qb45G9Vt/kdgh8eSMEK3yDvPwe6QRfdnko2Z
OKFU3nngvDZ6yTdP530QVdwLalgpjVAVlBhpFbLHg85fJP0jzynCvCkWzbmfpwQp
pgFjnXEZd7B6xNL+6CkRCUmKp5BvEAhqYU5j89rNoPiOvrFUeqggnlI9LmglRb+t
N90aOIDQq5N5Jmlmueaf7sgCPLz4/207IXB6dvlMLmW350Spn2Sey06pbP/KWcvW
8Gc4wW0x+iFP4LU1A6xta/sQBbcc2KY8KxCcV4xsmSCnmufX1lTX3H+lZd0IRMHb
151Zo8tJ6tLnguPsfKyDWHw8zZ73WqGr87z/K7SkhRMhxhPPJ7He692vIjLUjMEb
bvO+puQ2CvilNVXrhRLv14FFcmUgWGfJAJw/JvznYNr2mCvYDeclzJmbkt4ERSMV
ydBUQoiD44BE4ev8G2Wn7bn8gVFrP/dJKu0cRErf3G+LNb5j3RlgpZMre/yE4pF9
NSUGLz4/51+Q/Uuwqt85CZ6L+JIHIoNoct6rounOlHH3OXEebK18faw130U2DS8v
YOr8O3qGwLFiPk7M8bEG8YZQ3oezMt/UfYljnnFDnFvFkrTwYW/5RCqiyFXzyWx6
/n4TqIfyKfvxqJiqUhKZo49BzYgVVdztelko8qiv2CZv0tLE/KzXKZuo9gc2432F
u5vfkzC8xEgOKHwdHPzhS1qfR2dRTVreBhEPadp+J5nHPTNVtpGo48dgaF1JH9Iy
qEXVVf1UPzc17sy1eiDVpJiAmWCSKMCOw8451qZY2ehRnl30DxOlhy+NY/eWJ9hC
R+MnC6Szi7mCX144+ZjA2drCwPIONe8HJXqPBRaOWL2cTcCPKvNmrKvLQ+tL/Csu
S5VVswoGIXzvGGRWdwZlzP6LoASLxrlvMgaKhgGNVhdLcECO5jJTSx8TDlBLRkg7
ONerjdmeUspZ/9zTL0JKhj3JbibgTSCM8jK/h+gd7RcfjRnExRBc3wNvqh38LeFm
IvIRy2lSDSyTH7iPHx/YhW+hmBCL0+JayNsJd8DdQK70HmzynuzNtd0ZGVg7vrLT
WTuLP1xum5erYGEHZ7LFKITkwaMT2rmUjQglHtl1qCks3AxtSE1RbEoS4O8WRnaV
Hf8E/eIDJszwcJiqJAJ+mDyv3I6ftCo50S59mk0g6CSyELRK81jmtmY5P+UKQLPv
Oa+4A9uZU+6AxTlCxTYSmaCEzN/zZ4uq13iRGzalX7OH2ZBybbJ186mlVOSoykZx
sfq1SVhg+7Dzq5CVsKbyF+WDN0AI4CTm6zEMxBZvpo1QoNcAmQmG4oV2V4jGwbtA
7Q7xX8gfHPMnqaGUtZ1gG7kncH+A4lmwg/pplldBBCbQlfRmn6OT9nHc6Q49FJ4/
HUN0SnYd/7B5jQqilaV/TMkF9ta7bG1vWZ4nNa5HHillctuLo5yyX6LbksqgZVmS
9Zk8lcyFLl0SzJR4++WOOlHG2RnA2yvHAye/AmbDl1f2gcM1Wtb8oIbHE6ALQnvs
ICkfVqg6Q+81lJLekjRqPq37at53EnL5bpJny9o2gTJaQq/GQWpWiFQKmeQKPx78
313aUsYWiJUUS1jJ0ADgo/7/Lp9B70hYxQKz7uWAJJP8DQhp8pSoxdAnoNXgjyOW
Tb6OmcF/G3Ns5sFrg3mZmr30n1PgxQ0EnRyVVXheSiSqE9ZKbn0T4KeJKHz+pPAN
edu3LgwlWi0AnkJMYxRQmrwjbLTI9QNdCAM5b2IzgfMABy2eVY90Aj7S2EfeFsST
UdUf/PwUGfjmDe7McL7CBZ5Tcxf4wrU7kMmKXEBJWEJCiMi980EbPyGfzjBDI0E0
PH9AxwXEJk0cB1arLVCc80/npjevaN7eTISfGD9S3Fa42PC7kxX9JsIj7CiP4wSK
w1OlgN+4xQXMxkI0YiVwsWtu9gOvRGOnLgRtwdPWy+Zx1RP8K7WdkTO34imfVg9z
CdvPB0501qsoPWKrX+SLVSJbAr9B3kpE3Dt0qtds5azJ58kczk+8gqufz3ZQQLkl
1L2qpkX2zkTr+1Ap41Rz6QKmbIqlJPgOpUnPQJoUA81SKeGh1mnjbayvd8A/FtcG
6IFoMimyHRz866mJVmonp2vln/KvfMRpt9JSRRLekHKUV4eU5nGP7Zj3MHULmocF
wHKizyzjziki4r1lraRO51D2nM3GvxAdanpmzPnSOpF3Hl3zMZJgyJCoH74GJ5Ul
VJUM54Tn5m3pOY+X1+XmK1aTCa/oNmoa6ZaTkh2U0JmGoOC0jHqcCdWnM26sGN9W
rjLf63TCQI5JODbiDrHofhtTqDkjs/sfJ/j2mdTNRb/Yk3NL1juLo3pXKz02gi8L
VIdawS/ByzW914zMI1pyjveWxAlFg52hCg7MJ9L7GKqvo3YSeCdEYTTu/4m1hCnD
bfQs9xukYOo+i2zJbF5n+ixbFyLgSYAN/EAHN1zzbhh/ILVsE1JhtfHV8FcB98vy
knzb8YxVZcg4k1om/oKKxLiYrffYJdrh6vFibxnTv/6idGcx4nR86lv7qI9VCiIw
IYRW/Qig0wWPr4dhab/kdhSctpU59ktBcnx8W4UjCvd6EPZxaFKtU0F0cRxl3r7B
kCtL6dvbs7+hc2/aVWz+aVgjF7g39dnn8iflTgEUc1P/P9hbWuVGTV7K+B0OrfJN
qjw1OeTfESUgfDEXxX5hG3SlPOi+ik9M4EVk/LFtzKMFV+phMIwv4BMPN/sok3xA
tW81utvDb0qNZj6jrA7Uv4hcxffK5kcOC0mYiA2EKSlaOQFh3qSWQiijBxjEKcfC
vewf1Y9eqlIdyqHCvl33EqRVfYFCN6F/gTdwhu2gPoDOT2pytBbn2S6XrgNEY51G
HkkomTn1fx2Yc0jfoiQHGOIWmd6s91ox368qmS1Ei2uVqcP0aBjJZOPaeesrcE+2
LNeal7G8zSKLCUdkr3fqbgQ8Ulc8IfGcUmzaM+aqh6VQLJ5TNP8LOiiR6fc87iee
HkVbWiC3fqvw4zjLvTS8DBC/NWzRUsDWdG46cEDiPnI55EXzP+aQuRLe+7iSJQup
8eEZLP0ckf/G+OHqVvIpYn1l1l7snBHodgZnkV7RB/jJ4GVyLpfdn8uZAbC4+smx
NJNe1qQS25CkFGhCA5OjMSCkv80BXRmWkHkYL4Zu318w0EJ5eStX0m9bxNce9SsK
mt6cue2fVImolbLEDa5kO6S+tsPiyXHrFqcD04l4jTa42xr4MXe6Ka9+dQVjBZl5
CWhzjJLoJfbEQRJ3DRu1ao2V9CDE0Z0jCeAx8A0wUj3b0ZoU0J9fwH8MWCObWS+9
bZfdFnKXOrCgKdPqewtjue4vOrtfMrRNBtoQQye/dhXaOrfCWeJFztnTJQeblo41
anWbRZXfp76slvfvlQ1bxTA8YrM4Y86Am5CHnA6u2OWl5RQ73x40v08dIaCfRNvM
WemZNjuSy5vmWCqhutRgCyLmyrxYU8OjedTeuMaCDr3hPUcmGbi5AqhUxcmlsb6y
U58219umlLgnvgZ665gez1/2zGOvcEcwmyU5Wn6rXC3isqRcswH3usu9ZBcsN5gc
3CEWVYVStyLsBHFBuv1LOFMaI/zhVArCEzI2f4KH3SSiVLSSnWmW8dbW15yvaAwT
79DvnDNeLR8YGqvdQm974osk58OeBsnEaX2oh5iUNm9AA0Yasz0Ib7VAPTitJ6UW
JpcuDqGoMRaQaw6IKgenehZIV+ljEu0RRkRNtxWoxUrC/WW6yW+hZxLWBzTIWZVC
WCIzInoKX74PlBdJDwGyu3OhLS4AI5yh1b/ywGLotVGaPABX4OLuF7O+qGgBHwU9
pnMeSY/YLVI2TJnzyW7YU0mIDEBnT/1nuQ8E5YkErkxtkH/pJeScCl6kxNiVDEmj
+mfARbOBI3SDkoxXyKgKk8pZQzLRftH98iZSjcYpQ85cN+XU+1qJr4TrZ1cMFzgv
kIYi1WB8iRcGiAX+HEYRIJR0cyop6KeTAvIr5Dl89C42PvcbqreyxxFRlR0UqviL
NnFbIHR82FWbnTmd1xkteZj1SSZAEKMG7kQN+fJK+gSUh6KO+lLUkwMctz/uGaxX
qsNEw6zQq2qoq9ytfRCOOMjYonIl3XlVs5DiCnOhQmZ/O9hFriCGE/GKAs+84sBH
g944Qb9tQ7Xyfk2gueSankhzclod1ITHaVcxOIldbjEZDNEoARGTEI1+4xlAbhen
AKeBSa6OVb2W+71OGwCYlChudOh0msir4Q+Uuq4BLWg8iV+QNDwXgv4CZTEPcVU0
YxZ/x4og/kDW3bLo5mj4nExlRXXN5/XVM3BKuLBjSmiHAbW/ertKwSqLlM2K+9ls
m/7/RLZscv0mILDhV0iTbzhl75lT4w/Yb5f3Oh6EkppHy/GQrHBObtiOJc5cn7bW
RwRnDnlhkCbJ0P9vu6ftu0r+wjwmRPkbkKpnveBBaXS8SrDyvqrPpcQvu88FoGzY
9dIXzDc0yxULFPOshkbpTvUrqAqX8Rg/ZUiJu5+JPwQl3Qe+8LXdb4gWkdE6EL+V
rKQxMSAZ42qsoCcCP2J8uElpNgjVAoBu4x7cJNbruoRT5h9uYuUx8thMK9W9BB1/
Yj3GFEFd0eqERXIcH1IYHxJ/I9378E7aERN6ao8NsB6LitTB8E0nVxJn2Lwe1F4Y
NYdTEefBW6pLVW81zu7BEXSu0IxnMITL43mkRdMkzapZDlYgBus3e6zJHivdy67X
HbNs0sr2rzhus0U8f8YAiUYKTR+MXuv8llQci8ayhl4SGqDHDEonQmK2TTioeN5S
vkWakjqCNCJBTSoYItE5loWJSEZsQkO7K/3l1VrjUOpdyJbmgGYhRm6/zUSFISof
SMR6lEwM8VUIwSKYvcgsLPvR1iP2qzLapBqxdQgFU1J81hneZi0D30u2k1KLl4P+
AXKUq2hLom3y9wTwcif/YkdI6scQ7rzhjDM27WjUJeAiXVZ1bT/m/lWarGK0TobY
a8YyndWP8bonpq/H6j6E3d0S6GMNzU0CLceOKZ4EAjSPmbLAUc79QofamxQrMbIq
eHI00DXF67TQU+harAwv544nZcUQ6IZJSFWRip1b0vI3xkcVsm4C3wAWJNRnEdHc
r/Nlibq+BZssdwTzXdiHi7gBlWgPCYzI8F/rhZ8p1cGyTlwQyrWB5XAmAqNqeAEK
vz/FGubc0loanZRmWQFA9iV+0Da0X+jYI2TY9zGQns8JJRG5qsbniFN4iprKaYMK
VEJFkkWpNH+ezN6plx1r7Z1VVNJbrEjll2unmG7aSB2BOieC+RufZZ9AeVTWfrHM
AMggF4txEiesZ1DXxA3JGKDUvatcdEeAN2x23FKR8siqkag13lqD7ldP8mx9lOrZ
GGWGnK2KzqJngg54D6WHC9+KGO8wSyg6gQuI6iFyUYwsT8JsRcg8upuuPeznEgbV
xj0fMdR99uCMgMr6Dw1vu4XPqVOjPGbJjS2SxHfdjZsYOapw2edl+zeNAQPPMaHj
3Q9o3Dqx4z/XfxOV8IzYSqg1koaajwsh6xDui+qqVLTLApEmzkTQvN/Jrjl6s2yn
N3gKaNi2d2pc3TMlyhWDn7f5WuOGGfUuovb1qFuqQxOqVx/yjIP/7oup90hmh70D
aaAzXaAJWQE3XIFlBEimyHcWzthDVCL7zek/YFMAaTCL2Uj8p595igrFe+0C2UDG
eclExUJYNUb+UTotoihqUkZh72g97B6xawaNktnlDZJyIC2G2nx/div/3X6aBOmB
oV81aFmvCfvvvPCtqRxxcfTxOhqDKEWoGE1GeGds+jY+I3hLgUNaUwWxeGi+yE+g
zsGW9S1W3CIQsLpZC8sTQEHmJvSBmJPsfYTjEZ890FjsDKbD3SfgQEFgyZ/n/l1T
C8+1pC8jxPQce1p90rwk0nbvDVz+CcSt3KPCftee54IQAOesj5l58RJTfoa3wAgw
aAuoDXnMNXcNgin22Q3AdW+Eh8B7WSqlt8jRhlkR2AYM9fWZCMCK3CbUhfr8Je3C
8Zf0mDGrirKKeoq8AQlJU0yXG3acBhZBqfd5ub+yGstYvbmPVZpUW4FnobajD7Ef
jWB0Z0mTHDC/kAv4Wy5amTgJmdlpxL0OXCTmZ58JVN71KYri+oltVJ0lXTPAM6UZ
IdBJmvrBNBQIBMZBcChti0Wi2J+Xi63nF1pJiZtv1y04Bp6GgYLMMn6jBFxcPeiT
OW98qbqACr+VCWD0aOKEWmTH432swnfTpmaeaPkP49xIOS4czgf9fwQ52ucOmUp4
+zlD+oO6vuUxxfdAEKF5bVMpjVj92cSp8ZAC6lX+jebpxu/3IjAj7a8gP1cL8gUq
lpvivBEgO3ulcx/gPaO/NegE67RRQto75+DruRT+DOKBV0J0sC+vx4aPoaCA2Iuo
dWBsl9s89JO8/0mzWGhvmq89Nd8loCYr4B9OlcSg2Ug5IIshqawmHA7Ls3uli2CD
p4aCD1m6+X7hO/9cb2E72bqXtm6/arhoUEMeaIWXTdVIfz98GX6Z5n+kZ46ripT8
KH/ZPBCa8WemgSr0kiqrc0e9/W474YZSWLPPHWFzksfS+76wkg4hofnKI06T0m3f
nqyd3bCKA6y2wdJkBMtwzmQ5duLyBw50MWWF+9FWYkm3+uzma/xkK0daaa+bPIwP
f1A3zWyuCnPtA0TaF3vFsHLn0h1kI6ldQpo1KjdfcyY13ROAA7wVIECviGe/v+8u
FbgZAWS1oGgmC+S4rXiygGmdr+8pVAphgLKyEPTBi/9Fi2LoBIE0iRyMNUZKfXeg
k6pVFmBPevWImr3trF3hkLztM63V2FxcOowTFijLp8o6G5MkuElPDuD4n1glYCF0
mq6ro9dNicIaZopn1kmVUnnW6tjGU11SURlvgxq3fUYXpkxSuSbnhLyfK6K8zafI
DqobND29ype811Tt88zBX7QEwkTqRZiNNRy/iBLDeSNq9ONPiReIABd6kmq0L2Bw
FoGGgC5b7blP+S1ekb0gRRL2a/11JdNmy/QaXMGIfriesVTme5PfO0YMHzjuMSem
jZYLHYkTws2npLEKc4lY4knvdlRMZOyhyKQUhwr+r+DRCQTzrW5TWNUCvYJ0Ro57
tT/Pvd0MhUmrCAZ0mOa21jmHWqBSfwWAGVc9km9+iwhgMN/841Nmgx3C3GpZbtqY
eZlvwqX847556ZqvUeVA0G1tJRV6/3VBbsyAVIPUzfJUwUdxmkkJcpiDoFjCyo2N
cwh7C3opmhY5NNagpxyEt8BvfXkgrbcdHy0D+eYo5J2oMr+kiXGobnlLU0sL7UmN
cNCKHpvfBf/sTQK260JmvUP6vXsql8/qkJhGKymcK/TJLAai/xqmLTGU700ike4q
lLOgl8TornrjPsASSv3MzcssFKyn/VdBquB+dMZRC5j3ZaEyAWnyjvb6DIaYqn85
B9K3FIFIWeKDK1/prCcjeUxnKlwjw+YpgOuEZQTZOluzM+o36IntUdnEVHHqCbuv
mbR7Ua3UhmykSgk88x6L2EaP9knVwoYfaIclv/yrNTjTXtLkX+XNfv5yehU63TdE
7zDPDSm7QdQPiXhBWARbwPg9CRz5Y5E7tvVFlbS35YUnyuYb/7j2b15eP46LIKWs
Gu0k4YCHH4jyZICy5sO+fWv1oP8fIWRg+G1yqvU+7Z0q6R64pJr35OFwlCeMdxRD
vUcsxwdBD00YVxK7IMdpR4XfXUTxApx29+laYmF32ni7Jv2neGquWaYdEwFzA5FJ
qeVaN0MeWZPW5QnLvHV4+jYyV3EFgy/piaBP4zJrST7oeO2U2bPo6VdJmSW7R2wy
jyOcsLWoZMDDKPK4bcbuLHFcbBPCuV/6q1aYTlvBOcule727KTQ21NbgQtUWHKx+
e1F2T/805yJdJz8YIii9PMZFse2zE6gUZgBx1d6F7Nok0qNa979Zw8q8u6Vhd5KQ
JiQu8UH0z01mZH1/Kz54akyoI9X3jSHbmGcIQbVgyx6EZJEGpWTBDHONQOaEHWYB
t6npwTk/lD5wHabLYBmci1vejJsNXUGj0epr5LUAeyF3gbYuHaJLYcg3rbL3Ph1e
E2Z5gxwIhg5oBCxicI2/7t+2ZadqDghtHovVT+JfFCdjPk5vvgY3wHNHrQwYjzQA
FpK43BAi9Ym21ZG2StJY8mioDZYO+XKHu3DbI6Zonng32hRWb1WVSgtD4QXumAE9
F+/Arl5kCCGQz9r7zi7xNzEHEzswMeUYO1BldpqtoHCevMQlYXS6G3j0QWft8c6z
evqSJ477pce0/FUzQhLbfQDXsk4+mVYEfqHg+kmQfqV8K+shuLOzwNg1x7T5Jbne
08PfVH6NKeQAoWb5zWHk0bec53wmH/AOfSUTvZVmzjZ9MHr4tfZZly5hlB9jIM/c
9rQfGw2I+J87hUTElL0NIevAysKRu1J6yuv3iTS1Ai0ZAspXcC+Ltk4wsqRihQha
wCZXnKAGY1XrlbZ3624MnDgg8EuwbiL+sHlWw4tSV71H56vTpvJQ6KHDskPb45Vl
4jYjCwwnlBd3Kk7BGhPMCWQYZBrVNJY0yVlVePepA0onWU0MeiLBENY2zuoJTyi+
VZZE8GhRGn0o1AwkGz4MHDiyTNJXH2rIAZY2PmT+BT8MR/i6aC3zHGfskz1qd+dM
R5ZetmYSjvKyvo0Hc3+4HobB7UUfbu86QamdpRB92lmomAwe87iQcCC3Rt7bdlpU
x4cF8w6J2H8qprEI9qqpoLWr+qCO9SF5jLcLq4b5EBsn3MuPl7NUueqYMLxH0ctH
72KDeNq1SiALp7cvnLRc+WrqPlBnH2ITWBISMtbtXVfEgWChZX+GZHLR/TgWG4Tr
z2Ar50OU5XUgnGSMO0hJhtDOcd9uWgqm5kwwEAJbbyLbc7B+AybQmSW2Xsebq79y
PyeStK8sMHtkPyU5PAQ1xSpjMw4qb+o9d2lXBeLbdEJnr8WUCuV+B/JlDFTBpAtB
Lf14/oatYdxnXgStHZBhw9bq/HpKEgOq+1IWH6ZzS0WHCHfjoKNwh+Km/P8CZcff
B5mn/mSDceI3KNgvxpz5AgbFso5IJmX4EM/YVYsWnOwO2ywCMVbSVfMhzRjzAwJj
O0B0VFFp0H3Q/OHmR22/Xw0b7RwsNNQqY0HjozIVDwzQGqQzNryHIIpt9yb5jWxo
pstvCct7mRHqLnvhVy5hgiAPZjL1mtpAEydlqdg9/HuXtwUrCe+CL/DC4+c28EEe
XlxvLgMrXnGMxUyx9ubhQrrnmq17wviKYj1kdQT+xRcOt8z0F0ETJs4A4Qs1SqJE
BHwzlbHcHiq3KLqjsxdierFxMdGeHj7GquH3HhJIk8x8+lhI6thYlTT9hZV8Yn/a
rBpOqmBXEi6xFnrNX4oNQt0dx/X7DcyegeIGtI2TtBjW081NRkgWhoadav9E5kiV
9iyl0ztzbW3OAT1nm6VpZT6X16A2zNpB43OGYrAFJrWexHhsU92qzX2Hf/3D2EwQ
hOmqiuOIlU/RE2jtQ32qvalQYiQJ88XUNN4QD+vmFAQ0wJccpv5stPFk20/rw1E/
uvbyloCmSM+7qMDQFTFu0ysuGhkeLF9BKMuM2iXmItn/0X/Ys3Dhh2SBXLjd9vMU
xIe8S2NscH2szekOVLD8RrGI+cb5lbJsP/bkvYANdMRH1gBHUjLfrFZtlGe4/lFp
JOtE5vis4RiSrHnly0xDJaLtiwxhiqnd0mF7nm8kb0rrp87lQ2YiNvTktof8Uh16
pihvaK3LuW0s4W8kl4GrJ7g00RJPQ6D2R3F0Y/FP0EjxRlMPuBLhOajp7CReL/u1
NPtiI0V7PNFV5ACax4qAH0aiOU2mqj1Ga029uOktrETxh4d4zVlL79p1vTaZjaE9
PwCDQt2EdGH2cbB5bzenP/gfBRX/Q0eGDl0ohgDbjFZEua/6de86caYXh3S+DZfy
Q7fVh8xfRQ0aTcCJChe5bvOk3O6QACGh243OnoIp5gBS2LZV4/TP5zOR+l1qpdSm
I2LFSp8Z69YgjyhyV8fX1h3q0g5ryEC8rTBzDFprxE/zoygk+06n/Q8xGyJJshRf
BoQmKmgZK0vLMUg5o3N/yEHJJfKm6crSt1JoZgEtnDb5Qxi9Ejtd1LEuKC3gtqLn
V8q/OnVgNDPI07Zze69QdXZB+QdohqZr05XlNkgBp/sV1//HiSWpY6Fl4hX4De9D
pH7sSe8mfTSB7bvr5nd4ZtvuUkvist8QLWP8vc5VnihHZPXI3okPNMi6tPVkp3qV
Xa7X3c6AIs4SJKZOPBknyooHhupnNro5+h8dqhcVCVKRRH+RfOKwAyBmDVoKZO6n
5oBTN5IUTqbvpu7A0en70NsN4b9CFYE8flctu7fynv4qxuoUsud4ao8msifAZSxd
G3c9+wk02LxwTicwWiWllDRunih1PDFNVFglYAOoB2D975MhkXH/pToIRk1uWkaO
79X6Rzm7Yzj6diX00mbSvqfi3vSxLFH/xkeb0+W4+t5fOCk3FK4Mq53afhe+tmgo
xl2EUs+D30cfM84rChZ9imkKVNTho9zr7SBiLU+Wk4jkshzN/t5jSlVdLkKv7S9T
m8W4sjgPfQh/ST6yNlOVx6HIjdoghpO36qRT0T6HgKNx+ynG4u7e9IZqGRwb5hT0
HqaxfLvi1UqVMr0rJ4pN0wYvoY8lWAtDfnkAGSuoSn0y5VunRkrBkrWhpPCbTtks
tRFYmKyqHwm9nDgPeddKGnrKSq4Lz5nANAY3yiFizDc+3Rd8ieAtRumA0C0RSPOd
8xPt0jKdtnx4vJ1tbhAuKrDS9QyildOQokg7+L1IIftyffpFUQWf8vW9d7yexLcG
DMgxdj7flTSijvfdbEljt0GWnqwcS1GnDv/+Gy/QgtJIxlszzZPPfi8kS2M6idIu
JUumDqmR66SvGgyD8jZB6xfePRGLX9qlpJlKLVkyLsSuA1VDenvDDk7eO5Pcdw52
kjbLtbhMcjz6N43KTypVktH3rlnOiwhAtPcKt7BXYtwa8ts+smR2H/MJazfrNoJG
UlvDFpnIiFzuPqeeATXelYsQi1Hv11pXr3iiVBmy66B60tAzqbKr+cyP1VT6IyhV
+iZgIkmnkgk2JY96h7oj6RR5Ad5YHKRettupxaJqYzY3l+7XcDHtYu6w3lziapcL
VZgjejTN6Y5Qft7G6kAbkuGBiXr1MFlFvDvh6AvoLDojKIulzHanllRdtmRWYOpR
/fRCWCoxMjC/Lajk6lAXD+h9gfNx2jfeVH9GYAixvtiPPXhykN1XuDiLI3AmDkAF
btbv/NBqvSE2SK7MczQSVf/4dQgyZ1aa+AMQbmtU/tn3dpixZwWEAOqjfk2K4mee
4G+NJp2FwtSktX/Zcr2U29vFDlmmf8lL3Z0HZcWyFIXZnnjhfiu/O0dha387oGS/
x4fPcNePIb8yBHKZI2g8WyUmxdf85YayMiWk2XbWAwMT+J6S2B0uUEj9weKkw/N9
QdWChoNHp4aBYi9f4DBsm9LQXVhpgoRuAokXRANdZgDOw9SBOXk1scODL51+t2XE
gfL28nlGSuX1epAiuJ9P8/dcZcXcOYjDiobNd7+HQayN91+DfTzY2iXr5LIj/Cyb
M0iRcqARqn4gXXBrO+IaM0HoxgMgT/XQO3K1Sry/oxN5OP41ByylULFVpvWD3WcW
maDfY38ImUzqDzbgXI7Q6wV8KL04CyoV8JWaQIChB+lqLNJmo9I+01QSx+VYc1mo
x3gezxnPDp5Qqf/uBwZfImjNo+/dS+K6wR5r3T23RfbaaUOWGBbyutwWYcDuVpQW
+OltWBnLHS+aTfZpKAEVfIywmklkNxSOayTohYpybYIeNSaiYS/UKhZ09+/cd+a7
gHaeptuL6qfLUIaLopYs7BGfMcgG8k6YOfQGYal3O8yRXlE62/Nw+nPvzCwJVCYW
2T4PqpT2hUcVGIO6S+g95mL623snIYZfzLixVyD7I4mvRpnGgLkBhYmYCUFOa5hQ
BtfETL6mvkzcmhTU4jYQh69HWxKUjeDtiPvNqgEBpvQNH0pVDgOa62TD7xJR1hSb
G35MV/IlTG4u9TSFz8GKOSC4B5J2q50RiJzPzgEaAGd4O778Vz4gQFFyXeT7Z+i7
C+GxuajZot5eMBq8NfUdwuYFQE4mGTB0XaQc4ZjCuFfH0yzfQdCzrkkU8TRgw0Rp
BwpG3AUDfTqyUVF4zbuVTPkKHogDaUep1nHyJeqGow7JOAGPOmRyl7miLAOMBDoO
8gCPZuFe2WnKiLY3bl5Vf/Ixr3q6lXlhCzgD7yk8Db6Eb/09l6lO7h8jOaCo9cGo
KYWHZ6q6Z8/WFDDTDss6SiLGFH+HFXOMWkgZSR7k+24bX7jRX7jezkr1SEnZN2B3
ADnMEc2vUcL21Fld9hFbHzCKGKRCPLF0mySwkjKQ0bAE/HtfriUf39vOAXRPmhqw
yKjliTlxUOKJ8BmSydWv7XACcdwVRCr1lIGhORw07o3T+CHabT7RAa/7sfxz0ITx
+R706BGROMEqjad0Ycoa6EBVCE4A0+9K26WDVRF2Yzy2NNRjVDodRFru0DEH7V/T
8luSNVKec9NwlFxQe3c8mABJGy1D+1r4NI5v6BCsFc+TeiORjyoVXUjocN4gqWH3
/njBF4hVlh6uPG7gesGLUAqSabRASrPmLbAiCTKfXCNIRTdBgcXNkASyeQGHEABZ
9tOuIWR6rcli694KgZMGQBYTAU6lsbbGgQrZ+2UGJJDTOenz3Z49qrzXXUDc5HVd
EU3y6aRdPpga0siGeRfLga3eszEoUh3BlGOfsvSt/8CI4bv8usEfhvksOWtPV7LW
fZNmxoMYffFPRrtzVE2u0H9oVU5RbBeTXRrWuGXsBve7OKS/6wNOI521qRis7Jp6
aU7uppwT5wc/uxv9F6zcO12N6JRBb54Ve1ertVo7mdYiokL0FCZvGHB3xbw6zLg0
IvsdAGtFB4qHN/Crb7hnYMdVs1ZePb+I4aClAfmci261NEXP+iAAGLn6K7XPWc+C
pY9KjY7P8QRGCpU3eZz7+PWDl6if++9XDolgWocOzrnnRv/i14mOMla+R6oIoZ6f
73F/31fYql07yiX9C60njRdCk+pRtPjhzMyw3hfaDCmdSDKBYXR9+YoUtBUjTieM
RWE61N3MDsn3o7f8eRjkli6J5OT/fKZRJOtw5BHGogbetzzpDOFXQpBfznh0rEIX
Go3/morWpQl3XIshvKokUK5mysTsouh1/BpRTolXkceGmkVCZcJ7qZcq8EKTv2Qf
MBQkOV+B/O4LtkwyU8UKTZU9SxLFV2T9J8Sc/nA0FsdAxFgkehoMbobBH5ivREJe
oCkaYpxviAdyw9dg+yR1hc0bio7PBOkJ2/2PP6jl+yV4HgauBJUYDaWB2n1A70VQ
Ftw+Ds/q4+rEJ6Rvg8j7aA5wIjHQ95/ZZ2PEawbLy0Ee6kpnSJhzYoG7zARwYm35
wYyyCV+Yuaaign8uU5TiHCwJDdll0cdN09r/gBl1fDMl0xY/eEOaEgh99oncJHiz
pCZwnRv9OqqorNFzZTbN/YZJDxlguAFlR5yMFtVxZYReSskzISxnFVj45SSqsBcl
ctmTzhWSHLtoZmr0t4pgjX7EV9PaIToBSqpEQCuAQKtmOJtQVXhaSIe1FN92qOsx
c9/LrHijae9gk54OqKIKlgfEApyj2feKNq+sJtIsuA1t5B2iluhrEPl4y5t52s8W
h8bMBF27H/GVHGkQwRQssH1kuMfYqKg/EuhRUhktEEZn52pq3F1oi8j+J112aagf
XV9ethh7ynU3d6fD5ixM6Q0/6JI7XmvFyWq24AWFRP6d0YtQglwbVLV62Q1ieip5
vBpecYXusuc+OqmPb0TGCJ6974DO5yULngh45dS+SrjeXNiY0xpHRTSMk3BdIZsD
TT2XC4Wsdz62biSr2jULpp2XYpQZDTU68TnFfnugQM9c/VyeN/RKTER17ZYE6kR9
2gBtAcb5vEatJ4Qit3injVA2E14u39OBfQSG39EWBCS0SGj5/KNylh+RcahstiGO
9Ps1LMglmLw94YNpH2Lh5Lq5ARMG/bRRsgaslPcZv4CbJ22eva223UrlWDc34KJg
KlnGpwAJRR50Jd8AJdvyKOb1APCRRoaKGhnLE+Z07ntIGLynALZbJfNQI52rGM+c
WYhFKa5dc2ONG7m2cHM7sbH2qDPO4jXgwSCO+9KGmYfbdNEOz5BOcg2ON8iUq42N
WeHjNXf5JqmBb1krSq6HQ6/J2dA14H136rrwyzNw7EBqVt5DzKCCxThKeWmttUuj
hLsIbskfBbuUKd8wDs6md3NnwtilP9fD9ej2IN07npXcjHj6spWMeb57lluIb1bD
gOqz64zXY4b9GVZLTfnO04EuaSBhjiot++FsXrtiYS8gxSOC/VKUr4Mdb55wQDiW
GO/3l0Ex6dwJCjyIT4d3ur+QhpObo7Insj9pgugihrVqrqniPo1GLLl9ItpsijR6
S9j8+UNRSTAqdOU3XhBxD51JozuEof32wtzaSOEvmKUM1aQTuyaiPmQRnITSNXv1
EL2CTpdmflDmkvFMcraTJuNZbjj1H20ibfJXFCzTiYg0Ke2enC4WWHF8D/HSDNZp
IcUA4l0+Fsh2bqhRLG+KkwHea1B6DZqrJL1skRCb5ehZQ7JqdLE5GSIjhJLoasez
eSExQ9LJGtzND7TJD1NrGoifN6nXCxfNYaG1c/Vg+jguooFGZhVXj7pUzGe8m74D
+Va57XqpuP579x4O7UHxDIE9r5w9JCkTpr9f3au3rSYcjC0jkIpWEiLXo4bthQEC
E+xQN/2UmRPqkzOUz24xdjlK0LkA9huQ00geaHgC6LgHgLVNl87vWFxgHeHNf3Gn
GpGC/qlI/Fkla9cBUoAZ6ce2VFmmdY8X/LVrsKhu0wITNRFRqEA8FO6wok5WhDdr
0DP8asF3tukN7BF0M8cyHxDET4MKtLYSpT7iAoEunYj3/YlRxvYA2QcgyVfOE2AB
RjBZLXbCWzmF9YwfQIcMiRgOdHsYMfPEd9tbTr8ulTGlK7WKzL7uUzMoTLgnOYVP
/94qYGG395iRi0vbfVSBtAxF8Cl9fG8AGLqka/O1ABThIqkKRi61N7W8kv0lhC+1
45h/VpBsAa/80bROvgbbGJH3RzMSle46Erkyyv2CbbBd1z2WodVBrr7CVCTTgmyq
KHjDfuALhPjgY8JV0BPyv0QwBzN4cK6n2JiNHQGWsdiCalO9SPj5eF0llmhkiyck
dhdjf9k8AqsxBymx70TlhslHf+ZW8uweLv4W/vPjTCmtUtsJ7S6Ms1P9tsjXNOl1
aDS96N/t1yGK+qjLgTZ2fUjgzpOH9U7d8dME8TH8yccq31DZPXIFqwy0YS76OjE0
/PeGhWSudBIn7zLw8o1X6fpmDYvUtmmmH1NWeqrWl8o8y/R7m5nZcqtt4ZB6XtIy
PGlTx8OkqV86rEO6Ctq6FEky8itxm9WolBTBpJxXMYqtAQCKkZOuhFwiOObd4BUq
D3TXFHB2utirVeHtpmRmZYRvZt17j3o/FP2QCAa4a41UmZ0799Qluu7gFvHTyBu6
pmZTC0NItdWJkbuHFqn9WJlQCw/WDIZn4x5fpIwaOd2xnKjh57gbFoN4e7FByElU
Nb+AlVqWhtEIlUG+EjuHWYAs6IiQVlzH8Yt20MVTdd1JJRgqnzr0Czh3CNneFfD2
InavxfS7IChxmaVS61+cVmuxWSQfc6m6sQZkA6W3CALEx8EnwF4cv5N2juXTfzEd
gBZRRG6jIbiM1N9rQLh79oWD6xrIHCSL2QF2Harin79RJLTIEw520XozWE8kTYuX
0r0FzwL74vCEty8Z6A9OY2jGLBlT5ZCAHih3qr/OAiex2ZNoZ/zY4i4o6y+tWf1s
bsSaH+6b8KODkvukRpXggrvSuYfiSfsSiOqwjpKbOUfM+7L5287ejmRJGhI+9GhV
9DqlW3EiB5CMSVvPgpvWUV+ku73y3V1UicTVoV2R4K/Bwc6tNtn8MIYu6BnTwUMq
Skl9XvT+rZpEacJcHEN9qce2G3B/r5E2ngquL/EQ9SeHFp+4K8ULAANaaSyOGbuX
XgplAiGxdV+WbUdYCcF4+6Flkh+kE71HbpVIwAK3iFfWbGQENOY2ry9EJ8a5NmLs
trAVlEZJxHtYsssE54gWb1IMTUjjuIK/HWd9zCVsElI4ADF9NH0KJU1+lA8Gvi6o
DzSa0JtTjlQUh+fHg2kmdcVIW+wlrBx5pGh50ZqT7REInWmEqxFTyfWFraZz6Dwp
KK5o9EUco3AWhjQwx8wQKxgfEqB603zAvW6G6NGj2/ez+b76mfOf1girMyRR2eZA
3rrXw5zJRvjL5Xe5R2xEzF4n4d/WxQQl5rqT8fjdFJ64bB4wYFlutl3UYtiGooGm
h3gB+yxwuaBLOWZ/A8mIr+0ovisLLsexuq+udFDygfg39WmMyIYDV9aah/fY8lFv
FVyvI8ICsqD+PRKHZvZ/kSUSiUwELoUvWa5vZGkIrd7sBaIwoOHBJml+bc0qQhNZ
5E9QlV/jA4CGqGE4NKz+Y4Cr7woSMfRooV9rZBWrQPMK7z35Gr0Hcpwl9PEAxaRt
QTxg0MMaPFqk44HaqJ1Av4ibPekqOnr1XIxcczsfYwLt+TaajqxjO+ldpX1GjStU
/55bjO/1XI0FL6XWLRCBPyCz8mapuCIuNX1JxhtY3vlJC6gf3ltagy3EB1z+MYDM
tOz48Fo7l9iAGq1s/5rzwaLQ1AEYiaMl6n0Xap23QTbaJpQJnOIfer9IaPczcvGT
nqFPP373xf8yYd9HS/buH3hPFdIwUzmCEUZMbltSfLHEXXNTdq0Jhzo1yKPVEejL
iyZ2P58gHaqQXSa7eZHs5vBCHQcsAI+gU+pS5YI9DwCaY4mqrR7SAeChSz71MPWi
XkrbiS9qZDyBkUaKNvPPW2qYqnaTwdbXnmMyH4eHDb+jOsYUi/Ds3brn31NuK7HE
L3buDuAmQ+WZaKG47W0SqCPWFhTfmywFc7V14dFviHgHesPTdUgSOMTasrYrOHPL
sFM5IdCzO4vCIh053QrGa7Rgii/eKByJ9spAHstKbll8b91LyXmQ8o9q/ZMI2log
uPyqiFtjH2RDKcX9XqpRvAm805ca5/1Z6kMXwbJ0Env7iTJkhTqYfOxLKsDd+FB5
udVASX17uLhyirXvm8yoKUH1ieqqPIGqbLtrVJPabz6F94QTFYvdIdqJxFBJ/IQL
25zJYL4M/tRkRQaHuz+en/1spnE4U3jdIEyA00se6Bzag5BbkC7z6Qi6Zq5rMSls
1zOdlh5VH6CUrjZzVFQEx3KV9EpbPcswxgEF+ywY2jho88NYMutrq7SicUTrLrgc
fj3HhbvMp3wL8IP3Onx0fIAgmZVgUaQSuz135ljhHhwmCn3me0riM24SrdNOrp/r
O4U3dGqOfcLxYki70IZvKOZxdA13iqsKpYsODFXI8WyQvGCfINZwuVAa37K6ZTRo
N0Ewl2LeowxgjWoRmtD/FaZgww2l1SuP9ThaeGFyPoNLJxyI0zeDSTNWrE0LpkrE
EYVMwe0jX+F73zfx8chuJgA9nW/NGoIl20HkzU+99TUOiJ0j1pzxrCNTcYU/9dl4
tbHR4rWlOlRFwiTGRZ+hatFhkC5MWGN67x5WaH8EaJbYdtvv95rE/XTC+OyFdrxA
td1YtM5JBsZk8BB3kJhlnj5riS38dBU0iftuxAZIU919H0IjBVewT+maT1gCVGlb
VpdecWnYmSrP8mFtQ589Qi+lYXhJtVM8+WsAE+XHxgTO7DtkZngqJ7btnc6UWSnX
meqyt4e4uVIfOxK0QIAo8mlNXxgtfCDvkJcLA8qJpr0MM+dM5w2uovANxp4MDLEp
yXLDt8KUr+xmbyReRT8rHo/774Hgq0gAuAvaXMzcAsFzaHntR1FMrtFA8E/juJdn
zK7STyYc+tAXo51bkCD0eHiFNy1cqvaLG+UDOHXnTQ1beaSkycDX7JnB16wksXhR
yTv480YhP2g3pex1Y543m47p29DRr4MyjDBnCxv8Yy/H5R9AgTDtZ3qlY1jLcWs+
zyXZBHI9GDOB2SFEujd6PGqEWRuR6PqgoGYOuiXIxXXgCBb2i21A3cq7T5X9jEdG
kTWuEpZ8ttzu8dPmORuh/ztCntE5qYU2vMIUefOiqeX8D+gCN70hinWvhWkcU/Mn
KIeGvqQ2cIVxQn4D1GMS+X0yvV89CgZ3M3peFHPZ1DaiQ1Fk6Zjh9IPAxJk0iYCP
Q7pQ+VZiokFBkEJwUiEDJfB5RwWwf7ceKQuqh48+KjtDd5D7O3VjehWbKqVuun4m
PlMqxy+fC4WU7+glvamFKxN9mtOcyTEba67U1dlLnHegfhkFAjkpqK6EhpyoVoEN
esl1SBPFYYRP0mLARINxU3YMHWYAJx4lZtYyXqXku4Fgh6IDKzaYAI5iKeEWFPc9
QveQpUqq7TqlyR5fjIh36fAmPk3D60ZA8hemiQ6E4FKNdyJyL3DujuvZVGmHuDsH
0jH2jeoah+5vL4ocX1bn3bpabwIBT/fOEJ0cZAssdbNCYdLZQneroySDKysiVEFf
nlwaJ9l6IL/ciFwbnZDxQX2abIs5m29pMp60JAYG0NhHNQfcxRxJCbqMqFTDUK37
Zyyioo6BxTyFOm7tQma/QLF/HYnapXhMNth2GtCt/XtIBGEWJlqWz164F+A2lTXs
n3o3UOIY2B2vZcwZ8K+DXANcZ/VtOCERC7XRY4KDLjBi6OQDK6w/QkL9LYWK859P
6/kexFebb5dvxZyOuVX07bkaBwBDibuRIsgAEIzV2BZRDLNoGSrRJiRNFQov9721
CGQWLDBDFV4ZRDAFB9/FpcWdfvMgeaLU/68ptPQ0R6t8N/pj80ADPfavLWGW4ca2
bPCwV3I+S33uZDWUahmvqkUTAgKX+BjM03kCHu3JT+vlU+KnWlsdktJ/uJgUnMmT
522oT3bXpsHJzdNjCAWsEUlPesVAHsFwY2kYWwCP3s2Kr7H5a1Xo9h3QOvUGY+AU
GH5DDFzsJh7un+U2vev9NbJEDPloxd/hwvAow6IGin6HMWud1v/MYuPghtSqev57
qyBr5dZvgy7xYgTSFhJ7LFu23A2/7ze+20x0Wwf23uC+IwTM6KwUFpM4I8N7/cCf
18gKgCuiEc9v3dlTmvUHtjhMBOKJU6NVAsLR4t6XIdQHFptErkcv6dduVxS8BJQt
70dABD1J5lt5lesQS5ylOZR8imFfnPdk+Hihz6zerAQjRxavuIVqNVaJsf8xVtvp
pe2C71Afawz1A0jneLPwXvPJpjzwmZnIzGW9vjB7AefmjQ5XvOexKvxU9nHm5g6i
HPwdl9u1zQO6TXO1UbQjGjHHezrLHfnBYflLsOM56vOcXxVTlHJ0Re15RmhCbGeb
7cEBEREVUWxYjgfYQIa2FF4iwp6v/NOudL3PuW/l/kSsSCY0v+IEXW2FkKgcZkbb
xC4Mt7gdq/sdlKqHxJjVcBGBfPKOWC7D1tSK2J9HE87fAsVVyWT1wgdTQTPkPbmt
BuP4+UyiWXroztZTOlrrp2SDtd7Pqriv3LswADuUUy0G2IePjdsjssAm4x6MQo8a
BBaA0hCneqx86GecOIssCNmkG8n/T4S7jh0SSCJJFlJ0jPmeEKenHhpyHcOZk86X
4Sjp2VNLNarVXdQqWky7GTwMtxX4rTZTMT/AOtdbvCFy6ZPXBJBPXYHcUmiFu8Vo
iJBBtIj2ABMZsdKYZ44Yt46uw8061EAX0WNvP0h6W5jTKRRTGp+i8xnI5IYNhmFJ
WaJl7xqEiGl/G0gVfYXDoQsA2jVLjZAq/Z0eA26Xd10hvej9l2Qdv/+zxZzZTM//
cyD7qIg8TaZvMiI0O9x10NQCBJPicva60suUfUr6kI3Rdk8u33Ny+rWV8faMcYC3
oRdzq3aS2qDjCI3KN3W80qxE0NcPqqyrV3vfuxfyOOI6vha9R4OJL8FSQiEfu6oj
ctCkWyYzFlXGR+T1gPhi++h9pmP1axvvr9XGdcPs3GpJxgGWNndP57XVobopRyPk
IMo0EY0c+pSLiwM0a97+OLyFRbUgulv/x14d9L/JDk6Sn5bvWyB+VGA6tDqHv4eR
RudRjxDmEWPd6wXimk+q66UbYSBoGYPgVaDAI7k2wbjc47CO16z/ACSTMjRYgq4m
LYaHJhFJhiBdJ/9p4JpguCWmLo+Yfp4x5RCBYypJ4daRJn+aMVFviJbFx0h66oUc
+hn1fFPxbdDAVMy+EsuLMKExv4JuBWenxbVVSSQ2QwvYo6pqWun8Ovbla/QP0qzb
WvVQcouOeFU4MI9MVo+uTE2DNAFIwIKGsHMO8rNqnWVtz0Mt0mfHCBGR31zYzpdA
fzVGAGLeHV1tyl/6lspPSDZvXNky1YDvfbadgNBFuf9zKkVruGV1Wyc/m6Y+2g/9
8jx/KBHVATlGUZ8pZu7B5k0IJNwJiJPlRX8pspM9pH0kBjdmBfjutVPLCrnl8Tsf
MC9Qyp2Lm9uEyL3sfQY9VoCIe6L2MUyDtW+0KES3YmY+IQXINdt1TvRH3HDAPd89
mYdBNOYdnDMAKDWXw9KO8/dkf+9BJI5qNvkDMBAoPE98eMQ8lgjRqCdLiK0S+BBu
fhV/IT1jc2y+/FDa6n+EjW27ugumxy0LZXNeUo0tG9qwJss/butQFsuhTQUhDH3B
m7O2ZKRauBEOOabj7E4sV/JGR/aFK5bdHDvTLPqjLBZbt+RGDNJwi4gTWg9M7SWd
KeM7SGfvwsCAJnD/VBKQQrghFeZu/OqWv9K1AKpfdBUKZQa/NE8zXDZEVgxdUlpP
LZ377dTxOI4TCox3BeKBEvg5CYl8j6hZCTDIAu23yohpErWf3xgqDymqY4DmMsVX
60Ft02ixMn3o0e4xGLQyj7h4bibcuxxYuMZlRWu7tSG8m4uypRjL8ZbHHPE4f0KM
RXvV/hKcbrwFTmtFFosH1rVFiD7R1y80dArBJVYFbShFR2+/m0ZBiQDJa3JWr+Xh
fxebZXSN2WnUXinch6RiDus2zK+7PnIIZ9rpA0Ft/N0xSYFUYRZvs9ljTQNeuMOM
dJYrQu7hXzOnFwpNa7tGGXa3PY/GAveJYLMZ+vEGL94kih4ERBbOlHcUxC7cJctu
z36E8sPwalMIP+quPO5VgaGjsMPwAExneIxeqi4mXY+UkjX4BC8HGvMOpOwNdWhC
PFWQIEgDq79wD3L/WZw7HB0ZlbpVWelFW3PcmHs8fXdsS0CW1+egUSYOBGojhvXG
1fDjOFd8PwP+UxhRWj1Cm/T92rXNwvRSifS5TEpSQ0o9UE44RayPqdMxk17wDOHR
SEFtXj+51NpC7L3xGWIn9D3mzZbdoeYwMbgsJ484Sj1ZV/RM4qOiRBeg8CRWQgdM
Ef8On4PqldaB8A6cOXmyLUmFWL5LAQ8JXIkcapy1byZ3lqsneNLcqdAyBZ2uPP4Y
Xl/9MFBjwK2WY0vaPBICD1IUlJKxOYJfTw4e0xrvU3dzOjqnlb0sXGOBHfXFh4Sw
/dt1jeZ2l9Eg6q8MfWxJTXvv2/6Dz6L39Z67xHnCEjHSRP/xDMdKgW4gd0RYGUK0
CA1u1hv/bQrVRoKVpNwrvq1u9l2F3QlGk2zBCqPH/5FSBIPlrjkEwkTm9IcfkeUH
6Qjf3K+wNx6nGuTok9fjRq7k1TLrtcpSVqhZzYxPjfDXmOCoMOwiD1np5yHu9aVG
y166aNuiGawuD2nI6ouFmf2syEjl/XX5WE6+l2ChvWxFWkv5/rVzuzfphCGRfPXu
8R9fltQUnc5yGia+za4of42gc37a+V4lURGsrVU6Yo8pzqU1oaAEPJxYdjugZmVe
dwDydfENahjXG/kHRGdcayxemjLCjjQIDNDJWNJHn73QvH0mWM4H2UeB6wgix9Xu
mcZ3CvHdr5sKTPeip48MEOwPkOqcOgpYWk98IlKywUnkYYpN1ZXJDTOjgiSTbFfC
d1mamXfPWRj3G77wplHGRyl9AOjP9FlYKnXm73HX1GABPPtApggUChhnJtw7b321
Hzfiqi56bM3zC95CVKcsQHkF25Hya6RE/QbglRAVbWhewUugEpPoXStq9Ig4WgAl
PI5eK5U73z4deK55/Sn9KL6dSacBLqGtc4WfquZl+xUjr1151YzsP97/99bfDbUw
N/0/UGDI5oL47+0FMBggAZc6HdShp+05Ew+MSRNyQm21NtVOHx3yPFd/pG4NpY+W
OtUrC+6WJSxa9a4slXvFgP6FYrdwVHRGOtFjPIY3yb/k4tldxrgkk4iWjysddAMA
0XXOfc1m9DKLkenAs5vom526mZ9KYXx4BPoxcg7EAmIFr+hIQXN2Q5no14zJt5QZ
up4hSLst25WzniHeGLkuVI8hUcPIoUqpikLQRXtVEmSR1AFRcmY4tplNLPNmVRZM
hd22RJDfWOqi2ej2lw5JUviCnSuLp516QrDCtvXaI/gFgQm5y+kU4BQqCPsQu7MW
2m7f0QpG1YZh8m6EpWTFX3zlIT4cbPuWEUdumOxchs1cgvlnyDLcV/56JYKX51zx
TuTA4xM34sqJkkxlvyyWd9cuuoJQ7knIe0SEsYY0lceupJreiGis9YO5WRafT61E
nC4ChZpFy9F9Xb9+obguDO8kDxMnjRbAf/UZoQnu3VRU1ijQON706wYCF+iHWaiv
Xw7CwgaVoS+ymsa0iQPLFvb6yp3eHXWCpc7svs6d4MukKJNXo52JJ0fSwXPGibCm
lsmwm9orjwTiuQHAyCRl41tkXyRyw1N66Wzkyts4s1aIPrGnjccfUn2RJksgLLT1
VxUGbbvKRlRzm2WK/ejpzD+HYrhNhYiTPksakUWiiqPtsqANuINXzpXkYY5KCqP1
U2E2h7qA2CKNdV6ZZbQS7+LvnmNNbGsro/1H/iRvrifgpRtjiwy/rL+Lhk3bBah1
OJfYLVgRz+qkjqI27je5MgQ/md8DrwtSEbUQZ/soadzwAMY0SJilKb0kv1hT2L7f
KXHRI9ro/7XRGUogvAb0GQtErcTEvy/8N7gAd7JUS8aUtkAP3SabcYTy+lHxmYsf
hLXWA59H7AzN/GlFtk73DzUDHZrK8vpiozhu39sWNDDy+CPkh1np0pKmXQCa1UYY
6aGAPCVv1933L5dt+xIgreSqxJO5zq6Bs36EXJxPis9zDGtvLHyY5LBeXf4wD8fz
KriE0z8Huu9Y07jGggBw9DiPzmo+qkHrHZD0l7zEt72Vki1YteZnVK9pF6oYo/2U
dbMAXDQGBatMsPOhY6w42rDDW7W8K9WCTH7yI3Ike0QTHRLNTWBhDYaGg0bqNxvF
il4X8zJ/Ip9uc5HJ8C5YggUlrLq7+mJ4bZ1W5lpFfb6fqAa5/LIo+mrMKTfUYcPW
/8FdgephG6Jqu2uQWt4JU8jJZGZTzkua0XsVhJm8StPgTFCexSLGUHNdtO0Iz1QP
XBla7Ic2Ve088lcs5ZdKtXAubZ4QRdedkJlrntj9jHSd1jQsunKE5wTgGlt6H594
FNi12ji3XvqKPEakm1IomxJN878+zoUMSv5RNdF5eAMWVYZI5Ptuph2DEyKj0Wjl
yImd4q8/P6fs42EYT0xisOG7n4wl/EQb2Qy0Nd5wtlq7FI6fMrgoCtLITGBQ3DA5
HHh92PhJVp126E34XYeYxCzgHiiYBTnJ1cXmJyhlUbZ4Cq9xnthNHDd4DHe88Fwm
3wRo9pdMN8UlvbSwTo79agBdXSMPfmqU5iVatRNhAxLrlC+xn6rWh6B08j3lvHxs
oDMny6b17g2g5o6+XDw4IO7GLtTYetNWCf+/jS5Lc+SQhJQ1GdH2zSmuDw9Cht9B
tkExbboT8DyelwE60o159N7hCXQYLnsWzRiQSsU8uEU1FSXrhvXjbaLSFHCiqqRd
JQlUn2T4xl7oVvbNpQ2+iO5fztza9Ij/iSJPURueYemkJdP6JumrZktpFLhkakbO
qaxrOBjK/Cg9U1iaxp9hls/p0mX+3bInqBX9pF03pRgAd9o3AGQ27IGy454uIx3h
l/qzT3ERMbF2l9aV08G+dH8ROEuB33l958jZMFeahvCRoXSNvMk1A3mnEM6l4iyz
5bvktUVpaPhXHLbmjxI5rk5MeYDX4o2k+mgls/k7taB9gaFSjtF7nE3YlV3+Hk/R
xp94rbbeqvWY0QB7n5XX1t31Rxi2R/t2Kwz1e4cAxbVkV/WpTlYm0HIAajHOGak7
KWrp0Frb1KHZpCKtMyY6HX4OpbtRejNdxB4+yvkS4A0zL4DmAY37iKK53r5dQh4e
7vbJa9VXGzkoJoww200I2LzuODybGU9tba/Ll3ex3UWTf5ZL5GwYKDmIDb2DtIIE
514AuXNsgejNb8k/4d5lYxacKi7iljPgMIGjBOuCFvqhlVfweMndRvAJj2vjKWKd
ioVVs3ae6a0t78P8BqAgunTmMg+3esJQzIDqczdyx1hLRdovfYnVGkSZbBILwuUp
BC4YetEwTTuErKGaUAYVMp3Qj655ul0EcLl10E8RvUrtdiTibIkFQF6u+JvotbDO
rTl6OpnxxB/Jf9IdoXEiHEcHu6Rcxbb8/Lme9lefhmsmxeB34mXUrWTznvjnJvUN
L+NLzNh2a3QO7AGJ1RgEux+1JNl2IG0SM7Ntv8ZgPUfMgIxJDS+6IfaKZenreSLd
HEznPiuuSGigvOuLG1F4Uad6JMUKLmGri69u9+4LNSGtHLv7p8h6RYQSC0f3JzqZ
dDLfJ0FNjFGjnOeqj8SwQU3Zv5r7rBx9LPcJ9v7QPY7Gt/jcuZzxSw3d500Hh7j5
VPnp2wySnNXxFeqI3KUslpnYWCeKY7jq7gJgv5zX3V9n5WaIC2i6qOFhFW7cFhYJ
ogWeaQrgWvgWhIq2AOGJFJq8ev78Qg/aXlXT2DhgPMUJxv9FtgSAN7zV804wCOhY
vLqVCLrqpN+xdUQjgy5gVGBtkHRtW9p9IhILWtu5WS3fASLU4PeizoTjXadweoHc
KeTuiDwJoQCY1MaHwOSZRRHVh7FcGvcvSFmIL7QtOtInF3sZ6sxixmJWX7SxXYj3
60WqEXppckkyO19HqEeS04PKjBNQ3uczCRUKjTrPBE2pjuOpDMl9XcKXRFaOoo0I
PZ6fHHN+R3v8OXOnuakBY3fCRKh/tGLuhJNC3kvrCRRzm652oi4o9auIZeuw3LsG
gvr1ip9qq7ecJ8H+eH0KsSabqeMsg+x9tv5yyUehJAiKdp1mXvg7dG0yX3N9/VMh
KfzWLPKpApPeLkGhd4JJ0ao6QXfsooH0r//3N/5P1kxwocDVVHrPMladc8F+x4ce
ocKA6CXg2HKqZ5uaX+QmfNEN7NC7xWsv37KTzJSgwGkVygEkLGoJz7zRjgmSN+A2
5dMy0yLJuiDHvG8zANgOMeIAlhtF67sVzNue59JqsESXk7TR7neGHXHbWKJ3fG3+
uR+y/BJ+Eev0VMggooYtP1cpOxPvUP8Pb+FJheCA62reA4nSD0rPsJZTrMQ5+UYu
F6nBI4V+noUQZA2MwvcfYUp3UmRF3xj8hXCrDaMNbzMS9xw56H1JhP9er+1f2/Ch
Ogbkz9q+KSi5YJyBWQ+hHX3bD5pX2rl9nzvUtQ5jiWzdfk6XJChJyjgGXhepQJEB
4XuboAcq32LQF4Q3VJqGDGkS4Adzh0lTiIPG2ynpM3/fSWGbPCU+PXJuoKjvD+GQ
ZJP3GVc9zvJMJshzzXWGOHu2keKIiPVwzZXc6PZBxGZXID+7PyZuniK/E4OHpfhn
PFtv36pJz6c/ntcHDBPT+vCSNmixOYSOApUKR3KDmkbQAeWtd6kpEcD9rrgKueq2
PTLr5rbH67tH5a1rvbVe1xRrCef139x8eUb8UCafhoiTRyZiGzh9gyNyduKyn3nN
QEhhLQ6Tj+heiY2qP+Fb/vtiQVugyolMIFMA7SSNjusmWETleC7B0Qo2bmzW1f9G
tojYK/bKj/33vY+NEkGLMMCDxYS1Tq0M2zgxMqQPSeyEwWy3Wvn9g/Axhp/M27OV
DMjMa/Jnk6liOeM6wfe8stKG+2CNQoDgihZuCJiqCxrqh6UP/xWWZdCbm9I47EU8
4Qex+OeUN9D5gSBQzm+Sg9Njd4Q06B+3EZlqQ9XRqEUi0EtzHi9BDD9NSUDkJh01
6bpxFUYkp7x8OiDUzRjIhsAFGO6LK0rpzXiRv2mqsvVJ2/fPNJiqhGpoIFEV6xg4
tJ595MUp7vfnVnL8ZXCg5+TnbSU4k5DCJZg0R9l/b4310Kqu+uDvtc31eV+DfKUy
T1ZfomjHrRSVRbdtVV/pWM2BVNHCfOUmFG21Sh9rSUdoeyHD5s+GlOYyVmpyS7e5
RCTzPLdICQIfiSC7kqHf8tlA6x4CbQiBHJ3/e/uIVoChMJmqrWbRbzk0SpUg9P61
Ga1mVdutn0oZhKwpOoZYxif82+qms9iuFWtS4i54E5I1qc3MfpI2YRzobTNlH5av
dp72FaDADjODYB0Rvpxo7jU20MmJwGEpfnMpMSmwXLR9d3KRQ9AGHNelYmBNiIUB
ndgJQot6dzHlhsXteLMm0cg85HWtrsa/NNUZeL4g369IDThKO1/IDfA5+zwBTBNq
6mmJ869/2nbsrnhEZZ4s+//6FQ3SQP0f/eev8Dz2r+TrmzJhdp2QmvT1u5fnLs5i
F+pfMYjhn9mUVMZ4qitIHHIhq0YALQlkyi2bdnF63Yu43VszOD57rTfnrVEu2LkW
JU9m4K/+ew6fwAixpxShz6+1lHmUR7GO1imgeNzQbtI1Ar8AmFMLD3YJGbfVwUk9
qSPShwuOxCLNL9NvrR69qyZAFUkXAnEzY9307hNjnbJpQn74KSDbpo6GTkSKEXok
w7JWkZE1EZAMF5LhcWsVz5acB9pW68Z7Bi5jS0mOTGgn4KHQamAldZx61AtOf6qW
Zfxoj3TfExPn6GbKT4KgHf7H+/VV9tGSralQWSSYmUjsexCjOBkZEq0Fhn1VttiY
N3Yw3qQeC96vuZ8o0M2wsskES+KhjXxrv9TlcAoBEo2K5C2PEfAgwIeC/Fia+XtM
k77G7S16Aiz9yIt/3ab4ZAtDrnwah4NKgB+KKyYdiWt5a0nEJbgsl5cplnGYAo1V
B/52FgWn5MKSeVSjwZtrbOJClApirywvxNautIFjPlmReX9fhFEg4I1PJtWiBYWO
NvVPlEZdPCJBjlEqJmzYNMgliVFs2A9rVIwxLMfQkkV8qLzdGnwzeA2ssjfTdkYb
UHrLaoARjKyLvvvqguJAwNHpPirltevHn6f7VaiRT8qhjJ/uhu5bn4uTJ3d4e36U
Eg67nqvdMt/z3xHcce+Jukd2nVPVce+ICQTSUgWmqRXRlmS7ytn0ZdTnuOXxTE6d
NIJzQZjMfoaNHMIumRDzdtKAe7prDDobnxArzriZ35pDXlITBH9dibps7yYhFc01
UwEl9gPL8fB+iOuad1RvFCG15ZAQcCM3Lx9wY4pIe8R3aZOzHqAEu7y6tmX450Zz
WiEdKV/P+NRcqSEVrNagYfvlfsrOKSC+ghNSM7Nf59K/2ZU8xo1NpsQN8Hy0vh21
iiig4JUoqXm1liZnXXT/EQZa1JKLpyQmeiBVuv+RcY8iZ7CZDSpDxnSkuYbdn8M1
LvrtD6QZq2TYepEC+yBcYIaWJUlNXEckB1fUlkobP6OEmdykHcDgroncYOtgecKb
esYxwrJV2WhqpXywXo8ELuMWSE9C60t1Pd5kFh7wZF9NEuYHnkG0e1b0M+b2hsvW
AVkQqrkQWT4JbyBR2hQEApAaAIyvIC4mgy0bKzbLKnyR0MyMWSDguTurZEz4fahc
4xopC1dVIZ4P172P04blWmZuhAxmTynZlHDoIcw6Qw43zocjYAMY1w3/qdRr3wsi
K3szfVAkVvUx9mHOHUrVe8MAp7A9g9dG6ALeDJoj+6XmG6OiqhmOrmXw9vF1aQVV
iFo8pX4qyprLkG8Ud/u9/BTOoJTEPunWj/EnrrbPSPDjPNBILAXJMqSrREgIMXwE
mcuNimM+1HmB91Y2+x3T+yTcGYOFYDjz/l8nVpc30f7GpzVTfy+Nhn4KevANn0Ve
fRECLip88c3p3nkXRmSGfxViE2in7KVc4eiXYf4sP8xtXfrceh0/tp+3jRkNd8t7
arYNwdQR0wn+LcxxUdVScgseyycQuSbPr7o5r9Z6dltIVXR7WvBKSCimv5Nb6jb8
qFNuMPBl39zABQ9pxNXyDTflOSGLo12rmOkaL7ZsowcqLTBxei4tVYC26xfEtEJN
B2iX0hI9VDnnCrHHrtcPCiJXn0g+A01mDgASy2JH1BlUmLpJ/tnYp5ibo/flzhTS
6k25QYo6gTkfhRVt65jKX9JRxLaACdcTXfj7lkNIRj7NdbMALmE6DwmpqgtWvZ+o
Zr3eV/TMAB9sncwHASkLkZaDntzVJR3wsuOEwK0atnSccwiQjdtlV52fhR2gnuxv
GcafQAYY3zKg5CLOeUQyhdP6zISNFUX36peb3N9GlxvwI+6OFCx/4ct1PmM0DJtq
wDScsx0z032cC8dwnIkYl4CBCU5LmdtX0EizoNRIZkBaxqMCZ0QvXMIGi/hu6wyT
7NOo2QTtKmduY6T0dexw8RNxI6G9tlfqNtv7gLmTdMj5DhpB5TOH8S+puXKcJ0ww
VbStCinoA3dakMz8Y5UN+JNrBuj3gBhp3kNnx3tToe8G3Te16aYotIvCN+35sp5R
yK1H0f8Ce4fqDh6/h4Faz+5w2W0m0fMmVSnt8pXdzRLwcl0tJLemcZtXMCN01rZg
WrcLKSoLka1n4dNMthQYJaL4SrBdx1AZVWpipsPeKL9Tw40kxQ73R7fTfpx6pgQR
f/p9NWorohF0HFVkCWIIw+/oaFqAxTe3OUZJ645ufQz0yShqzVfnc0US24BafFQr
3llx+v0dEI9sPx8/gUEFmBYl4fVEiXstuElRqiQ50N75hmBmcEaxg4W91ATpj1KG
Qf0ROk+15FK1McN6DSvowGFtlYhJwRDvzWl14LuhzMxRBf5oWpCbajWw7l7nyarn
ex1bHTua+ebDFBD4Baoun8RDBDTf84FJ2M5W9PzdjG6gKn2FNazWTGzo1PhkQQb5
4vvP3eJvrUMTSNyPjjsJqgb1qMnFFZtwVbla0WGvirq0JRUMWkz1UFiunzYCBETD
efqirU9suQH9YvCnUx8WFaiOpEfjXRKjDuN3Cx/25xNyjpf+g5/OJXMNjQkhKvar
Ze8iZuYWGMNcWW96ZA2fOpz4T6X7O1Msgjwe0qV2J0LwmHQXXOVpawW0E/oICQXX
e5xaeqYdT+ujzgx5O0CPT2K3E3JVdGHuVDfRSeDqDqCbqTMdd6eVN3v2j13n1GKj
diGvShCV7Cuf5aCnryCThI9UUIFCbYBndwKiLPtVBEyIKS0bKvej7J4WA01/eG2k
BvRFJgAzkvw52TGgGJgbr6jkluDgg04cFdUcyygistir3PhxN78d4fRGzYpaxlGL
F+uJtGlLYAucYfxJlkagnsoWZz90u/4+BXxy/6aGrKSXcEoYHDincy1sVNKOB9gT
jnNThCbitTsj+L3Rr2k6E8ONCHrjP+YCcVTguBdZkRnnd6NHDMB1SHeg6Ui79MxS
6ehjcU0zIPjG8kyV2OG/uAsvZQu6GXwwUv/8h743AvceBd6Tn8hYDcqhi0qAAr9w
vFWLW+8cEbFVF3+LqyPUIxGuSavTl84sFfXk6boFdc0H3VL6+0C4fV3dYG+HeNdR
wyCuKoadtOV3weJTo//7I5CsMlbLVzJ9ceI5KJYHW+m/jsV7WV8bHuctlC5UTzyI
7BJG0skI+14eFBiy9PB0xPSeozjZbBAm7WdGhetpEv9IVqGZOW//0Z9EQD9ksSp9
1YWY54IbNOEW4jyjtFQDGEQizXWJv92/pYJOMVXIHleEQvZA8A2sI5ODBN+lH8im
njE1GGBvKTr3tuBfa1gKCUW2NTKWVICQzEHu0p+2MbRG0ZyBXG6Lp7OJz9Q8EBjn
GDaW4qjRpchrv43tQPf8pkmdAu8EWepIppdllLGbtYBexbmnv0K4eRe5+CgRY5vo
O8UeKk539VZhLYz5ElHbNTjT9f8soRWBBKX+B5CIFQeQKmW1LjkgXmJ2YrO356kF
l829uG5f8LmE67DMMkb0m1TNPnQDq6M2envL9AyK36UkcrD/Vai1kvIaNZPxxW0T
mHtAeZM4WbkbvAgI6RDhnDxytThZJURB4wEESFb3yQFjreYOkNEzYhebhQ28ytd3
LjdCy09SKwUbSoI0KVSExWpbVUkQSTiFTFIdK1vr4DMTrkWRe2tnVgj0G0b0nfMs
n2B3ZNOAVPyA+7D0b6eMkcXkX+vksZK0KAx1z8XYEfKQ6t0bEfajZSsiS9mU9Mrk
DzZMqXjgK+D/eum+xqsx9IwA73szLDKywRGzSyNW9aeKh5lkF9Z+3nIG4hRRIZgk
HQgjgOxEIjUgleSI/YnVPQw7+scDfPUGxpjt622VW7dLg9M8pYTdhySdPFVYiJpM
JMcA9atDw6WXjb3C/IX98jtHceBZHD3XHaUe3yqF7xqy8dAYaHwS/QZaZJy6wbr5
m28S7XeS+83VtVmlXeF7OxgwV/4CFuHG/+2KhRJaIug1Hc3Ud30dSqh/zpxFmT4X
LEUNKmd361l2fLH7LckXfNBCmDbCR4W1yu6z2v4Ao0jm/X6VpZzc7bnJ7anVHHL2
0KDCYCnRqD0G5LKYABToPKLssMQGbU+efDwo95xutWNStIwE2xKRT1mx6rEvpECe
u2PRKqc0DNerOOz/V2JLqAVMHbW4N6EOtgEExs+l7qe7wck9VpPMhos4/XvV9Vri
caA3NLdW8eQ03gqbUhCoNDlFNUGipUMEys94qrSwCErpuoCacj976eEj09iCSOTk
2Od1p8GodpiyRmFjK8PhodCGx4a6tZ6brOfgvZqzQLZhxYXxxluCEH7WncdKv3Bb
BVNVdlttW5IpdDlBPVCwd80yqTy440tKNAKDGSWxcjlKRZSOnWE5KpgPKgO5Qw+k
OnN8XEZ5l4JMmW+8dZcQpDKrKBzs2kY029szo/RhmzpHnXgAVaJsYURO/47R1WUW
hsF5C6r96+iraa+n2FvBA7CWwezWXLbBlPJ1AMmMYhpUvr99cUVL6JdqeBp0rccU
f8YaV/kV6s2I0wxm7/iPf4NTh2X3+sll6lgmyDQPBhk7dPB541GD0SxRQvlJPZy4
2VS3Ai9e4bSX7Ck2q+531QZP1oilC5DDYDX3tDi4j42uoEDztg8+JJhdHWlzJ/pK
4E+M37vofvVNmQEq44Q+/Q3lqjsC+mLzVhDf2j8GvpsefYmeewObEOGZrXHJaJuJ
u0WTCSRNs5+UxRFD3bV9Ee5m50TA9LQfk+NVOhVbWVMU86K+3xd7uHZP38qsMdSa
Mbt/BybD+x+50NxdAle3Ixe5+0x/0PG9KN3FfVjJm8ibqZZ7dkLDt7sWsdbzZ8OG
zQ7SFf0uAShrwLmv3QNN6SJ+6xoarCmEwiRhCdOWlCmgqjbyblwAPDKsZLUH9FNP
IGozkd8CxkGLqxgF5IQeYCQRDCMVyWdCOoQ6lAmhGhBo0QNOS9U7ksQ0hORxiFHZ
hqsD1TMvSa8kdeUjFmUAuGscucljkz+9Z/AwkpQ6OKYHn0FaPBNfF3Th4ICweP6n
uotjlEMIQnFyD/7I7thOTcFg8JpG09TAeBO3qQrgaptmfyz+beSvcPFSARGrAlJ7
GemRamLSNQcRRUWk2CaoB6wvxcc6SSTSs1FPy1s0YPtp2XizlAyq9wHsvO8rEIGa
d4Srrf0PSj908ouTjNj2paeZAdktzDfzpEcgCyZ4V3X4oudoniyO7HIM8Ac4cuZs
2DHjgoAyHJ+88zmf1bdZ3fxzksqK5ADvJGUXH5kIwXYyJPsf90M88lubM19p4WTb
PyQxwEX1ZuBUiKBre26MC7N1+CtXyD41NG/Atk09I49nI0B7pJgeqpsgZPCsYfDu
Q7TJTz2omGrBX56xvYZiqXees/XLBMNnUyY4YsYDhjcaOMSqkpLVcBKMB21z0mQy
j/h8FiH08vKPIhNAOSdyGVGTvwF5oIYm2pxQDOJFoaJ0hGQHDaWnaccB3/AC6Fk3
BtakxBVI5FgxuHYDMtl9hRgw5nxB9sdhgqTTZifmMaV9SYI2oYT7WX31xh7Jxj6r
UukNtrIb5mbJPnp1gXKkYnBk1IrKmZT8J/w+VqjIXD2al+mJhhEutXmWO9G7CNx2
3U4YTuBXVw33iMeWjTTH/ZbNVJ+UP5Rqr3xsmkUDb1oENrHiRewBYviLpSSI6nZa
jOCXYWaon56KSVHHul+x19e4840qepqLv1FvnugsE56xc/VHl0ufwVFqhwltVnhK
3miwGi29NBxGlDPIqUm0KgI7RZn+fZuAkO91k84+nM//CGqGg+ooAR4FyeJt3pLC
rj5AeFOwtRrj2QgnXL9gN5dMum1v05lwedc7drSoMf5D2gZJbTV7c7jOcgKBwOGd
19yfQViDuFyIGTyJr8kQ7Y7hgYLiIouj+ZuC0fwmtZ9o3CuusjAwp42Xd2LbkSte
tHL1HFXqPVGo3g58VY/WIk3za1kUAUTzKeHe+TAt/B4E0JWmFzbvzymIRW9zEGK3
DuZlRIk55mDMzA1skdBst2QUpq4LMMB+y9XRnRwKdd86Q9kUmTAaKk/LO04qmeUG
IPjvTMZ9HRqlg9KwGbd7tmXN0sidnXvlaGye+KGpByz8g32zZkas4/9Q4DvvvCym
XI80iQawbEONWpzq0Hfbyb93uFzvm704+Da792NSYeMpxwDHyOkF+je+ELAJcB4t
cR2HZNX15178Ae3phBAI93GF+GdMKy3m84U4qSIi695kCbsfROgPrb7hnBSrQ811
YdABtSRlWM2IGou2z2K1FPaiZmST0+CwKJuK2oH5cqSK2jPepr3Oj0jwt4GpfoGy
YmPErXoce7j184YBavLcqM80A6GQ7el/yKbPwl7vuTpD9PQt+CgQb5I+3WU6qCg2
X8dJd8XbLu+QqLYihQ3ud8rg3RqCQvkE11G72Z2ffnzUjMhOB9TQYvOZeQ30MH59
g6tD7MG7/a90k+5cgDqhwmyLmyKE2T7uSRJ6l4f4J/5LM/jrHodwuIztfLmbuV19
qnavahDyHlen7i9jHC9XF6VJRXZ0m2ZVbu9CMR6Qwq3P41THIpLvQt4AIV8W2nwb
+IfhIJX6rJQbCh2mvvj/llLgxIRW3LuItLRh5MTjgYcWLwo7crLgwZC9NTOtsgpz
1dDbxOCgzKXUR1iwky8k5gJ0RQ2D8VPvGSLST/ijNe3mNVAdSobQ5DaQ7dOvpRpj
7VZ55TtutfUylNArYRDtde2itT+OVd2JMJItv0DHkaeaRYqepEQec+eSPxlCNudX
R2Iu/6muJGCPPGpd+BmsQLR3+1r+tQD9MINm2fNqURD1Kxq3GEfkKcEpr9luiKRQ
qWCBTC4Dr9rjPhkvJBjkPwGPPmPPYAEySsc3zUNwFr+PGbMSuCXobecAL79X7xY8
YGblDz9KuJks4M9VQCHUDTt3bPVnKSatcL364ykTYeFQpb7e8YvewMHwS6FIV6er
dMDMQf1FGz68SEvAOK3q09XrMg8LmbUwNlv019RQ2jG3RRWj7tbxrh7QJ4zmB/00
uTv12R24EYuNkuggER98tgSDKCXD/s9Bq5AF5KiLrk79wnBH6duQE/WgeoX0PDO0
wig5k3ZUkWHaKezhjKl0trKbf1xgdwqVm7MqcPHaz5iMqeYl2qhWlcxXve0VxDSt
hbSWE2Xp602y2TkV87UXeJ5iSldJIKz47Pf1jqXezcDIfNJ5h+uxYD8lGkykN7WT
edM8CqDOe0wRU9yIV3qnwP85NxRFYtQE/15YKr3AYWQ7GbJr/fSpljJHFcJujz0m
LnAbs9tRIao/aXntWIohZPFs7SErffOUO83ZN6kPQ/DNOfbGJA7cyBDbIFlOg0PR
sClUxdJlOnL4YQsGB5J+j8DcVQ3zG+k726bUp2el4GZvtEEeND/nEwv+X60qmz+8
mM6ujrNteeUR6mSWbLPjBI74jnI2w0Flp5a03id4Tm4cHYEV9p4OwlG58O+NyZep
eSwbcL2586JCGt2wHHFIDvItcFuW48Tf0++k7Cdd8uyUFK2+SLNNVH3tlJE2nHOo
o0gtCth95NhkSs6hn83o+TQxldxswr6qHUAuDg5pJUP3CiO/F0RtpkP7NCdNTNHV
ahgpj7L4km/aYKRAavtX+D7xbcKWI5EQvg1ynCUD9m30fmtKwzcPnW0gp62gzgWi
wJS3zFmfHoFLrnH8Pk3TTvdWd7OWfnpk/OYOmAdpSAJfcd01HOw8vmLgs0R8qynh
0nJQnD+Su3WJOQAK/j1LJzNYNA6G45VFZdFvg+5hyCYOqjk/2FFursGJy1AC6WhL
9a3BLAuGlHLYrDiQL9dGRohWvBdavRMdwP9USpMdt3AB4NQo0aGo4dzgF19zCoBH
F5t/VqBxAwAAOH9Jj7FHjkHpKCrBp+uqcxWeJqbb1TmMq6vVwzbc8P62lS5EW2nZ
S4YlB6U1JBEheeiJs3VlmOcXOjBdiB6Oyh/FB972HXXFfImxEiJ3f4+Fla66YYLw
hoSw06O7pfiJYr4ZQlyPV8yAUghwzzeq+tAGsB8Ki8rIbcWF29leZkf8f1Fbem9j
jU55eMRK2rV7amUYc1ndEbLRayNdDZmzXSrOKiNYhsz2MT9n6BKB7Eh+21zYrgXe
EyybP2mpGPTi6zEbhTDrs1EDHVyjyUUSrZAk299XXt/2S/da1pgM7aPbopvhsh7m
qx4Gpr8BujktqVStIdtLa2xLWO9WuAPP25CG5m8EWnq1rMzQ+mTnygpH+8POUuIu
ODFlugDG54mqnDvYEwsjEumV6AFiYklPAtwVjMJs6LMxab7hzOMtU8x5563cNFQj
pUx5CYgS/HmZIbNvLx7tbz+D7StgUvGqbxi7VgkT3lt+UhonGbcIqqWd2+tOzxk6
r1WjjKO5pONtlHYeXZQs8G3L5qEDstAcpdAdjonV+R8zjOx9EtqWec0CjGAxPra+
N6o+YguqbySFZZQNvdiV9cbAKOY1OIDFL9tK5MroJQ75E+Vb3IlH2HCbhq43DPjw
UqcmnH5QKJKndttg8JrNKQMXImbFkPjYG79S6FqX1m0IqKAPAueKRvoGzWZoJI8z
qufK3/9iRVxBe4Hm5mDHAQjX+4FkXKY4myZ+StFRmBeLSXZAmOi4jMAjpPsZUEsa
G9wBkFFlsrikwAERvIduCMXSpWLUXezC/yT/5mpT066LlRWbf5Bgbt+Un321P7WJ
7wZ3RTAfyFs7+E+Sz/heX2KFMEPC7Ex/krCN5akLN3lgOhMJYbk4WtWi9D6cPQre
Q2gqm2ekvm7862bOrT7Hruw8TuyepBzvdBBZApWHOqOY5Md/dmOqa+VDqkUtdZZ/
TFJcs61SqhfhrcPPt7Z9CgcHSzkPj6kK9L5IlOkLR/EGpEp0jYqRLm2PhIrLC6Fh
XNgwsU1SUgCR+3AVObhmNzF0U/B1o8d/Q5W9xIERNaquhWh/R5mPrB/53Ah0B7ol
9m5cocuX1sgKP8EdxlJmEfp8MksEWVqwfO8I4FQPLxezCwOy3Wxz5rRmpG9Wyfd1
r9kmjLHSTaKPUzX+UdoNOScK6ni95X6lN8sjfLCKbhwjoUot0izjJ3V+1vM+iik8
/mLW973D41LUYsBB5Fq7mr4soOiV5DkXkbMIIH3V37+5dya1O/cFEp0OHYzW+6Bw
/+CKC9YickU/HEHgDwKFie5bTCVjZfkgougoyPkagg58Zvng0OrgFPblNLELMbNM
J03jtEeJA2rU4X/SLoVTui4McGe1ZkQp89gat9O//Wrzy4FjnIiDl+ToYFu1m95N
5wJxjvG/+H7wJVDPU1H21poWtJN/E+moIjexpRaozY9kK10Mx33/2TjmipG8IT6q
QJ5yQ1yX/ZWOWUO4L4YRbAUk0LRQchduxOxEIeRbhcKBaeJTkqR4wBHu0IZuaRhG
uRk7WbECIj1fxGbiAfNbmB0ymWVzkoPFanHM+f5RBlpGAoq6C4LAWyL5eyApczgq
VJbWm7j7jMZecqLGRViaz07WY/rKrrDc8nR0AqeFrV8KK4oitoM2R0E2CG5yNtnn
5/UBdna7UgNLqTZMr+/uWhlvnR+6/fCcD1JtsQNbly+gpEdJSNzb88Q60J+foBGC
g2gXPpW7Q4wVe2lN5Kb3xX0R/QHPV2B6wxHfXd781mBTC+Nk3FSPA1tVnse7n+Pm
fpZTGK7JDvYqXzJSdKvqmfNMaKXUJUknruHW1zqgFv44pjH0P+itDzDEw9tjMpXX
rtift5lBEILHNPYKkar40yGIv8AGyoIAbBqzR5502cpL3LKgihyhAiN5vXj/whZz
aIoAyzzWXwe9i9SWMi3jHY9FruBhyedkanT3VQaUzMB8FVLFvRNxqa80ZmgK+QV5
E7Ummc4pMjX998PV5Lu2+T2ZUniJJ/G9TdnZm37lwwaP8ZjCB73hfV+0OXFdaIaV
QhlgXvVlvoBPfOBVyrTV3rozP4HDKD7q0yIg+swLEvMtgYU6hX3AAlJh2ceYDvqh
XhpkjU1J5ZG7+UG+xCuzWVA/EW4xoEOEihjSPlZxl/jSASvy6LuE74/r/iHQhbqt
SX0rhFvi+nCdYUh5OWmGg4gyeFVaqy5O1bxaq0pZssuU2pNcMbds1cJWsIcv6OhL
RBn12Jbf9Zk8Do9e+ymC/U60yvztH/hPae6dlbIMJEKszkTTuE7VmAUxsE/y0/Rn
rO1YSXCg4jT/YKI0irJUjfAQl0HR+LgZJwseyvTgBn7h0XTspO5+g/Fs7PxKnRQV
UiqTG1XR8c1JmxPlndz+ht1/nBX+tlotJ8WyS98U7z299puxBPSupXvhMN+kC2bW
cV8499VJEoZPJnvSOFgxczhepZstHkkntz0S2lxOIwNehn+/B4A4N12BMSJeWdpi
5WLWBncALIKbcQaHydJMTe4AdXGQSn4yQQFJYrnVeFHNy4vgpgqynVQb4SEAoOOo
PxiqLXD82GB1eMDd97lzLwU27P+W29TY6CvRZTy1IhsQnjLfoujkMa9UdI04qhhA
0AnFI1+3kKlM92NHvtZjhaIKH9YFXMFWPyvpkTJ1gh41wgnYip6VZq9CMkhZJ14L
2x4ihtBjj+Zk5vwso7+Mu7ICP0AqNeTjPlkOOQe3W8st2ItP5VoZEy0ahpOAxZyL
puHBZuGQ05TrbZcbTkE2ny5TDwZ/NyoQkOVRI9VVk7wX6TkhDdI5U15IJcQhXcQ9
wyL1maMJ/gnaFXkcqXuf+L70cA5L5Ftvnjdv34ecB2+SiJSYgh7B0wFP4lfdXK8i
0a2VBluezHznvPOm7c+qAtoLInL2bmUd78e33KwydpDc7WrSU7JUl1/srIpzNEeK
l29ypkTVpx3Tcz+BBCJJcXkGATp+7VLzLb+h5C8HHx7YvU/fkCXFKozszl87IwXe
d3wi7RpaSIeLk0YGHdvhcTri3kY4t+VXliR/ZDJ0kbd+vychAEabeAz5S0iZewxX
VK9pFdHTGN3HI4D1zmku4o8stei2ZqMcykCYb5h3o25zgZrnIvQ9f7uaaQ7UE6uX
VU35dyqkjmL/9XQ4VodKVwhwMaCdz+8em9ch1eITrYxpPP5flYdS0ZigGZLRU2iO
wRzzbOgF8+4q1IiBg3paezHBnekU42q5KnZ6qKNUamA5YQRjE4KWDSeUDs7vE7gJ
8majeGZxjBK0oxDmLLCTrqM4iXib6AtHDpdC+wIyw9cqC/0VLKMr2tlVr3KFnOxI
blGsPeF9Ij/i/G72/2ob30abMfQdVc/Feo2LKxhmt2dZBmADCtsnxk1Tr/dl1z+5
1iFuY4Tnsite/Dy5JbDcIZT4R1raF1YZJEovz4oPwlh3oxPXk+qkW1nx+hqEnpf6
m0p9KmW2qXNohTrT/wea2/ZlXfZSL32GeXWTTSyglCDWioEy7fVCDosY9P7ztQb/
PaBBy50GglsbEPLlwn3RPEFT25Omfn1Fv8C8FSo0O6DK4x35PQWpzKMWvlx+Qg6c
Zj6SQOYG8oV4qAHHV5eTmPKhk2a3esDaiPsS8eZ8oGPW42D+xL0r09Frg9hNKmzB
UBqYhIiDM7Ic0qfbc7LElL8t4LaiRLyQTnNFL5JVTNpSRFPXHpgcMlivopAOTMB1
1C/fdrCu7NAU95L8J6NFUlNaZo4Izu3bYSwXZhyFTrqArSs1dfgOZ+sq+LDB9PuX
DEJ8tj5h4lFNorT/a0/U7XIFISEFpoiHh8a+Ej4ZnA/2gLI5dfkr4FA4/DoDFcSc
gL+jxPJxm7Jr9/0FdEdjFOFMTDxpZTbQ8ztI/E4PgL5LkiL263yxeCQqi8Dn6Jgy
6Ymwuee9AsQaT0SjjfBar0BzuzyH8mtN2qRd9DpkGW6zUGyRkOAGbMNYvlUV5MAG
DW6Y2H8xAQB6X3jnUEzkXf/QpHthSDUmi3CKNb5/kH9ekIUshnUyd42g2DCgaRVh
+EwwOskBrGzqDkN3Uz+SRSyH4jdM8l9pWLFVcKxl0pIO66a7tl3MI0mArMDm66wX
hqhwoerwa42STVOfLQW0N1k7SiAJP6fBMkkN4rqR9N+K/EymkHTIeIL/pZFfpNJQ
nbcSyUp+Kve5bbxMR0xaKUbCfyOPbwKmEX90roMbwl46ny3lAA/wst3wAQCZhJa7
MMNdh4hfzEZ7k8CodO0oo9tECQ8WO4DGBaeB9hYjzHRVLvvYoqdTyIXApZ9f3l9h
SXsl7FaYa2OBtFal6iFdWXXigx1p27Ba96kRbe59GupoQ3hl14UhtB1iDkeGvIAb
hTMZsfkKXfmidZhNlhf915ot6Qni9uvx0mZFWSLx0Pw+OReGpmn8Usx6C0Dj9P+T
bWDL6+2bdQcfCnsGiEFuGbmwMtoercXWvVPkpgCJaL9iZm/FyLePzFlBNgxbB4/f
IcivYugBY70MXyUVpziQ01Se7B2dev9Gd9ZxMakiQIayO8Sh/5kgeQdqBcUqDjc3
BJ/ovbPljwsVT+jyFYdJV1XRm854PkrouDDaKGafVEHx9i9mvtthijtishUVY4hk
dM2KbJ5gYchV/on6J7IqqsbPllRsf5sVN3zdLtetlVJS583NBVi/gTOxAw8YM4ZR
d3n7N6IHc4F/oIPiocbSqIf6Pu6c1qNcm1/cKOvft4wJeCeCYAop93Vh+bbiJBwo
YlwGJvkINmXdUNg8RwDr9NqRhdxY+Ah8T9/2h85zTL3/dK7gbKCK9SABMs6kUSqU
/9g1eJWMYIYDOTIAoLCuDLpG7Kn9cK7U7jY9KrIsuJXeDli/XZIWDiLwEJIfIkit
pVv2IL3osjqLKeB3LEI3El/OVdZGp5KvJezQmpaGCZ6URHdEuqafD8AF/WCbRStO
A4kC9izuuHRkgMqARAZ/90C2qSYzrRS6w7MoakvcAwIejVlV1HKxzkKGt/yQ/eod
ivWWqfw0DKrjQlO6CjWtl/0KCkHYLi33zrnVARC0kn6HQgbwSPJmn73aSfVYT3ez
lbxLDJosyV0eRchT11HyLQHsSXL05XFB2OXOlX0tFWljD533ClyFOzJ5mLG0LpAp
XpdG5Ar+2xdx+b9dVEwDK1xlRrsQybyxd2hIY+v8NwTOl5hZzH4f/O2m6XYFK/o+
jVpvBgXMXEwgCFKQdtB8/1L8UEynZYRtknniEI8zRupNWSP8KV4ca7uyPuRsQFOn
d2XB5EUUee7r9KKR6bd6Gymj4whOS12YcNj+5bVzqXJi+zwTI80kD0NIG4pFwg2a
O6STn9d57JGIol9yKKHEXEMg2jYiHLLYbzmG+K34qrfYcQX+2y0osaIlc5FjYsdj
ror7lzEIhfzLNfVmPKbisqhiK7fet+ccv3w5EG/4h9UIx7sTPb5v6psBTwDkzlpJ
cnqWZx9XhCcsta0ltoXtd6cZzciWRWmzn45vbSPeu0xAdvZztQ3HlS4boy4IByv1
7rr0H1Qo8M3ds35uPz3h63G9wCxWitwXILhW99aumNPO8uQaUIRohk6S3EfBBQfL
Bt/pPyKFJ5KhMUKyzEqajw/wBQm8YDQOErLn1NWzAvgiRTMIPT9nHjLRJ7Qf+vsf
z1fVHGvhp7KHGZKQ4LwMT9imHKLnD7QZzwuPoHd5YQwf7dw9N7z7IC5yPP79okaa
hCXuiuFCGYbfbdNBZi8mEcJWGIRsmd7v3tKIcLat1Tle3OUpL3U9ClB7XDUM3vfi
UQkh/470CusXbILPA7HKqNWdh643jRSuj14fbhlzGiEqS5ffOksGhRgDKZZqW/MM
WeUuA3XPGh1mucLPJQiRQcRUfGFRJgpZR6MNfgZe3mP7ANPv9O1bMmrcDJ+aDN9L
irO4dv8ZYsQ2qmTQxpGzoo+/N0tBXqOnyuEasm/8U0gaORqfj2Mds85artox+cWj
o0KJuLiJDBz7E7Ma6taPW13zXbitMu4rCSHQsAqfF/VpOPPNA9U+mrwEFaNYQoXx
6yzmFjoUWmfAkxzdGHbuJ7R5qb+Ny5LkgYCx3sTGc+Qrmcoe79geE2HKE0+RErkT
o6agAa7st+ksxOvYpoVuRR2QX9BQX+l+6gqXdDnaGBDZ2URRONY1NKpi2JtorcNY
5Hnd97e+0k0kOo4EfwVyDciz7eWBBx095oQcio32X70J1pyqJIQ8je1gf/Fmn1x9
OjTqjxD3WoYJOBedn6ck1ZQhczy0UgWPm1oRg9uHrpHzfodnG6bj6uLmdO8Um/WM
qVl5yQptiwbWGhG10A4pxeLo1HhLOzK4/8Gwpn952ZgrOdXwYLyGSrOGyTIjrOYr
72egVIgmhcoZiZtEEqwrGIK+dcwLbLWDKk1Cm56gn+D3125OF1ExpezMi6NyOReo
vIWezc3nPeu7+Z8gVbGRrRPf95J93ov3ZZMvXUV4Rqkv+0HeARrqoVPTMC/2ZlV0
Ud9kozs0RvLJVbEhDmmqGqwLFrj0VLOdx36WZU1n+NwX1TVp7J45Vjzv3Q0XgwWt
Kc7xzN1wr06NhtftIaLl1OCIY1uRtd/i4nRiV4+bxweTOH4GEETrpcbozjtxSWfd
jC0uG45Tv3uRBoGL5qc6/wHIjJQLUQYamLWw+LX2G9lAGvX2lmIPIpa67wcYapcg
2nwRrqMgI8s91sorNoPQhEPaZzCVrjGSKTmgBJoTGZBsZzPV0QCcLvcrSVNRP6Jw
HqlgCkY8gMmImF4rSblPHKmgcgQxNzeGbvpeVmemyiEgyGOOhfsuvIOJig54yKQA
d52ch+OcngGQGwqwJtTIgc4eP7gVuoYld7jIGfHHqJTlNvhhy+7umoX1zqM7XvAY
G6y9y5crLmqF2XGq8nrXAd+8V/35/ow4UJM1TZtuyCSI5cA336Emrtx0L53wR7Lc
WmvbDaDhB8eMQpyvpy+ygymvD7higIX1WU3OFqHTqEM2HKR7SVZHblVIjXCx2wDU
97umYXpKUqzcLa9yWtozivCO644RY6fOblxY4DXA4YCCNSXj9gwpHAjc5E7b7CFk
Pqcl+dG5AU1XEes6qZSawAHvQ/1b2oryKl5vadkyVm2yz++5WDSMD6Vo6sxD14HS
+Qb2BMYwsAJ/3/3mcF2l5gS9fKtKNH7pN9TWHeejplE3BU3WiX14gxyPJeg+Klje
8NnaaDqU8EnpKWsDrOmNTfTE766MgzJk5OE4YGRmGwIeU/4BJq2xa9kAO8zm6VZi
CazeqgqYxdIs+V2TOywea5jRmjqAQaIl52p6f6fJJ9js7hs9EOu7o4Pimp97Nm07
NtaaJZXuhalt4z7Djv4sDKVq1NjNI5Fo1LP5m7Mn0gJrFZvI2uOI5f4noJvjAnaF
IOCLPL9hZo/gdPjBOimT3whJW3wMB2FjDbxTZFDzhWC7sc6eWD+Mm3cYtic+kKto
drLrOnEEYkGp+tWIainZqnp5Er+Pam+Zh71SdDNIPzKBcSum3jx4z+2+ebAKvOlm
FyBZgTVGEXlS3UbT+QFV8pZfYJbKIyx3ROHYTqayNb4JOdJpBTVhSxF1S9fMHDIo
Pr05Jh7nhsvORERhVpbj4gUCjYgx9QGnFpzm5zG0OEns8nSYzRBEnWVX+Az89NtR
EYBtNOrXdmI2No+wNHFL0QsUszX4Y0d5OmSIVUoRwcB3GjyU6y+7PQ++y/rFrPts
MOsgxwT9mVxBJxHq0K13n3LJjTrOGSSZWxO4ldWDyIiz2e6HmUmPw9yNI1rf3qwg
f/LFtMrSnYmZp5+dV7jbAdGWIOP+VVSsCJtMwFmbvgE9QlbgOjjNM8K8OiA6yVXi
nsmOWd84F6TCvwMrfsbF6O6tBS+NPbENyeXciZljYnhg7sKeNq5OmN/b3y9v6okc
ayViM1uxUkPnog668iiMZ77zV2BFcrZQmaXbpTmdPlASYBYHRTMXqyAddPRX83hp
5W0U50pDE/YjveLgnHASYTj64e7yqlUfgNyvjT7QmUitUQrCxSt8u7bspcsizJCZ
kFJlAGk+12mhDDsrMnCUpBS5LfsAdGdtzYRhyyG7PGe0lA0IALuieW+5SxWxo8d0
5EsmgYWgTv2GxBlU0Z3Ect6F6MImV+6BrobnZSJE/EMWerH0rc3j9YysWwMPLYTh
e2PiIkoLT2cFOocprDDpFogmP0pQ03F5KcaF/Fg+cmhgH8E/GWL13aG7h4cLB899
sTBVIMb1RTMbd5Y5TiCGkCb7AURHtasRcSsVsVquprsjrucdHEO90lw3ikhQB8rE
jWLhg+iQex8zAziG4GUcMk2T86LTQumXa9RkDA8Ye9JLYe5bSvsOQz5IYgD9qYMo
ofnttndEeUfiLbHOe/O4/pfacia6C+ftN0PF4GObXUY217hrt9v5lW6iBJ+YKJxd
+C7g00ez5tTlbgoE0REqb/6GurrMN4prenSMhbsRPhiF3zjMG1uhFOZap/qnUZiT
DYaHk34uzdrhIhABombdkEbiVLSW0NOuI10rS+X05QxnlThV0u7VGaKImg4RI7Nr
MyxW2G/GOFrM+aG9MSmeKW8c5+CMvV8a6N60TD2UmdKll8iIJ4JFv7+s6ObUsPWm
EbaE4nHEE/merEvKyaDAMHwdixFX0P6wpaCwatRXMCmAkuhubaK+o1QH12J7z5zl
B12OBLqLKGXsgJcnAPzaJtIfZzSrOu+Ayysd+ma79Hv7jyVsUAxk+9ZOfEMU5tjZ
UemqhzlFFiRgztGBjEsFHcxmkSrZdyipAiAHY1bLjHLb01salYKIZZCTNZtkmhc2
MOsO8b1mNP3f8F8x4Y4DhR1rxFN/+SVQ8KP90SS++b+YQEdZBucdbOkt6RJq/xda
V+n0qRi/e2bt2+gpH15JiBjmgv6E46ae6R/Pqx+FzQU/UWGeQQM8U1C/2TrliMU3
SwWIyiFGxri3FRHzO1X4GTJ7bXV2y/tPjVRlxGcqqZ6KuDm8b/ELe3uCZ7w8KXWo
QnSwEyk1eee9QPrNHDVqFHk+YWG6JndNIS0Dyzw4LniNV0LOh3mie2PVoFo+WLMo
TY3BcjIdGrHIw18g+2CGJud6Ar1/O0RfLBINbImBCaw9GncjyeMpDR0TFssw7zTd
EoEJnDR1J2WmC8moXHTdf3Wp9ngTsYz+OxfbZ7EPCcUsGC5IvtENOCyTjNmy4snd
yZnJizyOz1d14pPvWuke7kXbSZwJpDKG34tSC9EddR5FhWZmIlQn9T+dPtsrTvRN
3OgmnxvSxpZnB8sUefJO+LAK3ET/5joWMBoun1Q1KI7D1GbAHZRo0VQXZbrk9W76
tVckBADBflFc2WLS80VcLDnPGIZaKG7CytyNVZ3l28DAT7ktZXKAjYGLNM1OFBv5
rE7bHwkRQ9H2zYnlXo767frzZCpm+lAmm2vWxTaqbcEW8fINSlbzVX1IWFAjrlSJ
EUu2pu1JpNXYwdlXRCunoBqBpAs6MkI2lVtJpRH4zHhlkGS/miR7vwn4QRsrRw+y
SFtTE7JetyFkZQJ35nLL1MkwbP1kJLHWppAmoyOmGhxFpjj2qrOGEOoWlE6/zGJU
uDog+m369E8mHSQfy2qEOG/Ps70UGi39pcFm+CoTnFoAFZJBEX8qP9U+ikWInTc6
6kzFZ5jztG2E9HLsRiXKK/Piv48cDNRia2svhKcnSQpAsRPBMw531SBvl9ZWWxl6
tQ950qTJzigGaExspgcdoNj8gnCXZUK9b3nST9snM3S5K4p4vpMsg87rAbb1rDX6
eRtfulq3Pzmjgw6sh5h4Hi5PeIkNp6GIhB5NrP1HQE2NJ0bGxz1psDRw1BXHYdSa
pTVel0ZdnSF+M0Q+44bk3D/S3wd24r3OGS/VuH66hW1dh0HPbWthFDqkwwu6W9TC
cS6ILx1pD/fxGasxEA+38sDL6FFCfOTbWhYg/aqsmGuoSMkXaKI/vcY64a7aWvKr
M5BORGoYrNYaiCb0/ajPcQ7Y6J4UGpOWQcp1ILORWG9+tpXqq/FHvG6+YjiDQ2OP
2odc6F9B15UzOI4U4xlSgKr3txAImb6kAGudHlY3SXH7fLqMrjv7QYZZtPC/PCez
rlKAtCzj1KaEp/Zcesvr8+g6jC61LOl1WClPJ9uOPTchasjP4kzZNaPKrdaq/JDL
Y/PPeLQDcXn1r0eEfkYg/oCHskD109TaGEGQxd5ITl2xXH1zGKmwQ6r3bbwMyyCA
7p5WdF2I7PxG+MPrV8fWUnpZ+NNSu+m/DuImDdrfQ6iUKl1q7GhDEl3u5MK7e3bz
442b8M7F3deiCpPk5Bf4SJiFupfNwrUTle6CjNl+IauXSwlqe7oqUXFZyRBGlEzX
+AaqEnY3nY1Qy0DEksk9jiUBuW9R62khhJHfvFDRPP8t1T2Vw5wWDW7wRUOGv7Ue
6NMCLw773y3UbruUbM+HHW0h+lgxasEzGhmvUEbupzemif5SfXscojY1IhIm8Ua4
HeNE2nzuJDsjxITubOAwvZQQ0wgNZqAZSVOYjLhQ+tZszNGMhDY8tKxjiRa5h4Au
/2MjL13NXT0JEynv0szTgKzbKu2YcvmFut08vZvHt/xqhLqkNbwfwDr90aCjqPpU
u+A+pbXibgYjp1BtWickMbi4ERHpsQKJCaSz/hcaw4GO7gQS6RbkBjZ6GzDcaB4T
glaRlxXCXfZMCkfZV7TU+vkhan3ol59w5mN8nco4jDtjjP4IxbrfgGrzW/ovVCXP
ck/HDbOMjoXC++mb76HGY52qHfZkDCyVhxTDzkO4Q4kt/7lwuxTuwmbiCP2IdIt7
GSdhPC57rc8XV2JP7Ae3Fn5+zTa6HvayLDVDDWOavqapPy7Ipbxt0jB4giEdh2EL
P2PENQNld53zeqayWuy9B1zjHK09UIMDle+4Z+5wBxbDWGUiuAYqYDjkSeFEeBrD
dMglFm/5UY53Y9tSlevJm7P6OJOJ8YWaGtyLIaO831EJhacl+pI1zv5kwrPl/neY
08ILUM82Lgh8m//4zc1FY72E8TwhLjNZqP2CRRBmrq/sTDwVXExkEydQlrjBiE7/
CaKAoyGMYGlmq/4kwUGcuHO3Y8xxRA0ZLp/h8R3E4VFtvR0EZ5zN1914Q3ExKoND
quaRLypTBcS+4ZEqdSoawylMIwQl2Lx1lh1eTkI3TrHB0fIpTadphP+U62NH8RuN
hneZwIrBo6MclFk5MiI/GJovEpGnTyun8xDlpN6XMHZC/jW1q+wXZw4bya9neD4Z
aO34D0BNLp7KxrZ1Xyc3OdwSHJGb7FMJYzXIfivUAzWeDySoo6ipQkHTnZNNtdDk
NqXL/eLy6xStuuKpiAdDipp+yRYWnK6thsbGAa1WrNG2Ce0wDqCGmb2VZ2KAvg23
MPxPc0o8qU+WbiZj+Yk9YSDZ+o3qKH/ZOLEObMz9yZP3yViw6TsqXoZDiLF7ZQTP
pidQNpAdNaI/OJU1w4t+agHIT2sYArysR83pUpLQPDxZ4Kkfr1XxVmFNNesw+lm+
NBO3zDoEKaV6OEMY/F3/XSTkhQpi57JlGdOrVw78XjzIxhPFXoLVLhCAE8dRlxRX
ioGyk0MaKOBoLxIAFA/hQzCMZqeod0/785hFLj/BBKl2cEiDPwD8F5kRTHIH3pA6
w7KsQmgwORNyFTyjSK3JyVRGjDPLu9ezbuSmCduOb9WPeBMpbhzEWF0EdTrwdBAD
RNLJUy1//RtcaET3BziVfKzNpPISpfSB0Vd9X1L6Ivp9ru5P+ZmaAKUzh6FQy4RU
B6eb55u80oM35MBpti88g6RbX0XWpFciuuRmFzC8nKB5bl++vTXQhdOKWjIKn3Pm
Blq3WcqWNySP3BqmVPWTqC6hxxN0Wfjg5fd8MpAe1MllPy75/Un9emGHYhDXOAn3
UXXpO49m59oHTzeIT5beBe8fbOWM3IMmXjdiQgg+0Lqxiwamq4uNehxtAImei72Y
mSI9AxWdwEllbUTGa5CdchGde50zg30YEIW3eqBHW0YcTuMUUOy8ATATsHPLEnog
1BjjZR5+4YSXE7N8OLIq1B9HTw+CO922LtsQoOel+J1tG4up7g12umXset6KOAEJ
I3Wt++I/5LHGS1kRww3c/MyeUDQ0nOo3eEGM9fy+hGL5RYFdsMheDJPKi245QUpG
TfeYbqt2DS06S3astj0QHFmMk1as/F9u2jQCOe+sQs36civsH2RhcYXdcvj9VLCw
T4SwlEs1Y8X6v37JKWA3y00IBmb/qXoYchFybcqkEtIiD4X02htxbCS02wDbp6fg
OvULxB3KbgfXiKev/kc6R9gNgW33Fj9L2zM1vLHXalB5+BGqduZospoe2NZ0PgMT
jVVEsgCeKKp+ujYFJabuy7mf2UVPx63Cf7RWMauJ3iUUVBbnI7XlaFN0VMudg+Wi
+d4wT6NCysK1Ivo3Ol62ew3/PAlmpOfZkGbfN6rtG5frxG6tB+PbKKymCQ4O2QBU
XvISkg5opi6TvyG/l7UUT+GtDk+EfjftiMefVef0NboyZvfe1X+oVLit2x/eiKpL
ItQaHgr1V34mW9FbFuImYewgZrAhtFyFFG63btYt3em8e1GN7k5vcOWma3gd7scH
Ggge2gTj6JphIFna/SWgL2j0SZp3ilPXwlsurf3rZ/Z2WXateRu2fKUvZzPo/Kkw
HpNe3pQHTzILdKPnDvN/3jeyBg/lLdyqD0n6qUKogpcxoCTIm/tco9n9BBeVKmB7
54WCE9onE9O4uvjEThsV9Mntd7V9Ajq9wv1ceLtrtttrJ1l9hMqPMMO83OvCtkc0
kqKZPX/7J/Hmbj1Z5sYhRM8sQH0mVcJ2qlNJnUSq5dWIl8z4mHTEOS1etNczIpBu
4/rbUWuF7CzDgSMCjwxfWS5reHcnyz669bIocG+pZRpZ7bQccwfyJdEgkUgAc4nH
q1+cnRvtoJwAKTPVqdDIztQo16ri8DvmfJ/JsqMVCBgLRIFQslhGl2Gnk4WS7l2+
BUNYuenZNj4rVBUQnsknLlWbC9bOIOpKrWjBf9BB7ZwmQMOincPcdYLzivomLgpz
v+jgybBddKC4FwKQaSK+SL8qLkGHsNC2xmA3fCO85ztcOExScTsbXfRdSN1W55y5
Fq5zeQkIjfaWGkHbL4wD9AjfdNMK5QD/edettAfgkZzxO/jDL4s/rGPq4WG4LE4G
hsZqIAe/z8TJK9FgoixbAbVhNFnZz/WQEwIoihPv3pu3+PZ9Tsk++c9koueowkX9
0az4JuSdeZgwSzWFa59edWX4e9N5ZgsCuF5lEXYQER6/g9tHWp72Vrx2cfoWGgqw
1VLYPTmgDayNZuBrI2KOSTPPusb/Y4IODxxMZOvvvWcgyzjcPHB16onoaircMy5O
/7juGSgB+yL0TtZ9iqed0rY9YUSoqqnJWaPuLQaDWNQjDAmJwv6UyJZ1/Bc8LIK2
PUgPGtlmpViMnaP/IoT0oFvPAA6Wj95ooJdZEBj8aynP2sB2INaYpxn0ggoSdSZt
uhWIuT8LCeggXm6lxHLKE8niEfmPleagp6OxwtfAE9TZAV7d+YRxb08XEKvYyH5N
apZvB+Qyu+Tb4Kh+DvGuOBALB6EvmmzI+nPEPP/pnI6uY2DIjDyRZ/qUNBTOa1ZO
E4RShL72U9GYrx79/FyKoudPJsLksKHlaFVEYG065wdiuQMJZLDuIr6BI1wGEqmq
OlPf9SikHEEBDla9/BV4TF2q81I8xTzkdel4JTYODlleTsYTUKfccIrUBUHuGenS
LEOh7NWiQ09gJitHn7vSfSq97cxHnYdsZzjxtpRkonnChdLD0wYODGK5ah/8V1JP
r0Wn4uWWtRfZh+NqY4H8z6GW21Q85jhn1jRNJ5xwPAEfzcOKcxelkdlmPZbyDxJu
C61ZCDLEtq/WDCdW+elKAv4AfxdWbutemhRj0PhpaYXMPsZQf0GhVbXPRJYfdziB
yx7sppLfcbjKENMFk05+HaOHFZmVMgdGrpAHXWQrNgDQeBSdBqOens5I0CEXsH0B
oQFRscVcpGgZB8MtkelfgkoCV95vpI2TiTch7IEvvG0a+rqIKxf098XC5jSBOGW5
NU+GI9aP1jAb4XBHHECgCVpXmN8wBBC5grLO7Uc1kztlx0M62Be8LaUP8YgQ4yyU
Chv1Zx1NJHmNGpRV87r6992ziKumKcK6RYMuknRN5R9C9zVwA66pzZ0ThmE1fO6d
z2upDwgE4zOECnqGqYHQ9QQa6s8HPO5BnWaVT1UziNobANzWog1JOHIRyr3jPN7S
WTmpx5BXW+9+Gvuf8dGRAsLiS0Ab9khUk/2EU9yrhuwVOsUvUA+ZQEsrXPvl/bpC
IFOem3RxDULpllfi/zqa183Ie2vsTV4E5rz7kTiXvtjbdOlRx+7T+vQFaS6pFiqM
upyQ0plkSdNGkdb/GF7slkyv3Mu+eNM16swftA7Nz3NuRi8PFgPDGxnYH8aXIvOM
7vKeJipgeDfngnDBbgrxZauMhC0+TRb7LGVXL6puX2wC3ReWrwUi3vcFkVOx/Max
+240a0c5zFIjgh+ve+29qikJS401Qztg09yP+FToFlAnDNjvrjry+VCG4TiTcmCr
gVaLr1cH2KP4Jx7Zawn3r6HOcUMAqcOdwS6D4SdW70vxAeF0iJcuXAx6JYo7AVVx
8GfwCliBjUPkk8zthaa2GxR6eI28kcVHWG9R2UbVxHug9Uz3MGRfynyYzy5f0/pj
lXDpR3gntHG3/OJ06J4h0aqbClIv0jr1FztzqmSt28dzc5IrjGCNQI041hYrP7EG
EG+S+Z99ppc4Li45SVvgmPOH9Y9Na/6ZU4Uc/R8V7SWhhXK2+wbCje+N1JPnt52S
UHpsC8VNQp/WXkp/5O7uDMJrDZ5Y/EY91pK51Qo533F42JQXCMeXvj1SKaQaL5ML
004/UnS+jdZUMwBgbYP+JO8yRqzrPkp8A+ku88jFZwn71lqpC0l4kRwZXuVIvLVf
I686vaa2jvkfuoF04bsV43/UV1BvqEmImc5Js21mkyRemVBX4T3EgdSM3wOuzWTG
srM1tIT7o1AGmlKs9Cpq9Dd8KyrUELyIqqg+Ls0DXOJa00u/kb2iY/f0VghGmImQ
c46TdfEBMyUhepDMZ/MC/faNz0Q4GmcNiX1phgWOWsum5EDc8lGf5WTYPHa878o0
ftWgjxyjjz6QEpWHb+8/e14z4XVfclwqQFCam304PZinqjQQfOD0Jceh75b1wYyI
Bu//se3GVkJgC4hry6TWJNvhYswTvkMtoMtMw1kMUGEnNhYEwD2Fty/nLV+Kh3qm
sizi5RuoKUEHDwgV8r7Oj3F1Jdgncr5kJuUc1ykX8+6DGbs/AkEuK/2agBKntzdU
zWnT06+z5iURibq6DZiOJ+sx3Gvk8Fsn5AegJR+Du+7UKrs7gqMV1M0LMxEvZiEV
xM88J9i8/LgxkLY6TBQmQyp0Nb5j+2/iepZslzDkVaxH4kXOnqbZKo/cY4tIu9TE
02ciVNwBp/8nAzgzHFizCXW2PtdOwyryrHsiJJt7GR9ugU+KkOF5+d8c9qIsEbqi
Kv4Ll99ohe5RqKg/5nmyyEDaEMF9GXb2b5qPZMleWEubFUkgHDvTQ7rxWMomxjTx
ybZrdxhC8Z0c7UDNNXLyT7vycVdRmSQz+Ft0QEVMyoDhXODpZH+R51EVCRc8oj4x
+AFmIm5LmJx6sdYL8tG0ymk1KhgjSgWuzcEL97D7x2aBK0SyYWFOlYlB93i6AXP2
17lFJn7PJVJPNX8H8JPsSSDgx51mm1jORdkUsRt9CJnnC8PVOiiRR0APtGVYEurC
w1Pf05cDhZhHzrKxriLo81MJI92kX+vwjAx+TRx14s5Cv3zmsbDLrdrcfh5n5CBi
GVCubbjHVzHGcQMiXjeNuO/Ir0QUSfa8mgPaZwV6quDM0Udyk3S+br7xh5E6uG6Q
mBIKNNwn0315kTkOMXuevDq1JvFp+dxDhX6c5MV7ARJIM7tS1eM6rCNmNLhMcVy/
YdVsZeDIi7LIJdFmMsuMUXye9tGrkcKrucsh5UKi1BYvB4nQgKcOySIHEP8CE/dn
XIuMSqDPkBda3iGoWne5zgRI0U3Y/xr7unqAPVvHOOwlZ/0DHZ0RDbDrouoxFn5V
aVF1JPWFeDfQasFJsZeWzpiFUhHyEO6RdcQo17t6oDmncZyxllYfPZVyda+nOI5Y
qSmGhrkjjqTBke2V8517noGrpqou9ZBIz2+dxflaj8ErSS12qGR3AaNVlZc/iuvb
Tl2Ock2cyrB8G6wKg5DBuwVsYHkLpXVTH1MI4Yp16KsLC01O9UIe5IvexL6aAdrJ
RDvUHy2QL1Nj9SZ1rVH72RgyW3j/w7C/7lSVcvruekJcCauw0F6Q02tEpchX8o/7
ivDZkFiV/d1EnoVpIXMUZLZoHfWWYxgFVWZQDbcLS+p54mwK+F37i4DhI4TG2/Tw
1C0jDfOmYqCjFiMCJ/zRsHA3E6+7jALGTFf5hychMxS0yESvX7ZuxngZDTdydluI
X/N4LGGs7INhKa5MhCDvfGreuBlwvCeWRo5QWN27qbngm90VEdwxylsn8n8jznDr
pHDoB0cbmUHI+onIPDJNvP2WlJ6tRmdZqhASE4Ud4HX+xJoTE9Fste40ucuZqAWx
DJorEO49ARTG1QizKzZNO1SUeCFPztJfIzmvy+orY2YMDTZueiMD68IzR5BvL//Q
07D1cE6MwtG7DwXQl8rZqOoplrLDam5N7r+s9hQBzZcO0QtJjDybXe+29kJpw/98
sjNIM2FbmuO6fAjbi5qmC2rA1ZxDW0U9rzFXInFkt6mQOb3TqOkfypXI4KjVXg6u
3Y6HiZez1/iSrJv84vZ/FfFCs1ZATgIbF6h7sWbRT+zoM4dD++AJ85lAaG8lvqJD
nuHWJT3rLmfbTB5v1Zls5gEi+zCPI1MrNZHu/eIRmXj/MOfYYGlgQWpC0d0i3iE7
ke5JnYNjaTunOd5aXJ7mxsYDYAGB5sB298kxrA1Dxm4mKJHYXfU2GCh5qFd8CdNv
g/SKtYarkdRry+vDdUs5WpJFPsHyuZVyqmjNuUhlB103rycOkc6juSfusnJ8BXVS
2NiYhpoH0u5HhJIwXjtlNTOehzOvUmwQhDBpoqFthapivIoPezKHQW7PevPmxuGo
srJ1lLwhkGkiaIC0tGTzLo0Pv57gxYXwuAUrXAdDziNtMpqJmmneqlG3XjcAd4+f
2Zs0muaDniX/gDR4+tN0B46nWkO2xws5rYQtvF4z8/q106l+Rs3exhX/MBQWVF5J
Wjza9dllsH8VHCdUMQqqFr3Bja/1Hnt2XpMxAC2lrEt7G5ZV1hKl4SZFm75zuYPx
wdZZ7diSs4cNpjoAnwhjtyLZY13LNpjRnFsJhpOY8ubJP3aeiadTfwMi5Skjo11U
Kmcb8jN0eb5qJ58UeUnEs1vu9tHxP0RsVZxMLTgC8jR1EuBQihDH/to3UkWhaTPh
UG2BclhOljCdQ09EiVxXiC4SBfp5z3bRYpOl/lTFR+OSEpWELaGhXqcTP96Th0i6
0XiE4yZ7LCB1NjZi/F1mhzdklEfrtsifRUBCDlGe66LhXJTotYKgQoeCw4X7PdpL
Pzp290uyPbUCWqA+1BJNsFxXKoVvvU4DZSy8oR1x8hLFv0qrNjC04ZTMdoB1udMV
kaLWvJGZODjNeSXN8JBR3TbIila0AI7CN65F+sJFqeEQE+FFq3QSx0X/ztlmxqdJ
Wp98RZR8QlUb2BtQtSlokFZOXvyFwlxC4F8o3TX+JgMoU6UelNMIfWZ9GFs85Zb2
LNx10IOh51mxs5qGAe/q2MqQXuo/I5ALsE3K+8nh4TTBaeAuIeQ2w7YFpytGaY8i
+irg36wNTaltogMysdAylS9CJZL/K6Y6aCPc/VBFg9ll+Nhuki9o4yuQoF/7E1yq
+mTAddn3iE+IkWYu66oGFEb8MpCLyQOVRmesLzRLuekEwfphNXQa/whwt4M3SbTq
FaPKeokv8ONxXZeMyP4YWY+fBKj1usU94nARQyH76t4NAwz/iveaEOY7nOac5TuF
RUyZnsM4yYqMnfVusk48yJLNoglelOYen3RqDK33apW6S6YTe2l6+VwuH6TXY28X
cznjsHKPxEZvrYN6DDcGc75uxfB6E7YNsm3OlODF2X9OzytcJTiMHXp7Jt0hpPYN
JcDdkCMyyIEQGWpKNBVy5pR5ZivrcJYPIwwDLm4wk/5Pi3d5SfH5+41tXvLH1Z8T
4R8KGZ1pGkPJPVXbR04lQg75IBGEO9jsJ3jNf/wKnZgOI110XuQlN0NIJ43ZR4q/
Ioln7SV1YEOEnjfQuG/+WrSE/b8JJEj5KruxEfbtHSqEY2976qdAM9L2RywbSes9
c9w2X37xAd3F0w2hvMcMl/yP0ciU9OlFf0YgqsL5ogktJQooVhgzmR93HLUptNU5
Sj/5x6WJyfkile+EWCm6YJWJCJaE3e17M1vJm1QhSE5zqESFLqEqts8YxZlQDwy/
VLV3WkhzCuSf6Tj2DYJBgbfiUa5aG+x6mYvZKqUWcNeB14gYMRGLZXd5uN+iqXVN
E4CUiKhtLb26neipgv9lbWsqZAYQ3o4lfC2Twd9pssTvjl2qFe6cqn75S6YH0viF
RqJrUSEZJ//OjztmQhaJ0PNln6lQKSCKhUwnHd9dwvKdKsbHQE+83G6qbGZSd5ib
u/rjGLm3lhLssPgjsyeNaoy2ecXx3irZzqe6I3Bem2bZ/40nSS6wC9m6mWvK85LH
82qK7WocR31axq4RS2FNuOv31HJQ8790Ltca1q0AsRbtbsBqL3Wy0WKk8EtsL7p2
jd5eOHs2ChOG9f4NT6j6etVFX7fylfh9Tq4M0bOcxD7gY9Q23VXvE3ffQPgdOB5Z
sBSLay26S3Qh1Bkz5BPm7h9ViTc6OKJ1xM51DFbUFlodLbO31Ft0Eck5fadAiFFp
UbQQPAUXQfUqQeObCMQKcdbJ7VrkM/CjEAoHsDYwytVw0x1w6DMkRvhRj0o2/+RF
2uKkL4zjFXjaW36z94SU0YR0Rf41/YqDLYnBzv1ESAl6U/wJCglEQXvEcHqOGeNJ
gbspHpUMHMco54jCD/0NRTTqNBl2/9FlWzywBSEhVQzJnU8hwV4h9hzCkbwZpIQK
0f96Ca4tdbskwO/SkYSjOYg9cWtoKv8SqU5Ptf1RLRBLKzTr4Fwb/7TuRjBRzN1Y
DBZ2DCkK3hr8nrWT8lDCUpcaeVS4oMYeGER3QLg638JmqwMe21igAH9Mu9KNMw5b
+SpJ4tKmhidJPbDdaV6c9iN/G9oOUgU4rbP1ok4hcnKUEvjF7sUoJjnAxYIB5grF
WfJFh/XCPuQfSPt3DpGJ77GUbRjJ34HlEFG+bcAt+XvvFnhDdCi22oWxD4+wSSUq
aeY+j6xHTgubt6C3p6XXIVh+UQpzktWiP64aJSc364tp0lDHHC3V3H64OvXXy2cs
4+v0GnF5nlSW09mNRVbJ2l/AL8ii5euqsbpeMZKz6jNzSCzBIBBM7u6FVIkq/r8W
bGKzuj2dOwpGQXoCPWHAvOTkSTwSZlRUfYHCxEzsskpIl2h6wQNEAc8pU5R7xMuO
oZ6R1LH6rf7M2Kl21Gg+aYjVJCCkOrvOe9pJS0lEJnFl7sS0W2UXvTZm1ZNYDDpS
wdyps8EWzPFD8XYZeYKBmFDYLScsY3yrYL8Utq76weZ2N8x1iwNbcyyYVMmal58w
4ZW1Lu3bXnPI/QscPBvuI0f9D7zDgsPfBOiaXJCErSgSJU18kA+NIQkdjbbNrBwG
A0cJ/Df8b7ujvcNmaYBoWT7hjiTdiMkg2vUci8nOLemUzqI6sHohfdwSfXqIVH/e
zDFIOk3AHPFIv2JMfaogCLMbNCyyYGzB5gnkrlHPg/Uk6BICsKDNTL9XOsH4s3nA
928hrYecvtxLj9UPcNeXxZBZQdNOCsXZf8jUw5ZxYscSMFFRMN3kMrhTIansuUP1
ggOeJV3550bH77stN0rxcK+pW+zEHWuSVQaedTppMSXQEexPhryYp4GenHRPQQku
Wrk7m7uMUFJKNLGJ7GrjTPnBK4JWgmHpLFlJ385jFA0j3vsILVuQ6VmwBm9Lcbu2
SYHJFVaQqUyPhZiikH+uroobUvX7RXaZkAXbdxJWfgzGpu5KbrAM0/0/QH34npQI
xqL8/g/KrnL3H89NRR+OKbTraaq4Q0PwvqdbZX1xuKmWtOtdK8xSUUG7VFnFzy22
KsSAXEMEMX3lprrP8Hbu2eaf04k6pWAPLUl+ITc9CrVE0gWDnrAMuU2roGBoZvCm
oWTfDpfSDtSEfsXvs9rzP4jqyh4auCwllTCV6sNltM7joe08ijzxv0FeXQZ3bpft
J2EQ3Kuxb97MM3Kt8PQD3RDtLiTWu6vlD+J5QrLlvwEIQzlxI9d+UKBI4lzV5a9Y
mKqr9K1lKteoq6E4Pml8h91KNTr8q8RrBvvm0npuxMYtRaGeA4bfHls6fieFnzQV
BcN385MQwbnfcz5o2zlXUfwlVGHMAXk5Kvl2NMofT0A1UBaZ8t7M/8UnL9WFJy0t
B6f4e8whm0svDg+HpOu7V0R28brzbllViP+nboCE+9+BP3UsVBIK4mM3XB+3yypP
9cLp/2G2WsH6zufqSfoOspgOVpOYGN/i6P7NfUxsGGmmUxZHunjSzQvlux8mI/yW
yabh6eQvszgA4VCxXL1Oy//EdG5nX1T7SB3Ju19NSHWOQat4jvRD28mRrIzwys91
gu5TxX7igehn01DFz8sHlQbHBSvbPgoElzp7766VyF+k/ELlms1pepnbQtRKr+YO
OnNX7Gt+LHXMKDV1w/4UqirqyS7B0yvo0AXVDNORfGy0/XAdJ2oTArq/0GU8cSHy
bHSaJtrIBxsAmb8y1rP13d0gCgHYxP9oE4Pxt6GIe8TAuh/ryDcb/7kHnJPZErit
O7e3wSFAm1wuHY91YuaO1Fqb4cGjd0wWBx1RmRIJ6Mn/vz8kcJTW6nhOgp4KWjt0
rdmYFHVfOayIpyIW93U+YPfxSmpNLv38cw2KDhRyfviOhyEOUdXK/AfEZV+p9Cxf
gqLaM4IcGfSMTxQN8EJyhLitO+QsPSocQwOb9hADbhLO57q3B2FS6YZnJGkqbwU6
rQtluDgzKNce2+M+KcnB6DjnSHhNHOfsEsAPOkudhF6dt0rwnBcXUhcF2LQK+0fp
rikkMOxRMfP6fl9RGavnVdvaQ+TogyY6jV01lDt34qWkYt0Ydc/3ofqTfGqEjXMc
5h3491/2CE1W+Ei1ecn4n06UL91w9yvv8Lrd96zd9kkfZxpjBjV5hyZyM2iDL3fz
FPmLH16eZWWq9rnRF7uaXx6iSR8dMmG2RTDLlToXEGQ4yb48Gqb+cefg5XbUhZWn
GlMfPPCVnNZI2hzyMiGmB8X6nbV/9lajMY4A9FXLw4NiukUT9eXQwkhdj/ozQKo1
dLv+zK99MRiLb2dhAMgGg0xfm1ddvfxUI/sFFP7c8aj4U5x4+ar0q0SiFxYDMDAz
OCXY5PLnBoGCQil/q8ayCp+OCq5Xexi3T0WHK8Ok0/69n3V+eTqlQWHWVgs1uZQF
T3JCwhn13v1qAJP7HR5xxez4MWCX3vkkJbyW6Bep9oUY3PqZJto2P7xcTAKTISvo
ShYWwoTR0TfKZrXORAd5pJkB1PwAgBkueMQBWkUavegkVYtLfh4tgzAT9OqLvPtN
xVZGfIEYU/mHyPcyiNuspk+YL7Jo52kyEr1xwrFgKedmyVJ/ARCHGonWJCn7yN/0
oSgSRiW+ZZoaQHnOZJFOTnNDnVd9h5bNu8ZAmrOjPwRO3zwQsILL6Tjj2YtGoNsQ
2jigSrsH0cP0ESt5Ghaq8oKZn5T8r8ZEDHbH4kHYSKymH/ACDufBU9uQZtolWn+T
3ot0QNlPtyGsBv5meFnFPeVxtgYghIwbyGRKKaP5i7J/BKLf7QueZwcbIo8A62am
J5LzU6lyC2wlOPgX3yAE3ySkGvP2iYkHztDVG3vNXqR9nBOvcgfoXCP+/tCngESq
u7Sf4Ds6Sv2scCJ6b+YIJgl9p1E4lOse0epGYPRoJaamxmlTVOWrLYQD00KLXqWI
0kspTWmZnR/hZIqYqP+bfkSXdUEHAvGoa9d1gTN6GaN5/rE0UN0YqXilMPsWt9tq
hQG2i5In+4DE0iyvEx+4jAefmdRwroF6Lla0GgrNkt8Iun4T602xagPGPH+x2Unh
cTsqoTQq/sCelFxHMY1fYY1BB8yffLwIJthsXx4TaqNZiVL1HC248i5uMdb0vwzy
OBTGXBakdYCuiO/TkyFe3tFNwzpUbZ14KRDt4RLgIweSI3tIgFqPLxksbq7L/zrw
tng7Gpxf+v+PPAWE4EUVogW/bpT+snTbs5HvveawLgrRz1RS+6YxUn+bj8o9sx22
aLoFg+KrRwWUDet3j3RPjoucm63C4QZ3Uq3ADL+1mZa/JXSns2+bineRNdVWNogI
XNtrflXfJJN9HKFq9oMO332PmGX22F1kIdzynJ3R5ET/sV6zBLUXNCafe/qRpMra
JqjWGgWQ/nNRqyDqNMlfhlenXhtUUy3gEo1Lezbw2qMIEzqT4335UmQZvlcOq0IS
+5borXqwXWu8HJUHTwSeoEG14khDlAHkRlhlyqBgoZFGPTiktbpkmcBwN75duF3V
KDCeJaELgJM6BrDt4JxKk3OpuEMZMXFER7SNZV0Gw/Boluj4Mc8x4LesCyZtO1TA
xP0QRriS5/EPQkSKx4C6elZUPgXsbpaKexPtCW+rlFul/FpzpiWQ9h2bUxmK/huu
BO/CM+U6rzOyrGYBfCQBVhDOYQq99ky9PRGZV6O09Ri8Its2XE7j+GuKUqfwncel
hq762TNlt6cFM5rsLIJ8fkIyvDYA9ndHcUuLg5iyDlDa1brLMvUVlc4KQoj6Js7R
am7mpl6D5kT51brNvymQuiPo7pVzyFi1dSoY1TQgaLxzV6RaOaNU8nZ5ZeUhk9Ht
RkGEvhkOK0zvK2VawabKaif0345Mi/MpQxmXD6U5MqPr4VM8Ez7XFlTTFnltoKPC
42LhfPDgZBH6VfNHa0wlwMf6DT1CjNGXrE9S6GF08TFXeaTdRU0D2Ap7OB7wn6S2
Wxupdmbz2rm1gE1gdnqZVTbYJMtZeIMwCVzah0V/Rdcorttp5vpm1sx/sc04i9Ze
b1edn6WgIjoLJPmHb8brpcZYOYwEokgg/tRNzk9vQQAkPEDyqxiL1HwnEPZoIOTr
fGaSJLXRAHWUms0bK4KsAxupmohXqdHfoZ5q7OeZ0+auLDmc7Bej4+16bsO32HQc
9p+O7KMMkCYOkLbkFT5uOlmG9kY9W64u/eTQHtkoGnhjJGpjQUjIRRbrtbAgiBpg
kjs1eDfM+k3lVH3o4tHhCGLA+3SHGYvLFOhMX79J9yL0dXu0Y96zvHvrIQ3DmTnl
qiyLWg5amfF0NMZSQseYTlzwIpVQDo05utCf6aXamjOedilhtLN9bwiZyIBkjMTI
hdYN5s6xMVwLJLkRs++/QIJoqc75VdWzcp9qm+vwiP2p2z+vREr19jbvFrqokr6N
Hv5gAk0TkDMsSAJDyhNZQTQgc0BBUvtwThdWtnMO5Ht1oordh+CTuzXwfZnZsyCx
uXHfYAyvTVDiVQQ7Cr7ukkxfzewCodHFosWTki9QKRD8cBjOcUrHEPHww4RMR7LM
RYvK+n+0plORhFtki0/Enck7zGwNjfbwZd9ZDFFgj8CDKSkL9aTzisb+XEHquNGM
G0Ij6lJd+G9UM8FjmooZX3XvXKMQ7dlnJaYSQxLetfAOIPaD21bqovrWd7dLsuL9
uUxD6dGP+e7UHSmragkZ6a0y/CtnSBJEZ5VdgNBQFiwv67dxLfs0d97DO603S7yC
v8deZoG+ZT76EXIYv5oxgR3DNs3Z2F92bVhL4DfDC6fBj57RBzz9ZQ1cq+NFXD0B
wzVLh04Hj8RuOYLrr8Smb9k0j9XQ94E6+6oxiGDPcYxnYVMwN/YL/4uO3M+FTkh/
7/EQfyrHRezetVYNy3JMTlF7cObVb3uPkFGSJSpLRpxY0BE6wum8j+yWrJUQWX4q
qSS+6MU0+TMDjjtz+JTuScrH5lT7f0ftrmyhCcnmNvf6xDnRWAME3tLF/amlpam5
Ao07E0UT3qeCGWWOUFD87qz/zTYDkKF5K1Y9T2+G0PjKzvKRvYg9/TfvTPxSIfTV
ic4hucaJYe6XrDJ2fH1PCuMj56bKnPD4YZbLcASlhrb6X3r0fuY/W8e1/xZmvLpK
Bdj3vPFfxDT2w1GSEkMa7U0Y3hV6M+r3CW8XzFoixIynXV5tytBdd71tFN7FAPuT
cIKYafPuCqGz8g4nzutZWm+c4CpWshc3SDAQeXDIwsYNy/13YtQgMUoC22cB0xjz
A0/Uo2aNjgihhPk5iyUglG7TM9Lq9G669NS4oWlbcDeIc6M0Hr2BgB5CJjA78HFn
TjgXY/CQtfgqMQz2E055RlfUmDoheSSzq2MvuawzRaGk8oQ9U2cGoNasm1j9qpHq
N2DCaHcn538eKh+A6wHSjgFZKTTtSomWroMHB9clGn+TwtGEPVsyaCYuz4Fz+BhT
q8nroVQTPHfa0cVxaXFgO6M+STnxtuqWzbWLR6kW6B2S7Yrgurf7Cs7fK8iH3bE/
mxXRZfJgnoIG0foJYGaxWFpr50NqICC7YbcpVGHWpB9Q+H1qrj111eZUpZuOGaPs
m9T1q+/tm0Xntlt1zx4mAgT1FXPpEAgYRX7bPPPPKmRYmmcA5qdh+nLgE6hD36ha
iUIqfUIMKwswgpKsJ5wxNnfSoAF0oRKfbOJcJCF1/mT9bHtE6ZN+saZJWrIMWJD6
z8r6huZfKU9dDVSxU7aKGnfJyx3sCcnbDMIkOvZlXl6826dmExGfuIpHil8J4a8c
pB3aCBPaw6DsV/YylZG0ioqna5kn+Uqz/jTOm7nfxLMlf4kIxG4btwGRaoOhI1Qj
fK29ldLjf5rdo5pY2LcgUMDEd37n33T3xvWnPrhuxaR4MnhwYgm4agPW56i6JIYh
ynjF996hT3UPzB4GzEMaZwyW/Zq/PWbXoGVdXkTkU9AUi1CLq27ZeJcF0bNCj/bF
b2mAQhzzNcoC9VrRbf9dB/AwUS2ex9F/mvBiX/3kGmTY7x05my0XoK/FhB6fmvmW
6b9lqW2jPsutfnslsjymqa0U5+ynmtQGid0P9gfW18yoDxSfHXbB6Cb+jkhTjyzf
G5MnUyNVxb3he3vixHwsoCp9PDrcfBFrCzBFsx2l/4F94RZlfvT9C40XFrzgcdAB
iIrFynm+RmNpDBrUCYfnECzUTQ3AOBLnqNiFYL3mC9WsQG56jwnHb9p36G/e6ar+
`protect end_protected