`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 43376 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/9huKRhRMtvnNqb3Z+UU7TahEoHV+T8U3P3ufru7l1O
3DlgtZzb9QxCbOjthp9+wDkjygH0eUfDrEl1ovhZG63Ku5b1qCWWsCHhgjNa6PmF
dG0qNr4ChYrOBr9K7ebHIIvs0gfniLJB7if6rYh5ruVjT2lol7bjjKoF47ADqUCL
TMagZAqDAdDnbvn1XOIPqMpHgiRuy4B79kxzjtRAOw7jsX0OLxcsU3hBcWZOQQ76
ioHP/ga/QoHdp/X9ReiCOfA9eslnZeTlEHZetctycLjd3/qULzIbwb7ttLRoJ85h
2wdxlWowhsE8Dg+WRKcZja7op9zd3PfIKZLEjuajJEc3v/HhVtkXMPAwRVs0jyzv
Cv3z3VjPeGlA++q0L8CZIkPRl0XHRkBJg8VOYrD2cMXO6my8KQxR13+qF2jInyhF
9bssghgKrQH9a88My/+3DnfiNSMK3r3YOmkEdzgFlmdt/YueewzunIZkFaYvH9Bz
hUgXaXRw2mOFMbfaZ4hfUr2ByqPuYI48nHXvL3uRnzKdu7XZF/xXCDx4R8n3RL6M
gPHqfxAnWWspXTHkyWstCSo9WrFVkXFWR/c3OwbbZ2UCv2vEF3JiHpFVljtwcaDI
8bXAHkADJzzbFMlWfeEYujkg81t/lRi8SWeUGlBIe2y13rLuFXQOhsZzkUcuPdWM
tPeduvX/B6mftzR9PPbO/ZV27jMNlwT6Gpa7nhTb4OtZ2G/m9Wh4Aabauo35vPMT
qKSvm8vXiVrQgd28dldpAcf1AHgTnEKCxAimszyQGP78lrS+CR0NYTv/eliiYEj6
bIeXv2rLP8iEMh+GIfj/JbKkZRzIJ/DLBhQJLh/densXYaA1n4BTZIKedqVuTzBQ
P7VnI8npkT1k8fYthrWJKvBd8fAZqdZ8b27kpytr1L4TQuywITGo95Z6o0GoCf9Q
Qfh6CX1jn227xqWvnAh/1mIIYqgM6LwRaCPgyiIYICLgOQuT4dW3XkExAswk+5iM
t92QVbQ28qt4rlOEKgisYTZkXqsCitYrkpNl2OOtiL3owYjidNdo9QXdzFMBfps9
yMDFID7sKRIt8A43b1fcKKsztk/QjmucjYKU2ZTe/zA4OmlLbZybH5oVrLv8VfX7
ustUWA1RRkB1jbkwTgMACDYswiNSMc4P+8gg190zdsJq+xPoMw6Qz0Enw27rkbo4
NyYiDoeI2KYVm0ExvgHxrmV9aDqALdvtHdNNlDrFPF8pv9gEJPnntyrdR7ictJHv
cb52OOP8P0NczUbV4irxi24ea4e1ltY07JsFXZ/6B6WGTfKSH2OuwLPUxSxLuZRD
od7Ssl61qPijTpwMld8fFyFEQktySCGi2xsBJfrTPVJE/G04giuEGl4ACJsVuDYA
INOan7dP59XXwV9VZnJC9OEAWHqQxenzaw2fnJnBMjHSrfoq1N/A8QqrkvQixpYm
g89sdXOEvHAxyyDVlK2XL7AnOsFGVuM4EEVgvrmtJ2AlnFHuJdDR/3saacnOy9js
Edh1mKqoVqhOf/Rzd8Mh0EDvpS9IEE/+N4LIm1GfaJNu0AgxbkJX7Ihm03CGmaEH
+hOIUlwD0o5wmGTF4zkTB7K6XqPI2du6uBAAtcP5Ryn093mRiGDyCdNuQWBKYSse
Bf1Auz3kVWKjMhOBSf+/y1W13pq5+G0ATbojkPDKi1gtyyHDPCBY+t6LA1o9a4ew
X1UEJl4/7CTgYS1q/Ybs+kFU2PWSvp2l0DfFwJhtrVzHxPwFGOXAyhqmlYPglVj0
uqqGO5D04S7FjI3yzYiQCGz5Ctykih0lIBzl9SLLaplMHpvJ0oLQjK102Lyn4Q+k
1dY+rA36hGKUKJ2Spvf/QtQCOA++GsZ7pv9mqrd9j8xvEnxUOnMvV8Hmpt8VALQd
KEaOIEvLNDnfhQnGIM2Co9Yuia61RYOtqlidDJdehqH1M0CN/aHsey5cr21mwbNN
iowfUmCVbIt1NKBqDK+OoNtqrEUr1g2lLme7zqUAi2/877gH+q8BK8HAdBbDDZK0
KAC+Arr8tO2KFhjBb6CkKpCg15TFQDuZQu6Aa8GwAWjrWgt0o+wzb4zSc5gCaC6x
jKWrRl4NQZ/C6eiHpSrRmE1vCNZZWMca6vYyWXHCk7QJ2Ibda8k2HnVRVxiD30Es
iMn5xMYXQBv0RozNyPALTFjXqZHjI3ucx8h7TRs7WTgoVA/gk+rXv1eT4Rkb+hLO
qmUqVb8o/oUyLgYIQjT3BN4RMIAhbRTubZIAF+JTNE3YgqZZGR9r5B0OO3oU5gxc
DY2mZN6BAn6R5pYOQE441c/mK5rQ36YgbXOIXGO1hgs2lHsXSV5zbmm86lL0/ZgA
yPadhvFBOLzDQB1HD4UkpeUtfJHnacNlsY6F+YMMoMMUj0ICoaMQn5NUqqg0UR+V
T0enQXndUU1CP5gyvhI/7gzjCkhYnu8s+4P1hSGJ3b7VHOVyB4PB/md4w/z7kkFO
BUYD/1Ly06uYEwtSjSReEeP6hc9crwJXy/ZCwkF9F5HL+eiRCFA9kN9OB/eXr9Yz
0aZe/U7l4oLcRUlNUWRaMKXZRyQ0cAoRdtiPwmDTzackYPR7rqq7xN00romXjeyy
9tmhv9xejuvYjuEjOJRQYVKOYzJTgD2/Jm+LACmqRXLAjQHMm0bSPId6C4ovFQRn
4WkXwsdu9Y9Sk0Aax2FSuJeAqGKghRrahwXZtwLj3L0gN0zplk63+kwAoHQo3q+L
tXehdbYrPgUZxyDg8AZGXCdjupG0z/ng3QIwT0wO3eK0J+wFDySEnuxSR7zv7iWv
usHKZDY8nopsYrXkLdgUmEbYGtpOYMdbx1h7OcL46lhacHOEb1QcrMtWMi3Q7Gyi
wUkz30xf36qlDOkKTNig/5tYq6cMPxmwdjS7DOVuaYY3a3stjUNVus5N+JCGTHQM
hFQ+G45G1NJ0/rR6yMYCxjyIgKaE1hx1JnqwX37+gfeSwmfTxFcHe32filFcm1V4
VQ3M36ooLJOX8e4gRqlvegnDKmX5MFEdZPqi01n3SXN/yEfunlkqXnK6n2FsRAWv
zGLBx6EI4UiiO78Cp9hYd4YbRQbuKnLTy+ino8+baHukYk36crBdn+AGvE5n/2fT
WBDf+nrX4c7uAacWw2t6oEoHgGdVlGRv+QnOvV3NjBsqLAaL4HtWVhzQOc1TooS8
fgr8M/l8+P7nWA/fOegdwQuvtMd4Og8yQ3YOM9zEda+w3juD1ebKmDXQUfP/Lch/
vfD/sXETKGehqw1OjWfJiyFSfDjkefJE9RQJAlby3YQKo3qjLtujzx5J4BB8Ww2x
rEvPkujc6w+zCN4BLOTqMf1feIFtRz8520stLWQvU1LUmtlc4onA+l58LEoJp1tT
kmF3e/xoHraqvnicSfu48d4ExQ9oq82D77iD5+2KQPa4KNPudKnKGjN8NA0QeQBR
nwIiAcQjcqJZw4mHfOU7mbyidfC+btCHVpOzKDEPPKVU23UFfm5tJXTJZCG5qnSc
NONjDakaqjno6uuTY6hYJlJ+QzM2VltmgP5fwdY+tgzPcbnDa0SFYGOgwtRPzVRF
Etpmv7FoWsZtO8NpFdSayyfENQjzDkyFahAy8M8bxG3VhDm8N4D8CZC3sSSVbRWs
S76+rKFff8UVPI4YLpILvXDZ0GDfOltmo8+91t6Tc6T8869a5KbMA3K3M7RcC2RD
1kzUdh55IJMZOMWlPaGT0EIL7HPw+jC37nV4qkNs4OwamHPM92b1dKOfu2MHMs8e
UVh00HCd9Jz/TK54ZYT36gOUHa7beuHrdFNypH1t53b8b3stgXRUPQO631V1deVd
146sXhvufNAIyTJ+1rVNKsv01NkV3INt4GE3NX7BXuf9rxiiiTxy57kCkv8kvvie
DhRnA9zcEV7UqgHpSzqPgZEPApIfHRS5nyUb+jnrIliQ6tdLQUgSZYYxsRyAOmVV
np/H9GDSBjN9ozWGjHHrx222stDIBwght+KdrYsSNZ3UP2ZpkiRITZjeKiR89EZj
Q7wsKtc10tunUvxi/Qn/HElr5eY6w/lj5axaeAeOg0Pos58U7AuNmRxgUE5tsn94
IwOc+cOMnqFThXC3KBAyodKKEbfD1InYkTpsenc1hCsCiQFQFu8ndrg4tLAhhgIb
l7YmoOLUHtAkGZWGZ+JEWBj44PwxyL60pYqF2nDWp3ZpclDAvy3k1Is/tt7wpFEp
5RrX2Mz9OjoL+3Ozza7ir+1cDDcefFbpbV8fXxE67wZPG5c4bCrnSlxLmDg0KCma
H6cUGQvVYE7Zs6pWHZbe1MTp2ffAJFmklSnsAtnt9mqRwpa31uJjWhpPEDOyM69k
OCqJtYdziVgsddY27Ck8cf/jj4GhG6+sU0bTbYGKkrSs7kT3Rk11lslospXsBRk1
z0vPUGJTb9t9XVZKqP6DRhrfHcTW1WGXgcryPjQaiko0AHN5bDDsP3LS5gGPLV/L
FoM9FhgRaW+34BRk97m+4WTCQYvKVUHvw0wbXl2EvEgIMuDqDJK2xYsj7ktfrn7i
j7mALcwGlcyFJGn382wboKe2a+aF7dWInGLpqJLfuI6r4RaJQLvbddBzK2skDaD3
HQBnGWhBqqJehil3KFx5VcXtWfF7/9xXM5QzxsAYSrm7oJGUcXWdZBuJjl49N47d
vTvctkejOJrBaODXiyxUZFv4IYSrBcOzJGPzpUJji2QHScOKVUGWpw1WDddso+oH
Haa3B//5ZcrlB/CxwSIh25BtXGqAlCZI1E/dQgR7Kgg4tc17jZLcB9SR+/sDNpXR
MFq8l041Z+GTZhj9Qh+dZMWc03H03VSkyKFTlQnfdYy2aMKL9elpoY++xvTcnQ9u
fD5IgrV4c2SzvvX5DuvgfkztZL4Xi067EuOHbIedw/ccLhxj4pgIjkoWm6sJYFuM
B6a21bUZCAD3ADUa+m0B/Sx+HrwGFspDWHcAWWXvRY1VQDlddxDSLU3LlAiW0FqQ
SXXGLlR9BW/wONR/nl0yL1/JsOPAPvwEVlX7cGaFcN/gGlQ6Ucwu/izWFSTme17V
dyUmRmWxQY+6B0tRyhjIRJB8rZVqt3mbWy8YbgWvCMXv17aX8k4UQaVr7UDQ83tq
+1P5ry5w/e08BA6vpiRhQVawshVXyF4KxMH8+/1Kv1lB6f2E1xw4PC3wFndRK6Qm
Dz7G/tG6B8Mz8LJoo7BWCEsTfFuG8tJCcIj2ZFD3jIjr1f//iMqI9L3HpWrP5MjM
eDAASemKQ+sAEjb7Z711cZbwVTCOLjvXQdqQLwy4yfRRnE9Nam6VEgWHvX2kQUUp
ykmf0jxn2si3//jfTmhUAFths0sNCe90eeJ9EGjftTBNAtLk3sO5NNZ+5xGSrRLX
WZcipqY+W5Mro5mrMbblYJhnTzDQE33j5IAtUZvhpY/zw4gcPMuCJL6s0TAf53fV
hVBK+bFmfELKN+4NBEt7Ch38WUvDMYKMVhy0u74mNQaLq7Deth9LBr3a1ud07HoH
FcRPV+lQF0M+Vkq1xUXGHxJ5lDp5H7eGigrSRWo7AETf/zIDj9aQeX4JfB4wx0+f
4NxVx2eTvmO6zCoxsjoBSKetMqAN3Wh6DFzHGkdyW5KOzt2CZ88tU0DqApp9D6c/
9lHpxHxfCFd0MVd6m69wehL0FORWUaUTlMaktyliEarML1uTGgFQI1F7+lGpZDTZ
yvlub9znID2Xp5kGhpkrSRNrn5eRT/eEEi+LR70bmqkDrudwRkWhlTjNmOM4eLME
ngS1o5tWolZcAfav1LHWDugxDc2yPtv9MPoqpRBaMoKbRQlLv+GOWpAgwmXn1um1
Hj8ClEhksv1J8Ul9UEnXFSnVNb6n8RZN0G5WnSc3qibrNftR8xe3BfP2MLtOeeqC
5TuarUnep7pzvByG7+PZnQEvHKEZjTKP+VOCyaiT8RWo4KMg9Ra/we1TkO0uqrOP
w/7muKwapZiGguQexLaNIZXWJX/Ghpn9IKNZC2zCzbdlBcBuMl9hCHtW4vkW1wHL
wVyrqvugG2m7NCnygHLMUh//Nlclj7oXmDXV5tQENj934lPI8yVn5Pm+tjnDs+ok
x11FFnVADTDByXEl/zQvPUIzsZ8bI2DF05wjc1SLr8eOfgZul8HafbzE1gjLUxj5
P2/L6GjBFmyxkcD6bdI4ei8uJDLJ98tM5BhuNX3/U/CLV7Q/S8PV86jge4j5CEwA
YcPfeS3fdElL0QUUQRKSuyeR7WlPWU2TabNylSK1t2oy1dFmBTdwNkeVEvnVGtEo
s5jdaw88e/MKk/ogfjYxZyCjXT1WVqYeI3lQKIjncfKW8QsswAQXshPaG0sKx99P
rNBeMVyi4+jiamHZZT2kl3GQfwamVROlL1ZEbHE6SXUGqV7laAwfF9KnYvnuOsTb
9S+/MfcYeb93xAQvHoplYBha4hTJoHBvLhQdcXtc13e0oXXLRiSu+amqY5W1D1zU
q9LPf06l3Ku1Ajq7MIHD5BubEVBIlJhYwJXNAGE9nN4vrX2QwhZF/UdlbvGWzG/A
3RV6RNQFZXjCjfGC9xY4c87BpTLHNFMtdj5r5W45EuOVwbKHxESBogM2kPLXSStu
4R1xe/Bm0PG23yqEV+JH19JtSrDMAfqj2xL+nJeYe3tvwWs+K6Q2n+uybcTp1Fgi
zOGzvCz7aIScHB6pISyyzelNXtMK913VBbT+TuQREBaqaHqMdZPAu/sYMOGG+k6f
xMghhTKyGZXZQO71+Tl0zBNi7fNsMW0MSN52vcYrltpMraiCLouaHzLf5Kse/BO1
3hdrVgDx8xmNrF+9emc1Q0iIbsLgK0hcMDBSIqVnRus+SrgkImEwIq0WNtg0v8lG
3tMk6L+E3YvSqb+s3QjTi0bNsZ1dYZFuYK87McUPlWC5N4x7vg35gRyjA+/n+1uR
YWJm17jc2hd4KQxvvwYzGH8DTg74XwJj6zdUiqmq1K0Gjd6AX1fO0jxBdGdYWPMs
YvnrtHMZ2GVargKDnd0eKPKn9LU70xIjg2aLuMAzN0Ny0sv2KVc1hEKH9MGWg1wE
3fZgiWdmvRLwxMlrrxbHv1gpbpcf+vcYiKKH6IFrsaO4X0gRJ+WId9W1losdazwe
IXHs3VQFg7kaPG4H3SLh6vIg03rauchVB6C7QsHQ37cUfMt0vLGc7rrv3qAmNtPP
H7DowUGuMHsVDOMZvUQBQQ1w6KzFiE2Puf8X1c4Mikh15xK5tWplOSz/kdqYpJyU
kYRRxWWEaPKrTxdIoIoYzBL74/hhAwgnjtjYM+vgPfT5/jklH/wzmJ4ujP/0ccC1
t9LsCKJTcEU7BTWkM7D5J8MPvRvUgk8IrupZYHBNF/TY9OVh2zzN3j/LdS90sjV8
NkSBGSZpqNvZTrq+5cjRlj1Fl54dh+6cMbZoSkhxh4ZcP7BqXzDqab2m60WsfCBL
75y3Qreyo8URvpkMUIsHK6Ce0URp5q89o7LwsFF+LGDBw2GaVkE4f/G77XBI9O3f
JdAELfOuWGIiLagkBOV9QQq2w5Qm/IYd6dyQWmXkymfQurr4f7LQ7ihwSMRz/l+U
7RBZFIS3MX6GM/o1CU/Xu5BwcllQyvGtbShHpIL6GvaRCWSM1508hZL7vgvsKSSM
wAwnRLbojeh5qbf973QlNZQ/Qz0TSyUHlwtYev6NnqzKWZeHcff5ZooB6g+yLLQM
qhtfZ1O796+EgRfw8jouEEAL0wWuq6ICS08FbFWlGNgnwdGcZKEFMiepi6v0V1Pj
gwD7Wlm8Rx4B3rUTBN0rU9Ex2nQ4gA76TGcdWzobh5IG/GQVeBTKebJnUdNRi9vJ
xmgKLMqRSq8HyxAHgK90svOa1xG1fnX09wtkbSm8CbegizeaRtYE+rp9CHbhVvFY
OnFJLejqLH7dvr9J0NozjwsG9BY7siC+bds6cV18AMEVcAfAgMKuUJdmvE1oHZBY
ITeDeck3eSI00UMLX0cmfwjr11RgZIp+gEv5+0lIhtenRwWi3hbXvdus9IDTMwl9
RoOcwfmEx7MSGDNwvDWfY35PqhtGIlWHV5hSFH9SSM9K6WVAwKKmmseP2QhS/J7g
ZApkZ4GRLRI/GSWYf2ift+nC5kN6yxrFfHmqiMimhWAc4H3j9h1rQhDAKXLv8ACa
ecIFUG7uYYj+/ct5oxz7CY6ZJeyB8CB1GWdF6VrbZw+VqzKqtOjH20yFfIw5ZAfe
3GB+yvdb+KM+uMz+HvESpMw3OsrLztl0mwI1rPDoRVkAjmYxRb4RDoPs+JQW04po
vcVuk9r9pGU3k2wgsaB7qZQqbBce3THfzAst9CizAOwGE3h1ah79AO8C8ZCDlm0Z
HKr5uD5PbhWbCweYkqhYl5w7a5F54HUiBAJsMDM0vxZVPbT/bGpLYr0VVVnSHYZB
HLnp46TFfrz90KP4FxMr3B4lS3AbZzrarD96EifSVs5c6KYnECy47pEcLtWelpne
/M0plWjenrNibk0s6rFBu8ZHAKqyJt5t4avef2DkPioZn66r4KKYbMCMawiU9j9i
WIKSuBbK3vujfuxEbsVYWBlx5WRFsvBseiM0JkPi7mKTqFcQJtnXcYEpRkgVv1NT
MoxeTUefWOVHeOpukD/bKTtu1Q20Z64nVfSSnToSUsKWYGq4In/tvJwV9SzpBo9G
dXBm94q4ETuxHpyGQ6SNqJvP52FEjhIjsKAKgvpx6zv/VyLZPrjarVl4a5lybELl
keqO9TZPMWoF7NeBJbIPGhg6fxGlvxeZukFV297H2P06kdA+2lvjCtPNqiqxaBCc
1YUa19hvNXukDtPkr+EgIxt5OnHwglrUT98zKJ3o/UTpm8coAA7lvacGgVugvSc/
eCjZT1NO3EspuCnZdliEaYLV1fZ/hCJQa+w/OSZymH3IkttFrbquTcN/57mEuVIN
lu41/KO0AvsYb3SSnWZH/rRWR8OuebhYmJQ0lmiIUq0V7tC3ZEr5n1Ex/9wFDgpG
k3rztTJSQogu0Hr70CVIgEiwSAAy7CYOkyrrD2C+5Yd06iuSVYoqsYtKXki8SlZg
qXzplxC49gaEDBMXxT5ktN2m5/2hd7yu7bOA/z/21w9UgKFCFGfQtDFymwF3DESP
SlTMWhuGzCEzDjZ1BE5QeYh5wKv1dq/EV9Cq80FF0XcWG/SpH69aFBpf4VNfm8IM
OwgnGVyYkOKvwjWNIKIoMx5w3hw3B6bVnYBow+yyr914HhPD45KKQYYGdXrp9mNf
Wgi9IZsPF58Y7ASg9iN2R0RWeRJ5equzSsMiskmQ8scTlCQNeGd0VJbSiYZbTU+f
Pubd9izFz8ZEE9EZOVDrCyp5CkN77UedoH6m3KtkzWQDZPSDubcxhLdyY4bcOvIW
m/ZljsyoIKRPTv7pP2omH3MZEsYblpN+vhbdcxfWlX+hcZzEvGAkMg2w3PlrQm2U
uLIMxhFCkS5JE86JVFLd5gBAyWirsh5pZWEUx4gqG4ffq7cRyhmU7qMAfcJlziu3
5IhWuyN0Nibe+5jRYLSVBjRySiOYaOX6SiwXV3q4k2pysMhQLbrGY3U1ScdAsjG6
M8NJyD2XOpz44Dr3kpxGp9xuJSGDd26hdZeIDwniLNxNo+FL5eltndojm5/ENgGS
6yUpPhnFawN4sLTc2hcK6KhdODrFO2PKSQ4YzA+59ueWheU9PT6dGlnXRJ1yF4sM
S+l/kwLd1oeDD7+Dz4SspxWUol3j/nRObgAq7mgXDrszOabw2vTULbucttESM3FA
uEiLYrLaXSoulHQFr1l6QjfHkfPWKzPpcI4hRzvRMkwuQIJv1YQ/oiT8KTay1y4t
bddpHMqwltS/O9pIwxQDAusjNPPjsR1dbamw4scmdK0G7mhVHWVocf/87T8R/Kwo
1m4sUQwrg9Fqkicj4YEckGAsvSyLNc7xES3LUtWmgeXG0axXoqmwu6ia8o2qW9Q2
9Omg96rqXxXeN9+H1hyQvhXeHMSChkG+jvlgMq25syf2rXZSQzJRbKOR1grPwXRQ
9GbNTtgxb2xV4FyklHlH/gQ0t/YosRILShF085mm/w+dTBmt38ttLMlLGcCxWWMt
auQVO9njcF4ERMrDolvuENmQu2pyG2EUlqxY6+ZlOyYKXIz0vk+0R5HyGlkZ7MOj
ERY64hCqtswU11X87SpIuEJrmJ3V6RYZ5aGiPS9wyzSnrBkH4kG3r85pcbYdSJsE
b+Qat/2Mx9/vvLJDiaqsKMhTwmRUGtTANxWbdlFc6kGnHQv33UBKtEdKxHydGfte
CTWidkxd1ioqQEYk7j2/ymlRPhYTlwDSkIA1G9FnwTDg/YQPebBWEMvJwqFWfY5a
2IXbr72eok5kFXcfmtwa7AuSlSaIRaZuYid99Dypp+Pgcn+ipXy6lDbJr5Lp4ShV
hlVMlGgYkKji6PByJ75uolUWtYWYkL1V2Njn15x47LMb2Li3CNZtjlP8vGA0f5WS
eSmxNkAe9frCZ1H62coW3cYOqIwvhz25mQ9oVYrbQea0yoOuKjmc258jAKpa/U6e
1YGqMDyDEYLJDCmHsb3t11vrY6Ii0o3HItf8qGzOXq3kNgDbOY4d+CYBN++cyhES
vh09LgvyLZI5AxC43yfLMA+C939rOSBZeIrvpROTa5i8ssUZvUdX+4eR8qx0VCeN
yFJ6eEwKSNXeqAMSyJKUZ4KngU4BzdaVyv1CmxjLLC9H7wUyUDwCQlK8NwGTRaMr
b+JC/penR7YwKe24+kB15WC13YYnt31PNJBOv3Qt6lRCUtJ90a20MVY3Pe866vAB
t7Obz+6PyxiCw4eN6jD5O6bYiNbKgsu8543BKdGXhFrtTCJTLb9D8nyQnlftH4GT
8mfJntgqTPKhqRgTVde+CwLBxtvNOgYoQps4SYS4++6IlNGkMEqBwM0vq79IDhIX
1mGEPTEn6pb5OB8HIXAYrjgQl6CA+LNLAxGFI8utAkCh0X+M9fW+Y5rVATzHnJOf
oo6FHmeNMDI36dRsP4dev5PsgpZ+Saqmuw6vgV0OTv9ofN63rPZVIGwnP8Uk8ub+
6dv9UhWP2UNAXLZLJhEpUbZB0GGis364psNn9NfcEi4Dskz60rdmgrM5t0s4AitL
mh9Aych3XymUdiwyRoNQXasdQBs8Ll38tr0bBun3pjhh7cW6I4hkIudG17l6k02K
M87d9cq9/D5L+b46CXaLfrFrTTg2Zzc2Jmrb9Ql25eChsX3y4+Sx9f7IkVvlLOSZ
pdMOxHHUc08YUwMoaCId5x19+jqPirQOalVQ8ywRCVAnGNit/x3qbElR6mKeZQ6N
0CID01HyK9Um+e7sg62YuuTrCEAnNaj+9GksNgNnN33iivoijgwyTpiG7JVHstj9
CUjADxc5cz/QIVr6nXtB/56lzbOL7otbOGkZAViIZYlGzMheB5eBSp6xOZzS/31n
pvH0vtuzw5uwLlpFERZcpma9hdXc8mC1m2vNndErDPGgoOQqB8Mzoptk3al15Shq
+0Y9z53F2cEDr5yqEQIaTXwhFz5bMYdJBK6Axj9zvpT4nrGyCq4mPQfchNLXROHZ
kLUuVv4APw8KmOF6UcXbLAzNJux9rD2tgiU2pwqYfOmCACzkjpD7Prt+pcIJCYmH
H3oqJZuLwPev9qCbAoohGDRlEYmJxrP5gRVgzLVHnqP1Be6jiM+k5xngfCzoA/XX
jbLCZEtC2GPNiv5ZPxdE6Iae4NhhyXONZlR5Tt2YtacPboiCgV93KwnBRltebFxF
Itc6g113BoGczQPTM0qayPce8DDU4Az1v0ErVpUjgwchpfQYOgHIUzwRS4lMusUr
zQgViFA9sdqUnPj6+i7WJV7mtvGLWD6NIOM1+xYySNfkQhT2NiD9Ydc8yWs1ZBvT
SA0nJhpEEd1Br9A+kEnHMh7jHIh/ORdBc4AruCc0316PJYxhWM/wsnJMJ6UmmsYd
IIhX/+/UyhvTWkcH6XIeT2NCxMytWkPSSDrlhMc9MVMUG6X/swmBWG+53vo9h8LH
5uMh7o+FhlkG1zGNJBsKB8sdfqq5qfFa3CleLyrZZQa7GM2/CGUadvycon1NMjBq
ESZni5UJYHuRh7R1f39VqNEvGcsadD5rG2tv5zWdWs8AQlOY+/rVI1xLY1vJgHl2
SY+kFt+2qrD4nzvfQOupMvBgh7s2wxd2ED5Lao/cJcJT9mTe1E7qTgQ1RtuhVpyU
PoMqCpQVP/fs+zT1mKJjxr7o3JA1JLkfVPcwt1mqHLdM7t3Eh9rSzQchVDPKUP7d
/n6kmu6JcmuapgsGHR0zfLDd1gwfysTPGnyDqPUgjeagpEyR+b1RWtibzDKmCjqQ
eFpBn31Pwq7J0cf4zoLu5m61D5Bv3lsLk8aumLH2Jy4CjUIGkZAI6uv+i3oQe11n
zICE0JHShQQvGA2VecLTqqAiihYEfrsZUAvAhUtbm++Van6KVO9BbotTpPYTMB1K
247BcoVrOR+OQDuV5Nlb/sQb17T/FcO9b6YrLfXcURcCm9WEaFkpPhe+cJkXxWW/
0PR8GY+0IUi7BwKaCoOTkIBJoAP4WPVDXz0GR172EpkOulyRYno8JUCW5uUUHpkg
qvlgzWKvxuIFDsAE5us7aFtQoattnwDKlTF0o8XRewUhf3fv8IA1QIYzHCGnv+cB
f2kBES9UcQ1wSsUFpxaZT0UBXExU+WG487BcIbfzf7s5ZcNsOkUlzQXT0YFij16K
PfnqpTskovL8jKXDBCaaGMfHBaCf78+8BGZoXKBhad3XxtsL3mgE52IaCpY7vfyK
bCE3ikguybBE9YoVWPgYK3QFLbmq2PxhPpVACdpU1HGb3DDaqFAb8fbhhjfsEQnQ
VlvGxL8bdq/VPMq9lTFu8lTl6WfDUx8tG33OMLSJBHrRMKAyV6P0USXGjTjKDekT
t8Tu7Q0i/8goGu7W5IteotcywZvll62cTIvT6Kv7HowIM9eTRWlP+L8SS8MoxERO
fP7GAjXAP/QBbBP7ZwkooDk53vm0iw6qs7juUnkQUbf3pofijRWvKJ5yln0SGbID
mvLCrlUaiEr9LiGu0IP6LIMPs94wbU27XZc2d3zmEFlXNcPgCh0mLh8Wy/Eadoy6
VYoKj4o9JOKyu1PmKPEergLhYbc0hmBp9qiDu/xrILk+poE1UsawHB3zPlCpAemI
8vO2dunohxz1waizYjcYmUwEREwktyrz6KdvWc1RmYd3a8QLzRFkPqbHC/cE2Jfl
0loQGPZammDNGzpxlXMIl97SRYN9PLhryAzX7FMWSRdJ0earsTNAABPt4M8RizNU
0ltro7eXdjJWiGEUiqwaplrzLoHFnxnZneKJLSvo7ashcnyxydr1TyZegVGzTYgU
Bk5h9Ankgm1dvB6XvzjB9lVjh6zRGbDwFukTxwOGfJejGLc2HWY4SW30lhKtW1zR
I4jJ6GDFB3m6hNC0iGd3udflrULtobiNcwGb1bkGKApqUiAbqNNNS2h3ssJtnNNT
2+xao30wO7MjGZxytlVdnCH5M9pxkbhHYZ4V/AdGZitF91kyjjzyGJwdcOHv6MbJ
pHLtAMcwyDteomiFZ2QBTRsYQgGoqoadCUtfZmpuA0KKl/kvvzUhfNZv8pRoQziX
k10mnJg6+a8PMJpQ/qdlticiX6FqqakNFaRQ+5f6g97WHvUhAcghSOGFI5zyauov
v11IXuqPDoM149oJreF0qrazRo0mefYc2KCqptjcWc8TPEvBS6wZOzwUFPQJVzsS
ym7tWdbAEj/5zdbsj6oaUQmg4aZL27cLtBj+2LDkKbZ+aDO1+gLSMdVMZV4HREAd
fMAx5d7szsbToyPq7ZdLjM4Tt7mZX6gLmq41ZDhmGhSl9+24KR2NYvWl+l1oxjus
mmTo34VLrVcy5scDlv16a42CYyGKEdaxTAUJk8lUUSCmRmZJskjYKXRl6CERHTNI
tZ/FfhotJBU0vfu0Nz+jFshxEYGduXSxonRgoFP+jcz8XCdJz/vldW8+ugMquNRP
31LNfKij9YyzrN3XuS/ooKUServb8iMCand8BQ0bjy9qscC8jsRt39YlWkh2MI+r
Cdv0mfHjpwzfIq7LMPgSiQJJSbTb3YguXUVwL66z7WwIbeCQm4SuPbU702jF710c
/sZUUIuDZyk98bYHPNc4taNGDKdUQt56PgfU1Papu9s2wxk9P+WzO+BBvfC21KEg
zyuThmIr2OCkzA2rh8BZfAZVgB2isu3a4IiS3myBk1p0uDuD5yOOOX/e2vaEcsFk
bClF8XIr4QVzSWvBdu6CMlM9JvKDt56ViGz5zXXUtuZWQqSeXzrLOQoaJeEgm1Yw
gXhOowEcKO2FHa6cnK+lYCiGu0aTdmPq0L0T7n2pLTUfrmNqP4SB/b0I9N9Omat2
Z2S1+30Aq0iOyN+NO7joq81I5gWp96OvbDrmY8yzOooEbuU8ioHGx2MFHEGIOKoH
RJ0QaWXqJ9oP+fn3WJML9Ybft/LEa2wz2rAIKlPEkonD9pgwAAxXhPxCw5jzDe7Q
VXl9pDhrL/H8RwHgBKc/wB7Dk6Sup/6saUq3mzdpSvfC+9Wi+XdnVUczPAn5UvDw
zfbD5XgtQ6QZiR7MgKfroxqKTxvJXyeuF1EZyzZteL7mxpis/TAOJpCammPosskd
kd47TFl5QCejP2fppb4aV8n3JJdxUV+8KbH0x/Yng0wSr2rTqkxiaIs1PqLYMQEl
e0XbTZXbYgjjXW1xbS0/SAMhEykpstkIDeFNDHF5SwR4xXc/F802qtnRDsVfvKB6
uoKXszEFygJIgewFSw2pUQpAEpCYTUB/kq2AhRV5vlw49iksuQ6rw8VMunl5eP6E
gXnxkO3ldgmmXAFd9Wogx7atzGTOtDMuh+7jNIuPFogpSoSTNqCcbGF3RiYoSwxK
OSCqPFn74Hf5w6QFSC+b6MiD47/MONM+zdQ4j7aXxwrFCff+HluWZH5moy7SjuC6
GYhtUKdZpVn+c+X88gSKnqxFe1o1W9CrOGIgChnzlf0A9kzMUwNuvAwAlDLOooDH
0YxCQ8DZEZFBGBo8yLQ6vzRQ6dHqf+ZDuEwQv6aZf9xnSnmZH79lmUBh+miIdkCx
rxY8y17ayTZzqiobeV4OnUmMqIWJWgi1q3/I1A0qFujUT8UeGe3Xo5nFwH1IxjO4
CJGM11fm88s7rROKgzH/fjrdD+dWSn8AtXHxr4ueaAqsVtcqEinvbwMWw96649zb
m/TEJl+miXvq3FGlcFtEreQgDFrEIoyj55cki0/Z4EWmtxuCzgPJpyJ0EYoWihy9
xNEHoBx1pjW7wS1PQja4wRCZLDcIZ6GMCD2QpnZuwIU0ASxuBpm4zvQWjPV3Vi4V
vyVm/knMqyOOCw6lo3UHY7JGtuYobmAaOqrYYolV340traRevZFW2W2nrU4/QCMo
BKPE/J0KASlY3O6znDkrhXPyhgaS4I/E2CAyjoFHZLYtuNoCxAoNYmZNLQWtGT+4
63Hc3WckUYVnKMa9QtIO+wo0gH18fFqyAugsoXn1vJzsmdasiyUqeATCTRWemI73
uSVgshOXtz61HiVyKO0w8xER70f+JSfrPWQe8boCqH9TpEa9cX5RITXCvEDYSEJq
cCJxilu3YZyxEz8aMBUBXOYvabHg5KZX15g0nK+gur2BUzDLY5gk+w7Vqz1RxozW
V6wcHg9FqYlN/+v02mzgWU+p9Nr9YZrLKJBBtWAxbGfeyWn+gjxwmkyHPHXQ7Wvq
/ua8uwiMWR9n6rFgJoWKXFEf5bbmaeByS3lw0gMsryD/hAjgQD0h8YrXqfVKhm8u
6Vc0ge+7biE9/3b5urIx+69kBB7eWzyJTFA990996TqIty4/viQ9ZFxNxXV6M7k/
W+brWqAZM9AqdOe3UuI/h+MQl8/vczBTNXm/y2f/CIABI2MxDvixhq3oNJo6mwJ5
sYYP63tNUBFkwjM/8TC4AQanRumrlG6jUlFevoHTh7WGQDeQwQG/VApitqzRM4p0
stvIosPhtPFeSIxsMORFTwcHrWf8HLn3u8wT6XPwGmCUF+FlFvlIjW4vgz3b192p
8sGP17zhiJAijHhIweLXoM2aeMa2bF2LMsJSNO8joJRcpBcdRmoMvq0D/YpLKmko
m6aPR//hDFeyZftt1U42poH1kwn0yy2lOj7Qf+GWlkPbzJ9Sr1/GWEAdWgeY5js3
K3yu+lrykpYCML3LxjJdnP354yyqWUP8JojviXxYSM1mTg8mqS/MLaJ0eM8LbDFj
1t0jcPLSR4D+YSJTE1cawvrQqIToOlr7gZG1xUjXkv6oZkETuKiacuWy0a3eFCpc
bDc4LAxhhJ8lzatEd1cV0psRHdrp5evBXOKylqKomadFA5TafaS8WGEcUZSFC+gg
Qyb6wbWoMO6JfDgvzJ8wJa8aYZmGtFhkb1G2kLtwX3jXu7E9vrOWy/SD23f9J6at
99u/K7PKJrmMpbhMn3vyQL/U2Sx09OdnHH0g5xUKD2dQAGR6UMNR2OOCT686qjm+
C0c3bL5uJ9KrVDpyNgDONkAXH7vq/nt11WMt5PWXdSYntcWWYTmwhLPVCWDMw/Kn
9OSaGrFSwwAHuJeEIWpTxMO7/nBgkllip5jUGWR/fb0FFOfjrTEdFwq09K7sZl4c
n6n+7XwsnQfgayt3qp6jilgNG4xORgdMfFm7R23mC/57EeqcfFF0IzcR7MZGvyfv
ER3fDOeS+Ofj3r8UKqDhsS6Ymd0JSnihCy/GGGOPwW7CyfaerhmXN03YMjrvqeTR
SMHJPLMS9WgLXUT/y0PccPECyzXXZCZfxgrMVXccUHTmPLEe24mAhRn9mxUjZzUF
DWkt3wz2BaNuxT3hpNDl71O37xvqHOMSZXQ8CJPt7RIJH17p5R4jEa0Px8rj77UA
Pf8NW1UfLVcPKrmS2KRgccrkPBeTghvMpNCBwo04DkBfAq3w6m1nDM7MkDErpEBv
zJUNNro5/ouy1TqA+qPfO7cMSX0yVtrmZtlLFum1Tj1w4nA+y1/wpJzMOXfs7/SH
/OOAzquAAaGkItDGRU31kt6zCnfEYtZmlK9qDv0TrCepvVVryzFVowpvnUK2UclM
IRNYnrLZ5CH3szztGMpXu8iq9yPvcBSTnZ3jmrAW+H/qTvwoEwqu6lXfmjAjnOQs
ewWRkwe3/1CfGQSXElR8p8U2stpj+bOChfoTIqhPMyfYAjtqFvjvszWofkQNizpB
WH/AXE5p0ysK4FLTHfxV+iPPFFLJuBC2f+p7UIhNqhjnZjzY325Ue9O7F50ulY6/
PZmgaljzj6OJsEy20zA/0QzpCIsoCww1l+ZIq3hS3ub2KGJuv6XavxwZSGIhTd1l
DupMKR+jgKCUeMwxhXDmp3UCYw0s60lqqU5DfmDwNlqYTSYJWxythURWXlrVcdqA
PPG+w82nWTxIuoUsCz4Hk1EhAGWxka1g+agFlQWPI3+r0PCOBPivsu4ECW4BLB34
zmzGhrpdSP8nm3myjMx523Kc5cgCrxBeiwNge/tgS6Eq+zYr/TtkLgKBvbSn11z2
t7KYW385UKQ3OfpoVe1QyzaxBZd8ZYKkW4mCGJxkn4FEwWxwJZusdGPqALjAZvik
/HVoyYsVZQu1jtMfMQe1+6MWRQxW1WpriS2R8uSY3Pg/Fxkxhb+nOH4ozsHfgbg9
ALIDFkguXunsjmONTs8V4Je5xf8ojxVuZi4n80L93AdUUQEb0k/csxQumxgsJKYe
4UVFEDvZ6bzBE4jb1ZqDqUaQN/vQ7Hlh4FyPB9gRAD11+I7XWETb4rIlSSTs9Ilr
m4qUwxcDWMv5PRvWWcnFAwPxWHszEx+bwRKc+5IQa1Suy1T4h4MS6GFxChMjlXw2
9/tHWApiv2GpkmfmDW3w/wRu7LeYmz5dXGa3xhWHWvhdMvJkiKefEFDxxVPUkqkR
VYzPC2gYwqLgrq6Lz3hlStdkJXQ/fKqRT6UWO/ItDb278OwonkfkKFuCl9Z8Wt61
+ayWNK6AgrTAOqNh7Aay+1LwE71XGSdONHu8fUhg/zykJ+ilYh0kU/ZtySeenAdk
6t/ss8X0bN57mNT6CCbqfOcwJcKfHdK9BXrwb1oz+LQWxtV9ZOmJOQyDsB6PwZYN
UFDWik3uS/nXYmepPgE/Swr9UrSa93TR76Tkce2CneEiqO4mKdbNHIOck+AUH/Jb
l1TQ8jEIlFniB3BCNRo++pJ4TNKt/Xo5PdOFXtNZofkAIizZZhm53UDG5K7y8YCr
jYTBJ1z5kYHqwqdmm2Ib8spzxiN3+91Jv5qqn9qjqr8cMsk+m+oPtSs+7YrA+akX
mon1e+g4ijv4aoImaW0fHj2htCH+P3/baYfvGiGjErtNY1YXV9GmVDzhReHX9xra
Gbba0XFP0FJV2XULdjr5mYdSkwORq72sU4o1EG+LY+zmzrKjckexEpzb5qRVQgmc
FD+jQnz8qHhhieE+7VrY0bEjFgs7vE6ObTEtGG5mWAXbo3DnDWOZThxTUQ8MsqpK
tbQt9MmIDkHlMtOtrIkFskW7ieffsyVk/RlEBrfR5E4GlPE3+myLSAfGi6fHZzWr
mPyivNiwQI6MsZZk4BZ0tsQwdNBtAhSBgwa2TBg4Pioq478vL2rf5/v7J8rEzWvt
ysrlgjtzHfNEgABVmcUHpKtjdUlz+JGMPwoyRvCJyu584ty7OtpO3Rf3PnXq6wc+
k+WcOUlrw6z0sWNZxXDd84Zi/UVtEHRGgOhAyhIX158c3uc3x9nkxmdZFTuB8Mlo
Bi+rmedNi80+BndTQtMqNziztljlHTt5BwJNFEptnb/S79aPMyAm6Slo8fdIw0+w
TpvkMILptaNBAxNDZKHQfXaocG2p6KkiCgznRJolDvVb3H5ezwmYhukJ/Kea/hH/
5fcEaqpLU7LmbvxFUIxW0BSmx09cpL8XUmwg+CJEqlThb0GeLPXoGEk+flJi25cK
Wpfo8uaj1nsC14aXhcMF4hA56xF7cIizlSWCjOgpw7b/i4uKEB14JszR2RM7/4Aa
mdXcabym6BM/Dm37y887uYQQqOESko4hXilhvhm5+rJVojCvTQGrW8VlVFs9mZ6X
khhWjCON+yWEQw344GRvAPNH7AhC4g3oO5mLyiabZjUDRggPXZVYNh8BS2m5FR3p
CqFomut5fqTU5raw37uH25fkLLPPvLX4htWjQ1SPFDAp8V4zDbL8CHQK0SzjDVr/
n83p/3l6BeTKNt3dIHVBqSaqhHeCLL3zHE+JJTN4iX7NS3ZAql7jizuSTOK2ejZt
9joijyTuXNzrqoO2beZNIXDzsZ589k6g+p9+enp4JPKM8Bgdb8/TO8mu+Shy+AnX
U/rV9CEcHs3xcwA7G5uJ8pNEXjLJuyM311KZ7PSOo0Ys3a+KvlwjVoLu3g5ucY8r
54IXMIOzP/VdNCNu2QbcsewAfO4fcn9oWPTEpXI5S3l4FKMJ5RiezoRiIo0ii6TM
3gMzR0vJirnZ3GsnOkMEt/ibPozpg8ZvZSzD1l9rZb9HA5WVCj9xIUtzagxAMaC6
Su8grpuN/gSEBFGJikVR2c1oOuMTzABD+eUNsWD93PWiZ4PakrVkxJIzdi1pjfRG
yHqC+YqgQKx0l0MYxtO+jC/oCO+dr70JKec8K9J9y+09cQZqLFUJcsaQV4UoCQeC
PKPEKCFoNhbhLOn5zLre4ahzYvmxYV9k6BUCvSEHNlibcS7JSwzTvwpqqKN/L3h+
Mt9q/NIL+JBfb2BZ0koYdz+F1+yz2WX5YipivFLvZXNm1moyXgSRBmoN9Am6+376
95wzhQyd2YRf44lEra23OLg3Afm/SJ74ZEaT6Tb3SRW1joR2vhu7YISogJ5/E+PC
nvIEMb5htIas/JHT30WkJT4NoJM34uHQe2p+jw8PSantFBDFXU5xBRoBRLu46zxq
HY/QI/ooYNWu6n+Hd/5XppfovRhr8zBwvhE7SmKaqqF++5U9JUyH7roAWk7IEgha
80q50enS1rOTtgvmGLDeD7MjY/kvmXtGesr+jqGgR3OfawJpTDW05uIB+NZLiW0e
xiDGX5+g2oVcnFdjguBwbmMmjs53H3eK41Ww+JxUlMO/4QazprHX6wfpCE2BjWfV
3d6pdi/94BSmNlYSB/PitGcL3TVFy8w/i6BQ26GMOAuZ9lHmcDabVYrsy/BPiXxv
toXCgiRE4YzRYdVf5fcumkKiA7FCWETN8PnhVGnFXatrgMsKTqojNW4lyAYwkl/k
MSn9GpPfX38cQWA5V21k7VIdQrvWjAP2aSPZ4aTgKH2OZNico41ehJCl/GoTylfn
5duLaDZeWGJ+EQz+4liLsuURm5WZ7ywliIE/wcL3c6tKYD0sP5NHEItqS2momXwG
5BkHH+3u/Q/Zd4XlLkMfjMpRgWJhyZXHk8eFM7KcydQwcfdfmRqiMh2gmuK+FQtg
yxgRXR6O2AHT4pvXbuM9ZdwaS7Pdnf6MF5nSklY/Krg1kkAIrtkdSSBakSH0mGqx
eTjErAS9RhpusF8ML42UoNB3fznFb9jNyL66gVfu3O1H2hd4nhzZuz78uLPoco/U
LSED/FSMdPm4FSDhls+3UnD0xWKG6WPT0P9186KixtonbDdQFqOxEjcDWCvaL4BI
5XAgYWeCsZypVzwkham26N+sRoJj5/vD9frn5CLjfs6X4kTPpIOUx4HW/vtmwr/7
prBfoz7A0o2poVHTaC1vfeXai8Nj+dYOBBL0H4wcTX+n8PvkaljiVNaTpledrMI5
Zr8nGNJKNptRb+H1t1wBkSuuAiAvDys6+I8yl6i5QpW43ioVpOcd1OK/OftHJdN7
706PaQ648OkErerje8i9MnbHb7Kv3EnuLw+W77/fiOhRxh8zwqcoVaQEXZT+6VVu
zg7NCcL//H2DEFSHU3KklSUy/Qk6vVphApVzcuJmElNkgjZ/jF4bYc/XnL6CGTZt
9jQAWiLhtae5XqqnlsWrNWgavcUOQzCbbbLDJCXItoEY/yQ7LrzrKSOEfH+hQYSn
Eg+HMerre7WMugNZXygr+SZSI5w3PvoqYqemH9CkoZ4P5fk+b6PsHULVU6CGncEx
N6IGZ8fa+D/1kuE2/KtPkZWAMhZgzL/b9IEH15z0YbjzX2ICwLzMhcZ5A7VDtTNA
WmJaiCqe2r39f/FCSpVF8IJb3FDqEWmvUVntPUlG+ecs3bQMAmZscXHJbr9WJ8GM
P6+UExrQmWyNtOn7OWhhMVx+DTgMn2pSZ1wblQBpQYfh/7GdoFZLnKgojzJ1pzPD
NbgnEIjU0ZJHR7UfdLEOzr5FUtfTUp6n0hxukLMhIkHc8hMEPDk6Wm8xFAZLVLEB
x9RRzVdfmqKx7dYk8QL97GfJl/nsmLldv+3VrWv+NpT2mRWRCnMTDblJzwOvo+Ou
in+ZfoaZeO4VTGDbAzYZknRIfcwpFGJpwp+9608sPgNMLZY12AtwTnHHzuJcPSTR
1wbGz/OEtxdM76XA7jgwdIu3nYHuBsuqzp1dLCFJt+2oD+mk/EdwbrXq1euShTgE
s/pheqj9zozAdVT3uS6PqLtaVQmxtjipTMAO8UDlzJTpxNGVC2ZY/p+Bsw1MdaTO
SeH13oA7FESq8rndkbBTC1/KQrLdeyN8JrIJ2IQMth/+aCrj0f0yz/hV6JZRMtEX
cQ/OC60IIQzlHPX4wKQtEmZDwoqWxANh9/4rcdLUmpRKhl35rVINLBh2o9okjfYA
yMTAqxJ6VcxYaNwbBirfcOySrzvfE8zMFcT1TuyBOrWyersO8lLm4EOE1Z9pSH/t
ALE9KbKhfZza66XJ7lgL4KkRhCdLpLxBCcbHwqCwBBhc4IpstEsZbngwzPKjLoPs
dzZOUpT/KGeiuh6ENqXpk/nfqo1jpaWSWg+iSDjfoHlJnuNoaY0sSI4dY/9auJGl
Fu2RCEC8wkl1z5KIL+O3dd5RKTMuCa2DnHDGjwrtT0pGXHMJ0JGvsVIMTPLAncn5
ho+4lMnQ7ysKlUGZtpJPD9OEahYUFLcRzie2fKEAJnW5rdHJPOE6/X4J3fkzjgKg
OPS8rw5oV27bRL6wotkfqBo76ENa7zNfvd0ndEp5EKvnrpIjWSURxPXHLp2XYFhb
ONPudqnxK5TRQrrRDV0uwJyhE9V5P/3hH3ZkRpb+MwSE2WpmD+ByFWk52AbatZ2r
bpmxH18gqyBVYzVY+FHF7RtnQTwfoENGiu/MIM4SIYhhmvzqtSlEfKVwTNuW+FcR
jX1DLBRZJ3eepJo/OFJrgc9T7fHUs60IW5Ykpt0kiF/oBCClGsIUsG32VOlHD1Uu
impzOM9b701VD5703XZwj08vat/GuQfAfQixO+Td0CYNWZXkMRRGT9jusg/sfVeY
nlQ8bzylCuL5HbskGDCZUSgMGKrRNbgCk81qYpU/Mi4jzrAo/aOYPSKbDwRBj/8+
oU/bR5fvOG80Pm3NZ4vQ4Csnh0UqrhvFnC52fkiJwlgL7zsDofPs2ZwOGe+gXROG
lowlgB9K2KhGcOnrt3RMjU/YpffHap8sOnF5SzLDrou9eTDpbAd/y8JZ/CXQe3t7
Z5+yuOC8tJt7pz23ZPuHaXnnkDnWoBEwmmjF7LO8YyjZMA/F4jX6RRxtAeFp1epU
0yQ/mdWdpWtqFbd2ZRUGa7NpmeaKx1D87N0k29Fxf9Wrajqgz+v0ajoDRcXmNX08
GRemlWJAVNHCR2af17j42vL5bykTbkp/TYpb+mBPP4978w/Qey4LVZtehPoWyYNK
G5JlQsRV0tf2rJ4WUYfMYk1nJCb5k0TetGn5IjdRGq0bjqOLguOts3nJDWm6mbXx
Tv6pChuHoYZAdrMFVNOc6sftg6rCTJWGu4kHWvCdGD6y9W5Ls9mvnDapRGYQGUyD
4quTkskFLpnA79RYkcL+3/r/ph1YGnTnMrJMMTX74JtRw9LsGPV8wql1qA8VjFuw
M9ZHiUPjRYTVYvM0Cp2b1/V2vS754bBB1/owsin9Yb8HQbeX5oEJmO0KoQn892OD
HEgGFfcf83Re8ZnftgQlRpz/eTQYkppiUhv81QouWn8kIVPHdMO5wp4kchgau6xd
4+beMVg5a+brd10jiDo4lP3nHjUuHXaEd0/99xbpay4NP/hQm4D5KwfizAgZY5nr
mThs0cy/PrSSzobyWJvPJya0t8N8tWYZG9cfW7tTVxpKiSdnI/cCxJBoEDi0pE3/
wpzHsZjKYZIQkbsRztWWty9VTBExaR+PXL41gtKBw9wccH1wYLbrIQpBIFOh3/la
JdH/HPj/1IGcD2gjBbt+oUE7M3U/pC2d5y7e5cDdmK13w7Zk4UQMo0hoOiFdrK6O
j57mbUP2vJyNdwLdOitIORA4bDpASa+mjXubxU+0fTnwYZWwWIghKUXQyjGwaZKy
W+C7nBm9thEBOvCRDAU5sKM7PO8kRse2OklqiR1S5Ud1caQC6z5yrvbldHaoNhY8
mPXGuc2xqfSnArg1eQnmwzHOaOFil2zQAGLQrW/MXqoid8qHzH1fLj0r82fLukVu
SUj0wu4Pgm8yGPbfJOJ9UIjEeioRBn6wkrdcTPSKF0KHoOZ0QX9iCEsk7/WeSL+w
Hs6ioHRlraRwbSGU2Ck42N7S7gKf5YC64Kih2pMr/T4zyZw/qUCFZcxPc5N6zfwv
Kye51RT6wpLtEhzdUSh4p+RmkWeacB5dILn97GhDn+m/ulZiSfcxneIUFqbowTa7
JjxX3rL/crV/vGIkNS05WUg41v8oFACOsuDd6sGbceNr3GoIPwtAnvVYrdczDGsO
O+Wa/B72UVArWZha5Od+vKRlzReCuZpiETqyBXL3sXH+O745eoZ9zyr9xA8lMaOp
yJ2yTU4I5B8QT1zem8q9At38A8EsjzSttIk5VNozLYY7P1n+n8lBeQvS3Aq7X7PC
VGWSYPmg8MAoVjF89yN+91iOzMSiAgmJ6UtF04wkAmwnrd8jgVN9RUFMvEVcryUS
b+IUzYr5MCavm9uK211ozFlkBbsEq58GvTPBr074Sc8a/6LyrTsN3Dhhu32OCXdB
nJndmbGtEI/coIFSETcr1GbjgoPxBtfidFE9zV5+DTjhTkIXnDU++nC/kg5XDn10
Y9QTKLw0Y3JVWke37AdLJOTcvtWppfXtkZ1yfZKMwNeo3UzdO5yKm1z6midc30TX
Rf1Qri+Aw5T4BTuDNnFZ3WqH/MBmdKu2YvhX5jZnjONzCZ35pEoKknN7EbHidmY7
sHaveBUB++5r6oFirRdUHmrlitpo9hv7c2ANzBsSaGjBfTWsi1ByqFRHm85TyCw+
YHaSIsZQHcxxf2lyoeOlPuByiIGAKUDxV4vXUXppVNuJNG8jLof47vKkt+N4Nx8g
RVaYFBfnTYzYNbItCdjhQsg8XcFc7C/ggqTR7FuCewwI5Un1qDRngotXOn/AiURw
PX4mSJXpZ0nG1VU93iaiBXKUxqguHPCvh0nWyJAOzrh1PhJwk0a9inWLxH0MAxHB
vx+HnYBy2Wku+3hNJfTPSLBArWbx9Ri8a3o3dufeji3JelSajx3jsOhvEtpstIx/
iRt+B2GYDLQf227E+MyP8TQL7jiK8eK+XbcWL5Wx1TKdbsKy7lzC486Gk+enFJel
mSw3k41k6VHicF7SAufjdMe3ubqAeuGbQJDkmQMKp4evVkrh2qHIB5j3AcdqwN1I
ZazWSlmTigZNUovKVUpZZHNFoUqbiEaZjwna95O+lfbSqeqJw4JFZTv5QAeY1DzA
4y9lqHqL1H/XANdXgZNMMB4UfFqhAR+3ExOnPeBhl7Dw0iOuE4kfIm/O8N/5O07C
RL8rM1q8nmAugAm7FRel9q+ycMXd0hrD06PRAF62SmH15ZtysyuKb3IhEXFhvJu8
5My3N9axxDANnsdAy7L+PwrnPFpBxPb51D+dR7tpMPC2RicoFsK0cBsaOX5e/A/O
JXqYkNOzMUbQkvEOUvZh3IeugCNb3LYlp7j5kZkv3NDgEzyTGvI22RJCtLOef8lq
QTUdgkaBZveUHmjdvDBCNgMt6zWdR5KHMkZ5gbcWds4OAKzOI+plDANbwiIixdgC
FU6Ea+yk04+2hxNFOSnNA8F4W5QVeUTtFVAGxLotUlvn6nbUk9E8kSxhjwfY78OJ
3VirOOW3UPMp1DrvefVZ6YeEtMXdJ5q63ZEwrtmq5zGcJv2eDnYJjth291ogq0uy
XY6Tw5hQ7n01kq2ymMaX11wjQ1xhlv2zcPIbOw3fKW96LFRm/7q/JyNQv16u05+W
WaAIpq4PLHZsSUQDrysH1gMjH1Afvek7B7UtVxTFSEooOBSadFzeXufCT+tOSe0D
37+wnILeRpiD3mfu6/SOhTvztltVFyendss0Cj3dpW3VLTIKsnnYpzMKVslVCR6e
8Jyr+vqO5u6gc5I1rOU3+I7obqiHA+kQqLoLlCaPxX1xrq1mBQwoGCW7NxDJCSq+
Uah1S/CdDd+YckNSVrSh+5FwGziu9UzAG4ZSCcjyrLORq49NzscdShHnGRPMqk8z
lka/3CfLV2mIoIcgLNZd/6igs2cF7Eh2edF6KNEM2ACbBxU0zd8syimuy1PJvUfh
7nLGCl3aitHOqb2N+1TjrV42I68qsCPnHbtBTOgEkd68P0FeOswN+O8jBlne1d6j
nU7rErq+vzHYURRS0nYZ1lKh/IU2u7njb3WNTw58VfHu2OlKNk8Q03+cCNSijl3l
sXoNTiy+Cx6O4pfXU73+a/r6sE3VXiWX94ARutnBVMfe751UZmiAPvo6dlbN3rsx
L3/EqvTDtOU6F0wvjLfiQ5Xoxk2jh48ULWxUtWZt1LRHciE2EIc/sFNUtQKREUWO
Hvj1li7yksgiQ2UdX97BOwV9Re0YplDUMF3X8pOm7tsbt1jlSuwkc6srGNCYsrRs
yxf9R0cSV4mysUEU6jNEwB5Iex79X4lpRuWhLCohdvEIpwrgoDydpGinP0A8p7PC
W+Nf3Mk+L0NWNQt0g2hnl5psg77tzKrvyHM6HbxNoLr9LPrHQDYlJLeztI418gQm
Zkf58/HWdXgxFjGtyqakCamI/v7ie/D0QP4xjPRjlFNkizHhNgTB9gDOwK9ry47y
gNWqWr1Q1bQRt76X9PHZwU0cS3uJq6qVP01E6faIXlqoWYBekf/a4f0mIMtOfZ7Z
ZHAGiNFhvM+o+iGFaqznj4iRKbpoRyuafgSXpU3zMNWlNl0g9YvAHdck9NcDx2jH
acyzdWgcvrofMKMeSYi0+SfoEqqjmM9kVT6MlF/hCmHLRes+WlY7ntSBU3A5XxGB
isn6wZf+AeG9Gqc3WOUmzystxBZtDYb6hMBSOxe3cvVB73c5Dcv0kEB5MlXMKK5e
nNkfGMlCUu9MhiiBmrC/FygtFEW8X/Ucu4Ru07BCbCRxfgSSwvXJWXpmG1HZ94Ho
RI12P+ui23efRjU9zRItmznbB5TXNqdUaIpU0xzuyRtvuXmiyMedlc7MqpYz6D/T
CujvJfsLvkutyMZv+HsFBQ2PiEKVeREpBcd7K0rJRbFWmAL/G6OOPiaXLYrUpC/Z
woLlayncQ7EK5jmMy9Fef7PE6R2LdaMu7nAClUy1imS0NuBPJd1FOQeeb3JowELv
m4xxOMZVSPzXhwH/8prmhmpyS8qS5V0dAkrAJuO3G3CM0JPC8GhLsC5vkxqc84WR
4JNslN6vTLoKCDwU4fMAqc5pb2SFuwfu+7f8m6A9hyfJdiGTkoMIhwZS4P1ratr1
WPUfzbY8PSKPwdB06NO5HDKvG15wpFgZwxWj/Mc1EW470Fb3PzX5S5IK3kLzy24r
pSLik9g9WaPiPBHTxmPOM57mqST2Ug51HpbEXAsGf/WMP+UdVr9JX3+atS7TwpdX
cKjD15lzlHc1pSsY72FtCt2se84qzkmxe1Qaq87DNKXJLcZXj+jlN+T/tJI0ptQ/
Hp1PZMT5dV4An9r/28+lmyWBhkXWaoD20+nihK/q6CoW04T+WoMiQSNEE2itCg3y
Oqww7pkb0d4yzi50ivOThKr5Q+/GRANomHbUCyyrRiQSqKiNMcSLX+WVBvh9kGa2
0ZqLL1joGGG/hk6lLtgjxmekcK8JqAFAabPY2iGKGKHG8zlVRUDqZXntdJF9K0kP
cxDvWkPeCclNY2wX0xQ/KFV0eOVVAGE5/Rq35TecZQ4xZSVb/sYYcMEv3zvV3pB3
aqFQEM0yt2BMUfMQdR6BDeNr16r9ubS0Ij0e9StqxEBRo26BYfE/ujQ8DfZHQ5hx
HBnYWiIyZiT2kaBpP4VEKW+z55W7+xV8lTy6sJ0sGv+hvLvhzK2gwLxGSs3tG/kK
5+1AJw/f6h0OY6wvTxG9LFVbcs3hIjgAtWMrQAtPrMkP6OzRwF9Kp/oWKaP6OnuP
ZiI5XG/s+VcCKPWXB/05UHxBTWlEaHqdVJksbdfVCsdC9QiPi+r8PpXffp8fUrnB
eai1pKgQ0K0ySmB576osgsifJ+5vj/jNZzfKccg8xGF/exd1KXhkyu2+fjB7HXVq
SKXTWnaNyZhG+Eaz8yGBouobJpHHon4enemS4C9mI4pWIeaBcQnqiX2NS5HCZEy5
aEHO1ITvmaqXDj1zG+Qx/m6qWnrzxZmyjcJ57p/zp6ZO7hFPZAb5gi28tEB5fBmu
vnhRHYZH+ch0mFvpyAQUyZZpvUF2jYNq9BsWx5qcIrI4YxidSLH1eyydAIdmpJNW
tpcviddtvh8hyvNasyHxsH68jJl74jLqJX+QeVBoAWtjdeDu1AOOP+t45jh5Uqi/
FxkjhmahF2ZkwoFgRLOoe+KOZgvTz0RGKfaww0pe+IFM6iB6UmqL2q+4znQD0HvH
Sc52l3lAgYFydSsgnAvTAYqYyk6QnzW/v1nrJiKDml42T1cykM/+SY+WiAREFq5f
6oVe8fTODFj+XatsabdaLwHdmcm11sdZIcmwlYPqdpKsSy4eH68fFNa7SZEW+xZr
J9A5iiQnZjHDheu9BqcfdIeq8qxUytwpCpMKCNiGfcjXizckJwkTVnizfEAeEDBG
IJeKYuIHoYZvVhYGVvhpOgbG/jSIgZoXURU11rEQXixMeKdMVNnq7/icPi7bU4KH
dwOfgqyz86brQ1842HUUs15DEDUQGCQK+iCGqeGTA88yQOuQdQV5BZXggBeFK2Ch
d5iZ7ywNPgEaw/pVQrKD+byxfP/zz8fWGWs+DYB7lgTKsUl3rMdB4Fxle/4kfpY0
YryOoGU4k0+rhNFPqvBNN5tl61fEu884DvjBe3zO1Vxf/u1+xrjYY+Ok+Ay9ivzq
zXPU3zqt9bo5/Kt2KEYTqaLvzcUIIqRRTuGlb/palb7K4J9bEF5vsF7x1vdubbat
7cozoASUzb2tMJOIh0Gs5Nu/pUG76PhyKxw3szGSxqPNlC2uTW2+5P6EhNsXyDFQ
q0JptJnasWCKRay+YiI/d7q1aILoxkSRq5jmWDX8RiwEgdtJrP0KMEX3AHCshiJZ
dyqVtgDuhmm5F50u08GKXemnhRQbpo04ibafMUM33Oz4NaFCKqcp3jaS7Zm5G3IJ
BWtbNWKOPJEnz5mU1D6sDOdCY52frpvuMRnn0OGP0YM0SqpZMy+6eZu6GTB5HlRh
clgmkHFIEHV46F49R/Oi3SKyplrLxy+SSv0pVnBJs9wZFIebaOru0HPnSaplcMn3
plQnAVMEOOlKAMLbHKrUeYyPO9dvWekVH7ubSlIERzOe0Ozt3pBEwUSGQb2NVFLV
4OnB+9KCGPjs+KDumOXv768n5dA/wK4jn22O1sbNuwJqH1yIi6TwMMCAADcsL9QE
7d+bMtSKTV4N+NdldEXcWqtQtsqHX+ML4kNc0C8CpNv2FQSSn7pB26XFzcf1h9n/
VzyidIoftsX8NifAWxvdhByErmYi6kYTMhb7hXJ1EThOOD8rXw3DNLYlnSpzdRCw
KJPpwRRAmzLqQ0i3i+zcPS2Ho+s5UrF7zlp7fGCnSMDBxj6yGzc0dZrZHJ+aivUg
ducG50ssnmjQzIDyy0Wc7ZWw966mgKQ85vrKZW6cXpSAGrQlCqqTXM+fjD1HeQDd
lb+ifIB9LSCtSFja2RXEAUXqp/SyjTc+pD9xAd7TpD7bFf4T9GM/HZ/DjOyzisyC
4oi0JcziIigKmjQZW6KU8XcPmedwpICUnM+kPL6uSItUGe7tBv9og6DJamSKgDoS
SLZHzHGWt1PrxgnQvida1H2cRGDhlO6KnmP3Kl2kZKr4qUDVrHhBOuNEEqozp515
Jq93hmV81fh/B8RAFbBh+DVBUZh0/LlVPDwNTKokogLI8mwpSrtcFdQBneAQw+GS
iGrOfTN3B2PTzZos3AxYnc8YTTZAf8xpRFv182firxNYGL3GW9oB7o5Zhc1+bAEz
Yle85VmkfndHJ5EGnC96mz1UywVAKMtaNStTHjmYPJE+1QeumcMPGnPZ1sezIzKc
+Gw+69Q5MchA9yk1llIbXnP69pwIEl0wnLSCTXIHLNRfHXH/KBiDUTKF90dCAZou
jVHSF4oaBtlqei0g9xiGNe309uGAYEf5iKmeOzbqJKwS12Un3IA7KWRNALwgNoZq
ZBBxIFv677kcf4imYOb5udQqqjhRHHVC6T5NN2ID+qlkAMZSUtQZAMFxp8Z5G7T0
t6qoiRri7A6r84dOeL1Eq7p4IazM+hyfdc9JIFcS4+IOS6dWwmHqJ6Vfs3f19LbW
hy00nH8gP/9BIk5Kqt6RCNKmpVB2gO5/qaKQZtAx4urYeTM8KLRwelMz3xC5gEJB
AFw9aLvz39kKEP4Uy3JhqlA/I3d+ulKbL4W8HdowJFK7TH3g5vosocnrf2SUGivw
dDAHsZCHyuNMi+QqqRuz+gFwRZccEDyVE7oBFN9u+6leDD0LqeNXEFztc9xPxNDP
BG1a+fd8LJRy7PsuEBDXaYRKOWsQEGQcv9recu8tJfB6dnii2vK9VyaIIQ58D8QF
xyraM0JlstZ7PIwQIwNZKX7dkKnpwhcvrSUVs4z7/Y4ZT/BbtLl+hNAUsJWxmMRM
fa4TfqRAs0cr0Gk28QcqL1XxYK/f+yyMN8fWKQUOpbdguTMmYywlRRxeO3jFe7MZ
zdvB/4rwC+wp0nKZSeJCfAn4QWGUrCO2XE8n/pJaJ1LPgvxFiP+D8ADxZkaMUP6Q
DXWdoXFZgT2jGlobT0LGFSYZGCrAB+OgFu/h+C4EcrMjZ9LAJbaaCQs/Q2UPynGl
mBvhi4+QdoHGOWSFlDiMv/NU627tA+AtmeHZX4T8eIpyKlQo9NiZ3dDgEmDy6JEM
VbOA7/M5aHZW/ZdSKGsujtlm1nmW7lwuKnEjFQyADxI75ceT2RNtcw0YvERiO2Sd
zAgiQfggDwNq9TiMferShcepBQFLuE4ls2YHnSzSa2dAsws8Ytw/nzfYchIBIKuL
25NEkihp56BQ1lSYCsH7oUxtTWyYiEdeJs0wS7EssW5YqzexUylPiLF1kZZKa+al
BqbN62jO/ZqKM1h6x9TCf0uG18MKOKxrvejcCoV0iFoSkbMedhjbxOA42z0KRk/N
UTG107B/JBjJfMea0CxyreIIerMez4jSHwQUOkc46s/ZlQae8ZQHRecS+IaNRZdv
GmTbmq2leKUWQrWxiZcIf0Zx4LS5fdt27plPno3TArsR0PA7ySv48S4aXY6cEjsO
wyx6svQXj0LleCpe8ZiW8rKjAKPfmTFzbZS0rqbm49GcmaayJMSFeHXSPqeKt3iu
EYuo1lmjaIEue9hEv2gqpLhLt8C9n6mGPmo5O67mJrHmBuubtgz4iaU5YGSenAJy
FwJRrze0FEonJ2wrvwrCzTw+r6rm9o9uW73SJaowIv9sk0dfmE5BRDHqo+2z/RJ3
a36fq9Sf2rQmadKharmRxm4y4ZLI/YqJElCVMvjZw+NFs2wF6LEALngegVFVMOe7
ryNaWXsLF86rVhweLJ4Biie+ILb+LoKJrHSkExZgcKoo9sEdrg+qzsPZyi8+xVg1
WWQPB6AOmZyudfMaNqRcWgFYYzaKqA6FpwcPvPUGrUSL7w9q1fNY2ncGIqifrgKt
14Yt/2qdzjFLNHbvGjwpzKYDn03B77U6MzEVdg3Lbvr7+9NA7DI9eEelxSQWG6/8
rp878ZF4GtfR0MLEguqJQBsrcN6DZhnZ1rXk8PLQxkWx+o8ZkPl8ToyD0sFVhR7a
KrMulN6h+DCBTxXMev+K7PCtnO7s2bVMEqJ4nopKxBlhOsX8oyb2Kjib0Veokklb
+Nxf1gdIqkYYvXgL7Fq/fgNSbtb87QeshCrKeey77TpF+SZrt9raHnEcITCEUebe
iNL+vAjYSUkQEOq/Hzoohr7GDfn3V2TPBUV03gi5gK91Woz/OPpXSDyPQlDQeX1X
eAftOaXw7kuQwbZJzDyK53gaxKIpChGkVR1iCJEaxUBSO6q9rOW5AKk4qpZYK9Ia
eLBfuT5fyVj3yw0WCG3Tvx4gGyCod1MpwZzkQ06od94/8h4tqeU6yVP4G0oU+kMr
oQud5aGdZc1C2ghvJ2NOGlkNYrWSGrEqsxIhNoAAnTT7pEBNHySqmbamLWam6Kki
+4prSGTY34fMAIXPwv38WPrm/z9e6Ce+54nHKDMYyjzJaKOChURGXagJgoy7hFxi
yY/fbRKO1z8EDgPIT+BA7YP0uGwvAiYf1JZy7XtaFOul4s5IGYNnjlwHfJmclDeD
ttI53VameK8IkoICvxmbePuEqG8IXsvXsU5UNkBcQ3ooc+29rj1ADSTyvdRBJw8n
ZFM6JkaJNEIGgZk9OFzv0yBTCoNFIjoDUkqa9MIsTmygHwUJgvhf1tOjqLNaV4fS
maAAZOizwrha9McVgjCErEx+7rI3CPHekjaEWqvhdY26xy0P7I4KN56vGDZBZNx0
wVKmFOMPAtaKeA5x6hUcoQqPsNYkOduOkdnGq3hjSF75e6am8ed09NxJmunup9In
LZI8N/4qqNLPYKgzMXeYRGI9uk0fSubMHR+JhgSTo/7OWb7FMNh1ucKEvbHON4mJ
l+GZD5lXgK1uiiHwUS1lnfKMgBBGT+xVfcOok2OVrb5eXhFEVc6a55i1c2XbJpPZ
69YdbyDNY9HnwD3kBsJfjvN5lhN6IYbDGMS1KzZ6kJKadZHN3mf6SaAT92wqoPIc
EfkOtR88kL1JhK7ykqxezZPUWm8xjdiv0vlG2ncH8S8LPlBpT9HQ8yc3auJO8Duk
9S4hyeAWaHFEi+4HZqwAxKA7QT7pxteti5HPjyx4mMjLzpfQzM55w54v4SVQ6pmv
D/zLlpiwKc1HX99totKbKVO81zQkJanILupi1OU5HgE72mDJQgvR7REjkAxw6BFO
l4b9ffsOt/jzkQcudD8jZLlEWwOmzmW1MDVLQR9k8Zfi/v+jO/NbahJwNPcR/NLK
oMGyEXdL64lTeAmBBGKKtl2LIP9eMOkuNRar0JxS6Tiq6KDVrPF9u5QAJUW09gWp
/J5OtNWZdKVvsMbl8EJSfoSjKKPnOqsjCc3lEnBqg8tkOl3wHDcECqBvbANeBT1e
gI5iE6KSR0t5K57H1AH7iQGJzirLmAPMHO0V1zBOOYdLl2jh4pcTUzgwLfry3lcr
wgYj53mk27A0uHZji4tZ1Appy9DORwSPOosWrLyHgEijhjvGm23L4MGznMwKYM0Z
13/LTA7IUNhyrjA1wP4WGSzj/jdvls3hhnQYcBIvJkNa5jeTxn6a15sRWIo2Qtpx
dHB3eGTl9e/jL775g0Y+tX3haUgYK3BB5VcudaqYuJiv4EUA2ChdT4yNUo8EyKGp
7fUERQr0WLy84FHPu+l157oC7KPaDscuX6R9jPh8yNqR3n1MPeQOMlOs1JoKw/wV
/3XuVuGq1k1If7yrnsD5fctjF1jQ682mFrAC9cHH+5H2/1X2/L2wc+5koG2vHJkC
bLfPfs5Sm/585vdcI/5FQswZ+BrCMHsgj89nbOEeElbAE0fS3pTEDNVB2lztOo+R
uwmZMmCV4vW7rMu8s0H/KWJ33UE2eA0o+5moptdYtRGEl9YBB70teYx/CJ0DttLU
ubC2HZRFcblojtfgeGmraO45Y9M6SLLL5uJ1j/9O/FT7nk3t3C7UZrk/M1M15caF
VpvARMl23b+fhFW42Lri7hNh5VLoCvtwbxzvRorY/RIhmi40/bcJrNzuVq4nXzW4
hGhcpEUp47l/Zy02aUpYOuTe1O1GJkBo5nkbYMtpnSBsBC6VYnKmwiVQZqPhvxAg
0dmgsYGAruhWF/BPM22kwMjRjvZcYzMvTBgCmXuBh0hTJn2NSffq4FOAynDM+RhZ
sRalgYIYSrfuyFvFPZJc203JgTUiJvU9SDESJdY0D0RuAe1OG8fVv6oopjNHAbt0
3oznw/xiFOf8vyfYVaMyFj7r3folBaBPZU7hyTXFO+j3mvnwsqvFHkf9BlVqGZ1m
9wef2dbG+3Cp+iBntsGb80BT+AbZ6Cs0PHi9LV8sO8pP6doUByHyR7mkvvBhlPlH
AQRsAf7w02luiJjezM/hW4T+fkaqek6UPeSHE/wb2CpaQgtYd4CgdWQTdWQJoSgn
No3Vis3GsCuIz/u1IsUwprWnQLiNtt35W7h6RVbkZ2YlDHYAQ5pMDPwDe1F9VCRC
RxO2WurRzbKjnCWFuhdjlx/lU7Oi0rTMuJT2gCIYpux+FGYRqctXMVQcobLtBgJq
ohZb5jB11DPvIgeBNst0Bmz7M4W6+z6DWOQPAMMHOUuy6p70r5nHY9Uwe/8tDBZy
O5VKpdjymDIcpulCmD0M0WrFIyufo4l90T9mm3Wb1/HsdKIkTj68qU7NMT+vKg6H
Jb1PsOEC/7wow83NnNg4vAsPkTJOe5MqnvaRDsQYVRjCwxuo2GsabLuT4rWyOJFR
Ly+79A1fNtoNuKu1bRKFUNf3wXa6Av1xW+0fOhhTcFPLyppVI4NHCjdw2hai5SQd
cECWcWN7Ut+Rbzk0+eVpKxBsipQFhO4WcNevsqDaBvjm9frXLLa41p2U8BPZ4z7a
kl5exg6IU72zqhpdXGbXHlMw2vwQ5LiGAkEbgXmkXO+EFB9QV0hXnvOKsrFJAqVV
hEgT8/YE72dCv1fc2NTM8WZbVShF0iXTaWU8PpvU4KhXSQWrCqzVgzMaX85/f1yD
gonl15YzBke2+X5wxb9Ay5Vg4s0iMyJlmyVcaN1SpLxu8ZucfwS1tMAKLIQge4RU
QV/2DHHh6JfwjX/habuABM1KQFTBqh3We8Js7CNaj0M69md6zt5p+12Hn2UVg3ZC
TFzofr28jTJbnoEsaVaBCvKzy6KVzvGS7oBRqAXv6o3O7PzkKomSKFBe57drGUoK
77zsqBn32AgrWdvC1GKe2axqUvPgQGdyeShxGG8c8ER8ZditN6Ywkay7n1qiDeYv
iGp8zcecab+WE+WOAgmLZsxVZNzzkZ40hS2L8lbwxpgjJ5LVeuAGLbZaYaun9bPS
N6xxGLJZCNhg+XcpaCLbX71xjzTXaUunIna1F0AD8uvO15LcQFMt59pG8r+qTyJL
xbkOLgj8WycCsE7WNWI2JbZpdw+FaUc/dD4XGLcSgW+WiTBJ8bYw0iNkIGnRfdcz
TMzqcc+cnlkb/BkeR9L0n6XXGcOvvWNsG2CxYLMjbbfkmVIF0QgURkB029x/XYW9
+AroFpBUOPNWpBNyaMMbTdWmzLRKg+cJxfr/hN/WiqW8+8Zbw21KwD3bB++e0ikQ
9+w3PS3Z8/oLPxHBICgfiBFVfW9ajupZzlOxfM+/Wb4T7ZYfWIjOg7JY0P4GC3Hv
BqxbOFGT2iezigrgeegHriwSgfZm9pT74lBG7MWvclbKu1ea8R2E9IZr50+OLftu
vRSfSnyZG49nfmXTEF7/WMyqAHkasRghPFOXms3LADauek727cM9BWjXgg7JuT/S
PhizODfxyk7nAGTDvaJ5nNKo8nsploJ7cSxFGAVOiX8H0Imu9Ie5qik6QMdLC3PZ
3zJLX4XQvJnoQzu0Ad4sVQEp2mwYEegpgg4dLY+6VLjadUmuaSA0UTQxmv1JAAOP
4RyPh6quFvg4BpUnjQM3uXN2b2TSLSLoWqv0wT1PlRILtRYSvauOsg2Ar+w3Xm/f
uXk1QHsoZG2yoSA8abrvROF8b4auuO+YPa3SFO+PYeeIJ9cdPz9aEAj4+TF3o2+q
L0QDthcW1cM5+9dBNZ4VE1liZfA91b+tC6sIrzLioJjc8Hit43rLbReobVIWFoDf
0sZrh3Lq1ucV0J/jhbQHZQWQWbji+P1srn7FdnD/Ost6vE5vdEF/wwkDictJUMyp
A65GoxlHSy12feL63kd5gh4hmta/SKul4Anne2cN03FzrYwz2l+DHZp39dJIb/Ng
7DHBWSv1uyH3Dv7kHvQvAAvfpBVZPb4Ssbp13JlVFb3dMH8HNgYAFwpm/PFtnQ8J
L0Jozeziv88NgFQPRZlW5CDTw+gznkP1aEr+8362ZvW9gVahXibV26lpQgo0U4r8
vI1mOITi/clNxCcUEjjcZNbimf6TAX82o9e6vQFK4lksyPjmV2RIn89IejeCg5++
UezHzXtsDRDr9pK6+phXW4qLR74iy8PKRuNoFyLrpDvZlq+BNTjRPbDWl1iS+w0X
A6XuRgxtNA6m29hlhDnd2PDK8mjpxPD0/Iqxve5KfR2WzRnao+DGcchooOqW1aws
z+jwZ232vF4x2CJJjJ1amHILjTF5cs9y1AuzkpgppFkl0Wpl6N9sOXCONU1RRzEb
pkvckUPdlBT1HoGDj0cpY7Kp1a7XXlMpFknwLFYgZDZqZN3joF8K1WiIwX6jcbsY
sRaMMRDALcXGo849sH+nbu7RRlmd6rrXTP1sWRRwio3KUi9SttI7v1dbPt8pD80M
dq8qb5Fq1GqK2eV8/x18DVGNyNCRXQJmMr8Myml/51viHk26cL6exey9B+T9Jq/S
WaZgV2EIoIN1Ia46IHK4yvWNvnunxoabD5eLznebECFG084LChSYaczAT9tB2hFV
8AevY84bFGqt02g3izbkgRmhwSMl3jyhoo6TJqTEFt/XRLunpYgZHckhjw3McZjr
E6wzo3UUq09FRyrNRupN74yUvY7J+lAecZr2RcDvpjC3qe/b0EupmxozuUYyRCRz
+py+C3KC/G4PbnoEZh3yGQHu8OIRH2QKe3+qS7Nc0fml07gtYk7ElqVFahOeTwon
GDA5Cdab/uPZF7O8xhT5fvtEuv8WDdMiu63Btjd0zDP55wLykb75euwomH5V7h1H
L9uhKQduDxELf6wIoZKJcr+ivHCNs6A0qC1+ef2Wr/D4iA3VZtt4/rADKLiSwqi/
Dwn8O1PCWtpSR/QZwrYrjeUbYcS07YJN5R97KZXOpry2UhYBvWGGmwS6AGUV6w/2
AygHUfASr/y4XetYXkPbgRzWZL6fPU7IlOkGdd43GGY21/9UrwVPOrHIRm9kPPhU
Qbsok8HHnBxfpQUXxSwLUjBLkYxHVTCM4jR6m316dYGkDmLRNrnefU01+sv+U8Ev
13zSc3vl6QOcXD6S0+zt8I02l+g0KbAJMv+VNkOHFE4VDM8BQ4qLSkaJWaj8Ct+t
V6d3gHpkotTzsG9+Z84l3Zcvmol8+14ijm/w7n7PdXDx7xKgdbKVFfNm6opVxWtP
XSWQRrlTgiksUKLvERx9fTvYBvBddUtA4E7KU6HWKnMAvruPtcSJ2cYwHfRoatH+
9HESO9Lw89rBZ03XuGzYvXBdU3Mzc2MpB0zICGjsPyuAERolg2Z1wE9aVrsh9yD9
iq4oIEixYFuwZ6jHkBdGX87eYxo2Zr7b5QVa3OttRDurLvjnRbuEtuVuYeZnHd2w
FhUdoitjbrxLjDxuW/n24nuA6hx8fVNmAvA3+EsHwq+iOSCgBCXdFn6oUCo0KhyR
2GqNq3ZVMLAFOuJ6woM/SNZNsaiTdLZwlO1VCSkWHWlVoUh0vBIFr0gb6j0ySozT
kVL0GpbcLjBC63iP3q0Q2QbQW5VgVslBscdMtabHnxUkUVZ+rKz51Azk4FpTn5lb
Q0wFGUyJNDn451YJ4zMZZNMajs6YD/soDi6LituJC9R7ZWVxoX/DmFbbHoujLsJr
fzWmbqtqHzmJELgRxbQOmTKT+o3sBWTT+DE2HHl28BJh6mTKJ0rU0K4ky0XYV2uG
GymBnxNR2IunAamZz4d99UVWk0T0k55c5EcTA+xv7p/fnoDJtgyjTSis5sWWB+pb
DxXEWk4qaH+eZOQi0umYs4lajS0W5pIKn/erhGT+RIkpjyXnZ2pfwRo5AuGgKGpx
7fBW6Hji2JfMw+uQmkgGBL5F0HFMjByj/r4fiV0frxZTPvDHGU3WUdPVfQlajvW3
/ewbcJHvEUzqgFcLwVe4NOTeJIAYu7kvx46Hr0eA0ENPYm8PnJaVoavPqMZzvzun
ywXJQRXXpicAimfOYciTJ7RIJi08LCGpAnkULu9k3U4/VgeuPpenf9NsAlXClvpW
GVCBMbh9nrEz3fw9ia/ieH+GcSeq8U5FPJn1x9Mldrd8RKZCfdpIzzRX7WG44G4k
Ywav8J+uI/urdWq45DDcL7++3qURoI/jaWVHtCeQOD4Ly0D97jV0+uBeBBkPzWHo
LycP3iJ0rBs2BevQLGj2evqlK+mdv8f2zUxN46Kob2ozbwlDKY9GnyhYiCc3jlzZ
Z42vZK21jme8PDgONVnUFd4+jtaJq15SjlMK2PmXUEflFQUKfwjxtNh6IIZEVFjs
3zkU5dVIYY1OHHABIk9YLSAaG5TvLP+zDx7LyDGAygoVU04GQAL1vIgyYIqrCdWl
SO42SbwhfYab4hEk1BQz42SpGX4nJ0V7df6g37DVIwfHpkDh5oEubHgLhy6T/Ren
z+cuuDF53s/s1pLltLEIqqEMvYzITe3BKF0bPOIDxVyfwTnwIfZJBJfZ/HUZHyCl
XDPQYRHoYXda7IPp6Qtamt+xtT+PH1DQf1PKeJB5i1j4YIFQ/7Vyry0I5NuJS7CR
WVycWENZPHIXbd3wJgHEl3bUf/rqek12ekRK/NGp8zhTA//XIupoGdFefoxOuP9m
iNKewpvtYuCBUlWiLLQdWJLAklWi7FNxpb93jSFaauYfNfX+32UJUa7JprJQtoCN
IcrzuAQvrVMt6ahoq0tlET36yQ+2uWOEcVD4Xc1gWLdXc/JXTycSmJMxPBWb2foi
CET5D+Y/z+lLRzHvdtsLvpLGcIlJUqdsEWUFTjAFHk6vsf7vSUpgZWXI/HScHg2K
Bff4zBdQ5VFUiV+a8CUfNvI3npCva84XVeVZZ+22C0M8L+foYDOG5AKEYknCB7Su
WQ/5s5F4QOp2dVIBzTXdHH50xJA0smWCXvBJu9lp/ybBYQXlJEBGg1vKb6UePgna
J5gLWSsQwUC0OrN94aTlE8ngljDyyjv1ulKhsbb5O/mF391lxzHreT0zbPQ5pL3M
K+H71Np17YosKHlOgoR7q6yyXSXCnMZnaf+101nxUEcF+UaYhvjsv6AMh9fiu1q5
b/66ekLCGcoCpqtvR2OPjMCSlC7iULGH1OZxSFOAOiu2Fy2uDhqZ5Tsetmi0IZQM
t9Mk4N+yS2yK4p97cT2vD+8y5upr8oGiN1veFFPiKaKlpXkapXFRay99a8eRbCw0
sPyu3odAIl3I2/zcEVmc7k0ILU1gxdi/iiYSh8/4uz/AeGoIrBMd3tc5slfyNEB3
/vjAyM11yj6GIfYMLAZr4SfHPGIa3F649teJUWcYHrcs6QQUxI4wnIFrAv3snHgg
bVJV55DcJmvdPaMdFfOvIVQ6rCBjTzLbVVshMfBKdc1YpJJ2p7+LDclU9Rv2iGvH
0BvmD5Ue4DA1tnkQGpest3uu9s8b7ERUA+ORi7dAyKBeDWDESQs6OxnXMbyhdMEJ
RVDWE+9aDe3GlDlAKbhna2zCC+Tc00kgU2RmhV/8D8ebXvyFJy/eVf9iy5b36Rb5
luBQw/SbLD729Y2gvoTFlRLOYm2qkq4+MGLCqKyFt/sVl8n/IcS3EqZt913An2/Y
w2BKwdX7Haw0QYb7gn7fUJcE2EZZTTkZiXBhzYSWGHdhLCisFydFuCEvQgilnnrS
aXLFnmr2mjv9YGznjyZLzmTMwzsEA84j6m7teistAM/jhEIJZLcp3S4QzEWihonq
Efqj0bcTH8A+zaewpKRMGZ9nOcV9KaAS8hAoKNBwD+SZeF5HdZ7++CFh8Snc6ZVK
K6G7X5/F6Rs14j/AM1fh7zkY/qneah5eVpXV7x47Ifa2TPXRJhumwHIRFxiHdK8h
X6z11azWsHw99E9Gu/uhneV8duVktk0XeyQu/kaMlssjZZ1MIq6J3e2oRkg3iGO1
e2xKpDGQOS9P/z8hOIaTMsCgWfpNxsn8+pWuqBoSdBhZPSx5Vw1cCJTB3Tmqlvdf
Ct8ogJ9WIuIiGprTLJ9ISPhAPo4epp7bkc6d/omK1af26+wZQXJMv59an7e/sdBA
8vB1p42iKQ6fUxtwwW0nKlWL6mD0RSbG7UPw86p/6oFDqF/6lPhiBMhHVc1MQCLr
XwnlybowOVVTFzI64c1A9xKkVOVWHO+FMLSzS092Rnn+jHGNgetDPHGycw4+zd+G
6vRCb9YhqEXiBE6CuN7qagRGpUzSrcO9TDeoUHuIBa5krv6V95+geNMTA+D+vEq/
FzgZgjXZOipYeXF0KUvB+aAG+Y1ZytdczExIeqwukK6HPmLoQShZMkMepHnYrddf
aZKK2uz7vQ7g+Eg39KwBr++clQRXKczDNB1DzHtr/OUnmIGiZZ358d92C5ORdCcg
4jy5xYLUTpiRS9j9UqsKcpvVLIgSHo5fhRug8xMOnJdq7W/1f+KmF6wPJaA0+zHD
q939tU2nJaQ6dEvI2oOcdjJm1HRjxS6wg5/2K9r6zd88VTL5ya8stcIBGwmewGWd
WSgJIT0IJbSoNXdrQGk4ltFJlgYLD3KuiejTQB90OgaYTUCObxNu8AXAANJPmsme
I4t6EXMUDBCgS76d3n9kQuxiCLoHSzSVx1drLb+dqdWEymCku1QBSdUoEzABkJcX
CdHP6/yv7gGnEzn2ih8EkMNK1sqRNv1JjfmInw4FT+/mLWCbRVyTKqi7ZMEE1P6r
V8lF4okyyN38qN5OzRZxmCmAyrJc+lgovMULHuTsrXYYP/lhYrSLZD5Iul7KfNsV
9NiKyb7VJyn3YfrF5rYUnmS889bxI0xE6ivjU/yJExKm1gwwBccp4rtAvz1SWveo
twVAJtSTuyffKmHu85g2EJoOYB3y9TDBZT8zpkYCo4jrHx2ZS/k1HeYY2wUJWieY
nO3lMdZCfzurN+fQWTdAbkyk0wQjfm0D9L4c1/BQwvznrXHrfn6Nmt2OpJuEpYTN
0J/6/dcv7yICLrBg+Jd8K5Rx6foBt4/tp38sZQJCQzmc7u2kE1+UTAH1XO0ZD8kj
LdEwIhFdQSZCVlMZGQ8lfGz76N4hpFH5T4q9b8uvs7AS+IrL1xqWoTVfuDVpxWYs
WgjG5bGl8ObJxiXJLQ6QoUOyJmUQoTSQSvCAew5BlQhIo7RV2AsXRyz5W2NESphc
w+xNgDwRxV7kE5BZEogXKyiyS1UBOQJlHo7IiQm4eYl2CBcnuySLplaBj3e3ys3l
+RhiS7J8X8RkseyrsVg/m0keyvIC49WIXogdMDXAzNmcnZjT9GgO1cyhXAoezj83
sQGLXRnMn4Ga53g8FpThkRdtFt0WdIKlG6lnigOFKEe5iHLOwg4H7d5neKPXarBY
muDKayW0WYZ7On6ailuKzH8v8Q84GCM03Rt6tWFvk6c7f4A+nU3+75OntQhbsuN5
6bXJgrEUtTWXGtD5QoRYU60+Zvxlh+Jiu06Vr4xujbh6YzmGLJljdevWS0oDkl8R
UHg5pm9EanY5oFbwNNzHKthZyCgIffIiK0l+0Hs4xPwOTrVQ1sGYZ6ye+tK/jM8E
p4ffC5gxw5RZSSs0C0G4+lef1+2/je41EYFUxqFxAaRHkBYEI1gIHoTCALxD+/l/
AhfuIuzARCXRB0ebaMUBxp+91TTcqSepcoEqvnHcxCgRkHVFJpt1D0glB7CBGeVh
AiKfxwUfpz/2KdWzyw9LnYRmYm+bFqpYo8op9sICmFzY5X79O/eT/7P7u8mLRhxR
n/d+uOmt+5Mphic4fFZ4is0uetScO6dPIqGrjsIIoB5FtJeTMDWO2TqoA9iNRtBS
3SvMJDlrkLXKczG3Jqran9gxuHDKAaSqUcM5Kw/ID/YPNYztaEj1kT1whh+igS/5
OgPkFTBO3sDJ2g06onsV1plL3uxk+nmovt3D3cllRrc6gd17uUiUiZpo6SBqJEHI
oBni9aP5Y4+ewmIg53DuCL0yVHjjPZPUWLyY86OAxWEfPJCccLi1/Bi0CXZaf07A
uBkMMzFsDBPChuZatK9V+bJkdhpSyUv79VtC/MvStop+TfzABod/Aq2NY4F/8as/
r1Y51mC7QgWSRQ0LTOO06fwiQoQFiTphyAXO9ZaUR51JWZrGPm16cv9gs8Lphi53
+h6ziMumtp78oHZBs0V/m4TxasGsMRHQQmHhkEANzUlxV4G3t1+WHvntjYxzrf0q
jIUPmgwUWKy9CWpsxhjzY79wgSrXrxDq4d5aJi3P9NgorY5RUrsk2h2ko5tlwGdA
h7BYXnfPPPriclsXnEw8fXqGChDcvhbDKPUKyVh/rISXUllPr55gBPAkztz6oi/e
hZcI1dbvcpk8i9niZTbe8gqejYI27HcnKvaZOv3oI13mIqiKH2kNLeKPvJvZZA5A
Qdo3PSAsL//zlQhoWXK0T9HTYesK4nTBcSQA8DeMjyI7HSfVCtpKLmuXOc21LIFR
OCwBEGn2pK94IXQLP2RWKcjc+q7o429dAAg9rVPpId1wbXt4odsZgy1+xAS3grfE
TaKTtPsht4+tH4H9Er0ePapbgw/gCIl7DuVRr/LmPEDUVgjudXODY1RSLv0mdLlp
bRePqXOHI7gRdJHiuR1gPNEtaeKarOuVrPQXSTT3SFG2BNO46xP3zH7qGkevfliG
e7G+vqpXLs6oV23TJEPlSAVkQ8NQMXO+//SSjx55KYk1wSeF7VSjSSsSJKkvhp+f
gNKq8NQI8chrXYZVn9763RCPm1fEcKBYKksOaQsdzokPtLAl1t6KWcLJwIRRnNNk
uLK7eyy0vFKFMxNrPZdht4TYcSGUzPgDekAvxRNbDvItIZ4ofQsvr1eB4xNQkPzP
ewH/YauiA66SGP4EIVmcavUKTQDsptzTzezYLzptkd85onFjlgeQogdWQCAP2SjP
SDtju7FCost+/4+cx1zoN9E9PMcP6XKiQFoBrK+wsbJzBXKSrov8kCc1ft3HdCYl
PNTuKI6X1dQrao8SEWqYIDlSs1pbYINn+FAtGr6hu6yWEoj5hcgpflI0cJ2aocIL
tOqCJg0c+NqSQDtlnG8qHM5wm6YK9lIPrXd77M8uTca45C4ywnZ7S/Ou5W7uf4Zy
kDWabx6FviJVC488ruLA5BpSyPOHF1gfmaVqkunPtnlqM6EQ/LlBZzMqzWO9Vdly
InXPOLT4d/8pihM+hhfFDjY6pQw7onj1LYizUWAiOyPpRk1E7SyrdP6so2urxuPg
4QyAeuEw/6mhRD5XU870usnG8X8mgqOxbg/cpxHkEYDI3SU3dzpYIDdinGkX/gIK
Po5FXvwHVmiMGJOUbQARPzh3m2E0MeehE2YyNdgH0Kk1BhQiWdtT6UYjTAsqWtlb
gE0SXSlrFzVn3LOweKmhCgXDqQoz3A05pR2w3irsnAyBUj6tTsZgPBTkZ/z7t2XT
q1ZUD4POInqpEYcAxseKOUBdD9VYUueVPQSGqsRQc3OQyn5CRFy87CnbJx90F99g
EQWa5JuE0310EBYYjBpWayZnb9Qb7YCOp16CAuUV+lC16EnDXGlhT/gaSBmTkwdc
DiCu+6Ftp38b7LqCqf/OgDrHZeyI1BlzTizlt/Us63+aQIK0kWVqFLObk1b8O60x
vZ8w1VnP9QgSdk36MOKKjqD2l3a72k4VhZ6L6wRvV5QxdnWCgrDs80zFZD7+tBRz
VsR/yrFvf1AmNM7ay1qgXh74Ok1jWTJlb3PZOx43p54Gd9tw1xuA5e+xrxlmS+GV
i/a9YkFwY02XdlvpIlZNaNDwQ5MjcvMYXKHGob+3A8Vo0QMDEqAjEdEQmi/t98Fy
XQg2y7zGIChaFneLEf0IgoPdoVhaQ2WlCmeSe4b6cdUQHJR3QOf9Dnou2T2KOiTL
+cpURLFKE9673VC4y/ZsJ6d01MsiQ+Nnq2ZJe+ugoHZaAfpDMbb4aJLrOTodkA3t
8POU51S46HS198rAJY30SiTXT7bXM/mnn/UJr7xYxvBP53iV1Dq5itCDibu8YFs3
TrF114vW2P4nMZWHKzHh0eh8zb60DIuQBZohCvY/mxEacQ07RV2yz+EwUEJcAB1B
w/l/ruiLb0UeDLXA30hvmzmRupUNnkfXaMIetjT1C65aqyCYzYlDsfA68FuRlJ3q
I0ZCJH1N1p9kGUzR2KkyBSHDBd94LboHxudKuJQCTunXOOZknlxJOlPtOp6b08XG
LFuWmU0jpNiMtEFqnXqOBamrMZKwp3fH+syvkeRw/YDMTcuxpahS2PIkVRYb8BKo
oPyynTAVTfHfeAtS9WWzd6Gmw+ulSiYivzOJAWX2jaEm6PPZF2kh1YRbL+B05cV/
H2aHhirZ5XIj2HDg/xFrzypnROEZuRdk0Qgw3shEOIvQxzCkt/ni5POgqgityp9m
dJ/JBcOYxznreOhdNg0heY1VAnWJ526TZoOADcH0mtd/cspdQkB39rf+8BAGwnnS
p0xSdnn1GJKpOCiggepkEcbiFNPiGg/2vZz7yFP3mbu5/SOHuGPymCFFObgGV5gL
1Ja1Mz0frHW2EOwrjvtC/OSs8nqPZx2IYrBoCBmbEj9ASFMeGKMmxL7HHm3H8Izh
JMhNiw80aMjLXH3/7RfxWfP5u+bZhugpAeu68h6Ghm0D9+DqOFFtzlZUIvVi+NVx
XXO9JUugyvVtVmBjmXZzIMZQUU+4y62z30R2dkEEf8TpYgtHWRS0oGpuInrXr9MT
NEtQ8NvqCQ+PzLQ7+0lmgIZbW2V4OGUgORKSmnvGAJBc5GcR7Ma4jpRxWHqu5Vzj
elUYdBT1YLd2YfOaLX1V16DKSjHVZP6/NYCnyUQTgnTFF5ke20QWDFuB2EyZNlak
GTIBDJUbLMLvVpghe9hv38F14TiD5ERDm1RuTDAmmquYWndDYP7Gn/AHA8cJu7h8
zwdenxN/W7rmUJKBeMSpZgJVfcYfRsMbustiHpDTRzzE9kEORLIc1ApuMbJryiPA
AOpt600pimIbceQutBvcPKzUtk4fGdyEC226h3VbWpHYfi9DJBmHkWjL3GGP8a4Q
rF96Panz9VHuNPhUm42ROONRg4P6IKTpVb/nNNjpMpGrRFnuylBCDRvWcZXlJGq9
Hr773YPRdgGpu8QaLucXqo3oojA2Zkcxs+yQb5wFcn5RulXKqsSOiybC5QDxyulY
ZjdzsAd/78k+NkDzlq1NI847IV+md5ahrLaAYFj8Effj04VG3SybTF5Ic1XPpzSp
pBlyUbRv51qqfQIOPwuUSTF6pcQ5KHLX/ttsZpXDWRW1CvS5aGLYRHMs+0uwzCoa
k9ZupuoLvCNs6/56z1uKpv8tkXNvM8irkguegSuZLppxqaeeB4ia0joCIOfNXX8m
4/jJu7svrvlC/SxowM4xmBLS5VnH18MSlJv467NKW8eeLyHDWvZTla9Y0zmH8Ayy
sXYwgrj/ILmMZ431+p85vWSgfcushYym0kvRIgpzh4+I31D7wBUa9gduQMpQMA5F
RbDpdIs58jv1qBTcIxAek86mmRWD7O9cQzKkNOChhcDU9r4tyQNtERebfYymZNzJ
TJ65uFvJg0UVNKp2uRCmlOSd/2l5LZxTuplxmOmsVF0Aia1V3lLFezKhpWpI56gS
D4uXC5bQg41CWeZY98SY8EgyPtHCOXb7QajAfN0B1C2eXenOjdUUw+upQjmZ/qU0
L84U5/kiWceIN8HxwQNUfV22mXqSwAvljbAr9l6AsNE9MJfc4Bfq+Fu1v1/83XB9
g4A8wCrXQitRoS8JUMhbGn+1ItBqyqxxSmNaSmySmuJMoWkug0UrffFDO3LBdSth
QUU6K4aMewdTqr55T43V1ZLXdDSaLz0fB/g1VxKO+sW4uG3kinBHByTMK84Sce11
wloMqrzoUZkVf8W8mokzuRWVpmsNTWDR7jwSyjpQsIpoAvmNGGpiDImd+R4Rg6UY
lVLhWYrMxlLXhW7UsAK9v3Sd6nNJkenk1M+GfwhRU9cK+/8NUwS00xWH4r7zFjoQ
ilHwSc2BR1XrWwyXcpJo5MJNbczStyWyrQCysIBdeP9N4RHA/xSx1qa2wsiKmgoo
fKnuvxqiC0/Cts88TeO8zw4KhIDsddOsnia1Dy4GaO/stboo8ypGYzA48rJsjrJh
nx7tVx13BhEBPEXtVy0/4wV7pXaPolH33TZbfmznGTO3lMXu6+efGF1LPTZ51Ol4
vNB7udPnhxPx8v9jSLmP+a3NTyPTFq7dkJj/XCr6x6fRxmDYAonPmcEzIWBQvEhJ
0ouc7T4fXk8jczbT+SbgvQ7EM8SHxqDFfhI6ZktzvwWt8RTkyLLnqNaUvibD1s2R
MV5ljDPXNmznkUOmBhI7LT++KZdsVg27mYrU9IdoffQ7XPxmjhgEnBOQkXc3JDHe
61nNDRgEEIv9Skoe8cIRyXUh4kibzejhSlK1XkHRb9Dl+Hn9Xu6XiX1HZQJAIfbK
p358ZIVAVfPcl0Bh6wHgMPHlv8192wPBS3z8DwpN6H2/iZthnlc3gJX/xeyZsRrA
MWRKsBGZSG8qtwYl6sd004Ikop5p5TzhprBLeFgL+xWQLjvXG++myFjBqHWfvSLS
7Q3MfeGBZIcKRiPEBm9y/hluBTuJZyg0D3/wX1OKc4xSkMNscw4q942/1Hekp07W
Uf249lQX23epz3IMgEO7KTXiw7lNP8QeSfcZ6UWt9w0e3rVdrFObnptfZ5ir6ZE1
JvjnB4WHyM6QId9XcEe4Y32LneUle0CBaCFfXXPd8nX9OB1PKzqJmlNXdYV6BaD3
d+e9+h5ps9WnT0Ptts4gMxuJweKbN1BXFxFs8CJ6vAK4NCxk1FRvNk7AZBA+Ktk2
Rz6af/IB5wLpRyT5lhWIJ+DCAU0Z/0fAFPRRAqcV2OA9iIaaLkxJAnTqDuqgkmpw
kAtZFg3xKoaJHLIc6odJgoahab/wIj8A10Fgaj2qqurwXT7SKgwiQVOLS6eARjkY
YpcjMg6qrQcSEZTYhWc7wAxyuUqhDKWaTboCCY6owtfFi05CztJy59+MK0mAR7OW
Q8wqXB7A1uKNPqVjTUgf4Y4mi++odS5usvOgoxZitFdgdqMeiOQJk80VlRqlVvQ/
Qvma6o2bc5YmTFlUSjxl2QbF6GzAymSYYahy+GZ/RqDDHIjritzkZohP7isdMwEU
QBoROxs8fHSaMtcyP6rbv/nyKd0PIQhiGwvT2UcCYFP0WzXtzAqhF6dlVpj/ttHU
3hUzT0PTXc7sDtmPJlabMskebsViUpMC/DbR/QFQ5z8PzRXOUtXiuw89f/IkDcAq
/AyrKhv6fGsgjEN67n9WzJ86ULA5As2hkw/oPzAWlHVykUkXlEWZ1wb1BIXJ4IzL
74Cb0HJmnFlCrwWcA5NrZ+cs7qbHNph2Xa27Rt1WYVKK5MsX/mQvj6g6yoUCS8HV
+6QwNsjDs5ByVRgXHZQQ/ny8JJD9tJ9CkuiWDQrR8MYAr1p/dQuAuuGc76HjkmQx
tIGseX67NEru57dOaoT5jtWQV7gxP/ClEqiDG+tj60ap6pjoVtofJ8/nlWkt8JDW
E/dFtAAThSDc1Hm4KSan9hd2CSeiIrJcoU7almFJnC12zhbWsLw6WCKR4AmYgHsA
+rnP35GpEoL7cAZUii05VbOzgYDTUzOJ6SO/pJxYYnaS98BvRXdBJpQibnA7oLLj
uSk81UcQ5URhOXD9Lj7QkR2sdSwaP5Jqoc9H1ET4+oklTxVkOduySvKenbNBvgYO
r8wtFDyA19bixuCGfj3UgqgH6XVPYubZQjvAs+8lN8oMn7oenrruVOW5ys/PhIvz
P2p+sNo4jR/p3EKyth4/2v0CFnpV/oxHfowJsnhH4tNpXDFUo/f7duklG8Dj+4Lq
EUn67T0PTA1Yu6hEkRrSvGOB0c0r1D1xw1U4zlFuiJl5d8KH6h0C8oXvVkluUtw6
bzmVh/vaVtKgKAPEI7f35WoVfuxgXT1Bl3pD/Tn3mhHqdcnpwsXkDHGDG9Z5fXm7
eqmsbPY+PBoWexER6V0XqYYTwV7/deYTTDGl9dG4MKHs6f0uSq91kW+087ObxJmi
158f0sZtw+1MmyxNFrRkhmWRIyUr7EPJn3tdicuWEJ8P681tansjZMf7jO6RM0oI
Op8sXwZTuZPkaBtjDde+nXSABTvN3oKHxSS81+0ieJfCbvI0woIxJvOj81+F+yNh
QUJzFsGVehDvk9T3b5dteh/s183A1mBl5GPyWHhMgPxZWUxsti1RfSjd4WWRYesD
5efyPq6S3Eqlt2VFa6Lk8VGv4VpN2ZJcpBkrlyv3g2Q12cvXxp48U0hKa8zcmgKr
C2kKM8ebdjzT8fqfqi4HM0TTsK6bB+Pn05gRtSO/nabFYViSvf3nR/2WXyZ3xhgN
9N5mcHVD+SRe37jKBxvVh/JHzIujgg56WTP2yiN8AiY5G6qvsb1Up9IUX2l6kLz6
6rXult7tmXDOaQ6Ezum0ZErtaIOn52hprZO6ziKrDEkIe1H8FfIUOFML2spzasUy
BPTbvSIMIMWiwb9nZmrP/dC7skNWVM6aGcxruCY/6o9H5FNH7Tce1QIXKrE2RnJi
PXRDSzUx4Ykh2MyozUu8INhj17oDKd0Qw8ka2j4mDDi4sD940NiL4dE4vlcXZgqC
hMF3rAaeKCMZjMnOwT4kjNOy8vEe04SUQAOr93tUOw1UTO5zzQ1TogPEsgP+oRqP
GCpIAOwtbWscrt/WR4m4DlevtbWmipnJZoTMzkG3eDL9+jN3p92d/seYgU3/i7uE
ec/LwMukUcz77qPTOpisJx7QzULOr57uoQHbKThvC1iO+bIYvVHVFogZsDykyI0X
XgXmOjJETuRthlRiQjdYtVbPnCyCii+v/y2jssDP8HhT4OpWEhTTd0lD53VMzVj7
fGRaoNPjqvIOPqmnXEsUASTKIeqC9vQzhkKPuInmS7k1O37Sae1ryp6+N4IZTmTL
XPJtojksIwOgPwT1Y47OXQwQB1HZQkEaPyZ9sC7Uth21dNypGxdrXIsO/FuJ+hAY
imHZGjh+ogkdIoYfXssnozupx0QkbMz65XOVqXdRtUb6ARVZEbkLL9Esw6ADWwDa
o2uF4D2CK2Gur2cu1hkVpC+rB/O0BXVF9Ox3mwfZE2GmlibCdFYTwmU7yddyOkWm
kBbajStzC102OsLCamadjY55cLXfAttUSeHFxdcfGs5645ye/8oiIhNnqD/drb8I
sitLumeodwTUp6Q72gsx/QzDly5DTLfE0jbBPW66eYgrd77B9pdY8nN7wWFyk8Nu
Ua0BRwTaZxRNh3pKDVmbI7WtpR+MQgJ6QqqddGUVxsPLWYy/9DS8aV/73zbyrHkl
7Up7mMpnduVRLL/Gf5AyP8zY+pIYqXnISb7L6y1xJEQIl1X0NqeV59XRTBptOCsM
vb2u3crde1SVSMitx6Hw/u9Tf9VBGxhL6/OU0nEhOv6s5RvwEfBFKhF7hmtWs9wn
2XoEyzYbo1DSZ72SXeEuJhCdvcgKHG8+Hymp/4Hqt1MVnxpZZn8s1OZf3QFLrtXj
neMDZyxbLtd51VTZQXc7hyfq8AtWEliLPfuTdPdtePH0Lmx4EjnNNR3BdVnKS8iK
kfRSzBAVeCKiU6QQIHwt+hlGsjcwC5KQWxxBlRPdDCuCj5mshr9FKQC0ebmWKqnN
t4Qgrryg4TbZD/V1/ErTEQtrIS69Muvtb/Ds2sYMaF8OXKhf7y2g3ZWzsu5r+u01
TnhLVtwNzjwoDaEAk716SVJcvKEHyKsZfIPxg5cySSRtET0PN46HfXSnV97k1i7N
giESHCwexpFvmrFNRzaf7nq2L6AoCRmWjhD7KBL2W+JTPkH9vWpbIXVb84LK9so5
G75vBQHFxfbkC5m96rSE2eMw6CXqWqTWKH/egEMkZNXdk8LoOH2G60JZSLGHdW4N
XU3HjCorLDwBzPhaExOcXeFyCtXrG/27+WaCGPvruF5WVTysTzB4iVK48af+PkDr
8Tz7OcC1DiI9N0Mlr3EVl0Q9bd2JhSutLEA3BosuY0P3IzsViNYnQD8IAwMVgEq1
ACyEShUfQ81FXS7/fEsJH1IyjwLn7TzCMHUlKSzBP+3ic5ZYE1/7bcB1gDGX3a0b
KfePuZGYaC+SwZsnnyslo/ostOwAY7G11hZqKdJ6TkU9Q/zEkZogGdpPSeXhKn3f
awflRxsEAGx+kZGYPbh+Xc+QSo4JinirBjSGDWqRgDeGADnkynD6fxqvf/SFSlxj
ZJgOb3pAwYqLB9MnJgoRmH71ut9/+oPXl9KpLJjM96MTNP4MxLwWz+ZNUZHBvrwh
MVsGIhVRE4uwCSavethWV5VAkd+S+VCkV5lK6xh5ZKCIQUMhEBLeo3i0R+97L7SW
dxkdDUgptyN241ry3BFZmTy95eVwWdiUdtv0WnCieM9nQubeanUOX408AA54VsSK
pphqqIUoIUdjIlZc1jOhGXSpeUoif3CG7Wi09DqVl3EYtwTGbfZM4mRbKYm3qP1D
2pNdPTXr4L6o+Y7KGcWN41UX0Nr6lNHdvJ/RBv15hHrH1gDkUZDjGvtY13+SXbdb
Q4NizC04ojojxLz2ELPnNUH6TjQuWEgsPZV8pV3bMJxn+aRU0NVaeLqiJGNb1iPA
4QhP6H4JLr1SLY2pd0jYMsWRjfZtctR3qmUJFMsRwAGCO3mhoEP8rx2MM5eVx3e3
NGAlBPsvWvofl59eSjqAzwpZiJiOkHnXl4083tncpw2S23w6dHb4H1JXYIX7SLPi
/8O9ed7faMD0SqwqlBTaqA4gKKplsWg69x4Taq7VxtChFblrmgtWHdxT6k4ltayo
j2/+YoJ0blQ/XBGN/lUpForJ6O/QCv6wPvBweZoSSPIWISv3luGnwM2TjH18QLtX
g7QCnJdghCiGiVn/b3bjNbZWn5qKAHRgDRq0U+moCisN54kO+BviEcFE0PXXLt2k
wFOXmgC2k7fYLGb5G29j0djqENfg3lG9BA5JoDsdKFxbek8x5lyx/6v3u09yB27p
Az2rjHhShPUKFoHcNGyewjsMhyVGJWQtzTl/UTpzEwRK64/HXDEAsyGDZ+oBk0Bf
4OKeHyVb+Z4rt/+XZD6hjohYq/XDPM2B6BuEF0VqhKPYTWyhJ1iU5HOVfVuaFThG
t/4h3n22u6F2XkAaVKAw/FzTTj7ChC6+A96rl1LoReSXtKnEw8eeQgvcFYRhm16z
kCoaOlEsjJeBWhQ6A/cEWxZiyx8jXpXa0ihYK2L4cAZCT90IdhJXhl6/hOIzUHrb
WZk9RF7DLeht1gcAfScoYtisvBD4LXxzCiUeZraiTL5XC44ZV0uPSG5JfeLXub3q
XW9lW9ne2kFkvwQfM7QsLSmSNzZbh8+SU61sgldidTeOyJ2fE1SvFpE1DETBiCYP
syO5q8g3S6QJZGzhKgZfqGMBzpXKdVs9n8T+Bu2HF0B1f8H7suEYdsBijdi4oVP/
K/JL+1WtR/L1Il3xcseJvg0FvBO95HijqdlYyOHPEFkkVF7HJkSMVdOYoNGdApm/
fFwur7i1e/Y8NCQwaR5Sv8vsbHlWlS/BHm2lxvcfbIUuhWJrcsWRR1G8mmbMFLLM
At1jdlJpFGJXz/o+3reu7FGbvIivoGwKbwjWcgA/zCExuewErgVSjywXpYwHh/Lc
TKq3lifrKFaCZTdMRqTEseZGzEu13CYE4kPTUokbFq1898ZRO+E9kAD18rb2PLcu
4JUMie5zCO4bLszxfHKY3bOQMY/VBiL06TGpAizyLe53J7nHdvrKV4P8ovRWgS5Z
hnyRZggBA3SIYZWJCmNBvAZw5EQ5RtJxhGRWiAAc5Y6KnD+uQtuVOvRc8J9a8B6V
X4dq3ESjKnFN03t1JkTPegCaKJl5hgiH0gLqWz1zMj9jumELlkwTeekyKr4Fh8ki
3ehpBdutdPVyAareIhu6kpE74UL4W7Pvt1tUr0a/JcMwUmbRSEPsj0MDlZLOPe0K
y8IrrDcRf4tB9E8pwMBvTr8YIAqcHUqKyjrX5gi4DfRcrMt9JhrunjZQi2/Cp2k6
QAj21ibE8UCcVVl7wHpbSr1c2Mje9esZUuYNsdcFidZZfhhH44XfJgmW2SEN5J1H
BZb4sAqUqN8KOXWbhxfXA5SSFzUh270lspMdRXtNIDClyK6A3CXPDWAfUgbYiPjF
YVL3jfv921pugH2+MTuY2vP74ficXCDATziWdBhHcaAxQJyKSy3PwCB2kEiPXT3x
SSZBRoX/TtQdkCc5uQmJOMQQvIDZ7p+xJDOOgNI4PhMmvnZSVykTXXRwR8vvU2l+
ZT1lNzgc9DEA9QwbbHuGL0WlFAODX8z6nLNLyN4up/UlASaTMt0zxfq/MET0UOW2
r5fjfRjfJSsceXYmVpO0s1w4eHWJYgZgt5vGC4A4eIBFVPDQrvHGVa12ISW8oUcw
FHY9m4/Ogh3hXOyOiqs+291aaXSMkmYLFZDs2+roF6Nd2C08sU33akel6BMQnA50
lkQeCBkaE3gtZY/oRFHJ4LWBIarn/SyyzpfOlvKoVkV/CAP3eaiZwcn6URd8nPPW
x1nMCOxLk/AQxDUjwff+7b6G+bK0W2Adzyms5xX68GHejG/HcXUuAaczYuirNPja
0suWbiA9TVzlNgVVzD9xb/DlvQlWyK1T59HggsDcUXFohLxyYPenTzPt0mLfhMaS
MPwjZzqJqnyHQ8G3OXSzKmidLfNKQtn5Lt2HsdbuEw0ec59Z8UoQDcIq4aXelNho
0qzR+/AaSZj4JOZS5PjBPVglKkPtnqKfOzP/J8YUtBvlWU7s4VF8FASUzKkeWlUM
A+zp+anX9VUsV52hTmaQfvB0roDW4Hr/lOn2KBouqz7ScRik4Lf7NuEf3By2zLVh
X6ZkcGUKlLPFT5gQMCalsCvuIcTuuMi8p2ufUsfc49HMJHREO1p0ELmRx+52f8CG
T9t0LCbgMq2Je1l9HifGwHxF7Zs2gPNyCfpYhJZ5tfEVSYMVXyBPniPdzshSOpIL
ClCwGoJRcziqs/ZZ/W4j5r/86UyG1aJpT6u0+XCHmM4q+QaJqKlR30ZkqD9UGwth
nDcnbNPlM4V4cL8LPJRKO3q0OFq8vi2PbOQ4HSQjyvhpQN4buDWYx4CUhj9FeHkx
liMSyxTY1/XRQp86UY85qvWN5i6YVcZOK0lzOGyVi6gRC0e26Zwz4dshOHBJAXXX
Ye+qNylOVBrBCg91I4OpNVDs2lCdn2JClu08FQRxKV35O8vLJy7ynE3mJlN+N29D
1Iy2ZQ7LU/jxeYgx/pnxZjQCB7OZmMMV0bf1+JiwZWXsKJ6WYhG8I6NqKmurJMJC
YBWDfU7d5b9/jer6lPixNrm90zSt3a/PZd9GDCbEq/DfJ/0yWmn/4DrBrqgOT7Oz
Nw9vvRV6GCtWdzVpawK+3PFK3l6rWjqF2ODQuBh3asjtIjpwX4W5SxRhRg305LB6
ogwExOhO26WV0qo1EO4gU8vv6LzIZlPFyyaM9ZcfvkFQzF2uTADh6Mw7nWpBo3jE
XdzfvaA9doLc6akLgWy+3kyvBqDI65WRpIqrpIKcgFJfaMY8rcl2hongoEMqJtHL
95H6AUzAT26GewaGH0pCnXJfrzLD42b6KBxUzDUbT0rQ8NcJpve3eYj6DTdLl68x
rzw9bPjN2TucBaXuDoTcM9C3KUHnJV0DZLrwPX83W19b3Fy/+ZAiMud2F4Gi/911
lyWwYuqhZt/TjddUD9VCXT1cjsJDaEBZ3Fe47wHiwFzGDhWPNR5jV3IODlCW1mMa
zJdT9aJUFF4tpBO5jxC4hHePfDgAvdCCUnj7IZqf2O7mBhLVnA9GMfHMC3Joig9F
DkAMcKc22zAGZoQzOtA3jLD7c0arE2640R6EoDpECRzw4IFz8mkMDSD/Y21s1xFC
2dmKOf3ZZUD6teQZSQ0n8RiX90Lt+8kY7YKYF9LmbypIowNvTcuhNIaBBStfRKnY
TG3amj9+jF0yEZ4MwhIbXjsW4BmSZx0MFG4jaO5FOYxMCT2AaYg3bYTmGPi9djru
e2QsEN2BDQfLMoY4EU0NfVk9+PdV2BAgikVkTMmIFVZYT8lyuT1T20ja8WtTEFMm
q6idWI5lFVtHk5L7jQuBdrih9CNjZy5uNS0E8eLy+PoHp4Yxg50itb6/tzWviqN2
k/4vT97DFmHzTjB4DKCCrrW3CNTGC890yKCpV5Eet2ZF4m3DllCUcwvx9G8KG7K1
aa9F94QLeaVlSx7tcWjOUGXrypZU53o00t/Jbos8NTejv+DiQZKUqiNJq4DDM3j0
UTc2qOc6Uy9AriLehRJBGJzvlj8uFMQyjxsrDtMwoZC/kRN6qY28JXVxBwPjqECp
pt4fDmQZwvwoB0VDcBtgeWNDtXO74O2zY5HTUSW9ZwXboiUCR1MvyRMdxkG5Sd0X
iIJlCKd5FJKX5nL3/91G2KyRW+M2/nIUOFFKtITaIGQ1f72dMBLgGNihzhKjBLqB
f5k0Y8vA6cHFWFXjPnszWgaQQvA3IBAypHQQIXz5QNHOg4ZUM6atJbRnySLm6o8P
YfDj74/PZF0iQT9uvGdBRpYWcOcnywTPQ8SKHpgRmFBFFMjqwPqgai9X3B58Gvv8
sIWwq7fWyfN+lnl3gwq/BklfkQ4eWEkw6QphG0I8n8HZM2epLEbYeKStPr7qJzVd
YEyxxkgTl2RDbJApUZSewihVvOHgxr6tIJR5kQS2XwMmsFA456ASnRrEZa7yvmW2
Vv3OczxzqWdr0HZWvY5zXxGnekBuwJ0c+nqGffP14BNDi54gytMqki/np6ys2i+L
2pzzCVMDQzVBnHa0lOJtV1Js9zxru3WSntm+r/v2rkJSEIHMHJYZSU62ogOqz67w
4HSxuJlRfQjtBHOYPJxhwls/0Jz78IbKJQlcsrlT/VCSXnDI2EpYD7LHzzD8JKd7
1j6fGimX/2I3qwQqQCFl+g7LrjW9i+254hGEfbbt60lOgCvWerfUk3utXS2DG8Lk
YaG8pVU4cMqP/fzv/mcAOAaVur0dU+iEMPMM9UcIBsPYEb4imP9tMWqgfYVHQgrC
CZBy+ktbAGeci6tmpJkdrp0WcOGS2ho3/0q/zpOV8FUg3qsJ0sjDqC6nfsVW4Ey4
jOyAHPoNSf9i/ERFMt3dLtZ11dqozfn+w9CQVLWrBMoK9nxgyJxeo//QJK7KF4Yj
3ONPyS2vb6lwRIl06mygNpkNK7i+QHk1O4ebJcRkysqFcxMZeFFWMgWH1SVyd0N2
/TOUAmVcjtpzkTX8Zq26Gk86yPeKYCFg5jY5hY7do2fKIqnobEYnVbtJqAkbvqHK
ySUqrf+aTNPQ+czaTYBICBz+EeVM40mCdNaMIr5ViBSnK9H76aNudcaFC8kxHFYY
+JsxWvm6QtCVRpWHaXng5rNH5owxi61YJW7HIyz2DYK736RkUfN58aKFc/jxotAr
qkikNI3D3bzkKmOkydPS3LNzN/CVpLDPzojdwaYNV/GEmc7PJEiwOw2z0SSCXAvK
IYxwFtfywuSKEjk+CzHT/tDT2AnChY/riZQa0K8Y9Z99GLsolDU1kUVHpiyfMk7B
46H5VEZJYH+W0k9pP40sjBh6AgBBY6iYs0xhFZHZcjqSger4InGGZdTEWKhH+Dkm
TksgSVmCVyTg8T0xewcNGw3VljwIX/UZsZr3vvKOErT4Ndtei56D0rXdDkgCzfl2
WXbrQZj3hKrXl2DfzfFB2pr8KFgcmMwf8mGyGyjzvZlwPjlmEphtoDjoQXyjtLUe
jAdTH3u5UsPqE+sz4lUXBsHOMwlG23eRKIEBtte97cLGb/eTSZW4ExbxPlZK30AF
/HPizr2pwbhASX/U/P7Ueegply7tuKs4c5TthvwHQeXUywrtCufAWCii4p/zqzMX
J+JuCIpIWCjyBqfi6+ieYD7YbKSyVQskUd5WtbYFjvYU3UlQpsugoeIrJJQX+XIO
+oHQ64CjkQUfJzPjmcs+3kw+cGfdM0vvQGPHeMpwPfwNuEe4D8mJcl2m1p5aGW5O
k8GxYLDCpPLIKze5+OjiTdD2NI6L3I1Lcwrqdc3oyLjBpTPBDu7jWlkQh5T1uoe3
9uSS63VMyytk0jPKarMQ+Zccz9Hl9TccEej/oo5npmOoO2YBTPlx8mMFSuCit7KL
0jrwuovcWXPXivlNmE69MOnMMqDZol2CKp/grwWySA7Eze6P6UaAmQgs8oU9G/KK
nfkpdZfKtP6dN6sM5JURfDCFYW06Bzb83ef5Uirn2Cn4w4fQaprKTEX9dQUDn9Dy
14QQGL3wnloQGIMnEQhqntGQN9lYr4uigDpeCea+2f80DhuHmmY3k8ks/0GT3jWh
q1IMT+Jwae/VmUpbcYQp3GuVhvR/otEEEvfqJ0lQKpjudPpPHi3dTWv/P4BLjoVQ
omKsQKGLwKCnPUddZPvtNdbNx5zWCmYJfN9F0D6bwYWsouf47O2ry8HxpypOQqDL
aHPHr2RlnnDTgKVad76Osbflgiij8rYwMj01YmDIu90zArj5mv9u1oayB3+xse5L
WC13YzDi7WOU1cAduG/hZS53NEYdjcxoTOIwWdti9yhwIXceFvzuHpsIkBu+pKbX
JILq35TWWQu/kosbZ8+ubooVYYZfPgDo0e5ZGyGk+j6wHs9ZccluZONA5RcSTHJX
xM8YOEIsUm7Hcvw9JGEGkVfQNTLumJXOPGsX2n/esA8jBkzXtdAuUVoYlqYuyl2g
b03zSTKVmrVmOg2kQrSRHyZB8kujKVFpsLMjBtKUQMaQRNyDWHFAeXbz9sjqKXcf
pKQ18HSeLc6vi/DIMqmCyhVAyVL6CSR0mjsb0BL/HvSqFGcVAk41qNDhvntWXny+
9QSz3xSPw8cuA0wFVStBn78SRsWwx79kU0mJAgH6enasTTJWhnNLnmywE1Q/gHRt
nJQmVCgAp1Mgy+DBQAfKKLV+gdtYm0OwaQ9wRJE7cY9ypsYy0iL6kdQhRCGa2utV
eh/EWvfaaIhCjlEj0GeHaaWDS0nhDjeG918mWPXz4oFOPm0vvbqKnW5NX1b75+JX
Yi/o0fBTcHlOcwBdkPbu7x2ccPMcnMPqTgT+OZQpHnhMvIrLKDLYO6qmtfjp+eK0
6ZVXA2S1ufEq3OwWuJkAk3/+26R6alyvIbLHhJTsUWLswyj2tmiDOkiCT2t2ZqFV
ZjlWxXz64CNtSJhKLoVavLfcBI9vB+8aW6lHnJo/pUc9g/dhaSNH0vXhnlxZDyOi
eP2UaxfV/4BTc90T4kdCSjv7j5w+XOEnfhpiNgHSXHPUN763Lg/ihDQNm8zzeE03
49oOZZcBZcsCHTYABYf79nPZvUZe7hNDFUpWCXpCFfu9Bj+6BnNY6dfxKzRGrbhz
do+Dow3kleMCO35T00m4sfBgZcEn5uWI+s7k+opNXui81aFiRxjSYIHekBOigoKa
dxtGlyPlQfAW8+PdZRE7ROX8pqL4bhh9rnXfu1LxhOPPTx55tOQbW8OkQ3orwg6Z
WbnnG7jrPghilPEnbwEt+6DyXa+tiwRmXCCe2MMn2Ky4gszYLyYkKvQkuIpvrDAI
4gdZwcpeynbG6NNzEbkCVkDjOCspZOtFvKP12GjeOzpNpA0F59CZAMJXNgVrm1nn
9p7HGNrSpzUsggd+Q8+dH0adMbh7Qa69Vtj2QCHF5lthCDXqCEXHuXdMI01I9oK3
h546NnqjbpXpxYEYA1dpQVc2G6jIPkhurMvr7UofEDGVz1PknfNSnF3pJ0DUxCpk
aoSX8xr5XXZvqzsxKF0f5ykmDHT/Yp6gOdcufJfYzkLhWS2n88h38diDEike7ZVc
tYg3KVReUqg2MWPHX3SqygkSM8+6v4ZgHOao1mUKSVD1K9TwIi7uXtzvjh6kuYoz
YWioacy02aiCgSvMY51hKuJRfofvQhy9l/BhzoH25CnrAzm1pF5BNpLSN+384YVk
btjysFgN7Y7LJIF8oXUwciM2jdoXVbL8jM4TIUVq7bFIGFH9Y2xMjaFI0vrGaL+P
4T3bmG26Kb0GeTYD8eyIUyVbwhL08qB3pLecPw6pug+L1aj5LAs25mK16TaFpe2v
dOd1LDFJ6RnZJ3r3wltqdQwYKoJqu6+UB/wATKET1JtZqMkISIeOV/yzJDTqC/yN
kKJovTlbG+ePmrNVBpQSFPbremAXwL6vUPGE28SePCjXP/FgHX6nBOna+Msg4bld
TL8ye8VWpfgGuFibzN02KrzefpOoxCMroEDshAhXgBFYt72CyL0GCxX+FZwd5Kne
2M76XTBVX/s+fsfkuUzwUp6PT1kDvxF5ta8JR6bHAuKc6x+jfHBB3IwC4DulGg3B
S1d/ZoxANSfT5K/8tOqZp/48XOtHoEq+/GZqKI33ZqiV7k3dJSVkss/tdObbnjSX
hz6A4jwVFN4YV3VlaT4LVWHN8HLqF4eHAhR39hXxY6VZG1ifn5mXpdRhEZw4vNAC
wDyHZXk5avFWMlFmI1hhSjIvMEsx7CdzMksB6Dd8tMHkMnL8SwN2VakkS32+WsR1
J4H0mC8ZQHajlo6G6P6hQ7liTyS//hVKij0jXUU0qTkJQ1Jfkkqli101dAVRh6+s
4cedSrbL8XNGauQLGcGIB1a2dM4aw3vZkLYQsCuBnBhBSz0EMffH18NHbWlfaunQ
dnht2C7uQeAPAzfUpv1jdon9lyMzvnb5wy+CDBbTVkI=
`protect end_protected