`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 7968 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/59UwEX+aE7FohaWu0/8IpTj7mav863zUNIsgIH2BWb
Abd9opeuBjbGF/waQMI2vMJTwD1ie1YueHc3nSNpEh4OXp8P5ybZFY89uyGz3ztU
W1EsuUnchJoQgbHZ/sLbgtGRgsrAFn+ZoIeGN1d6RAF2wAESJmYP8zw+p00RvjZ5
g/irlrcvR5923+bWtjXsf6RvTQYyKqhsc/P2+tWWj2OFuB0OmQS7KzLKS7nDfZeT
bKwg6JRonOdMvPWhCqK/8Mruoz3bARxsspynuniE7crIHyi6sRL5GfBBFPpv9UYA
9dP/ODKReWYfTDMfrMEFAj2xCmAa40+WkjO4lFNWJfQQ4VzTDnBZ5vx8VlVlzih8
MzGulUs0+uLKty4lFmLntjrGEI6eZ33sf4iMlyBsbn3arO0FWIbdtnIsd45W73xf
jHDctw+qwsoPtEkRpKBgAxWzx4TMqBRgRLcYQXZ+OiRkwXJp4y1XLTBRvIjv7DSC
tvt+tskqHPykhNjUhsXK92D9FAQuHS9je99ag1Fvooq5qX7n8JYae8QIkIG1XOMz
JDuA03r8dsJPw8IaPs+1QgRQV6nu5UAwUkwZa1peEGQpD8xo3+IF+R75wQTwv0GB
H1LorUnrRRFm19IoisFOaf2vpyzYYADF6A9FhpZ0rPf45LY31G1b6UTT+Vo+O05A
klC5BaQ8tuQiq46+shuqYmQS6XqksVLor1Izdao7UQ/wB4Vtbw1vV6h8J3jyrTOf
Fn02AcH1zZfiAWNRrVv6urQWmUM1EG9asnvrKCfu9JRgn39rNwwLCeOaCvgq+GoA
NPd4kKt0lMZcvg43PZV4fZ4LA7cHptoSW9zEFLUWuZUW3NpMgBdt8Ra4rBtrCRHR
YzWf3gVWaXNBuBe+cyxTYA5USkzp6beo4k6rr3VQR7XeVW7TIy4dC+2jblj10b9l
xOPC2Zy4DIcZOH0rZ2OYcPNAZN7oBu8YJ/85WTc3ET6C6YL4oLPGXxrmdIaflOL7
uqeT//EYtJGlBTnSVV8Qk04h9ZpsE8SmC+QW5AacZcz38uzff2BIaSxJOaeuJ1EA
HqnIFXbth6iZ97n7ObuIqeTVxTXcIer3Jg+7hcnmX163mMB5NJatocu10OD7q81H
5vRFzm0miG30C710Hs/YHq2g9xd7wvlctE3c7d/1x/MhqA9aY57rHNpk5IbhdFM/
9ZEuQk1+L7UEBaHyAJ6+FadmLhuvhYjRZzZeD+P3ILxBbcyBngfEjD2qYpco+DAU
yuvVwR5/XcPe86GmTSQ+8hXqCPQwhj2i1uiuTWDdlP1q27LKb5v8R/elmT9APxhQ
U08yAo/WWPmxSlgEiVBcdSp/1dQBnfdul1GHYN6AkBUVqMAfNuFAtTzeuJmbA72D
Mrafb9oAYhIt7YJx6gfFf0eWuubiY+bBiLu1EMuTWX20ZNHrWW5jEpLFmTW09MOA
sKW/Wscu5eDzysy6E4EHGH6Jo8NMKTeCdHoNS0hIRHiaOPRqFJmRCgOZIxj6JdnO
ccDtx+XH3IoMnqep0hFCI2cIvE0AlTbqkddupbBozT9rtoq/M/lC0xFS6VXWkqIo
v0hcR9o9s62FsdgxTuNXQ2vntxM2vIcOflVmrovePiokKjn8/xp6o8aApdLpgvtd
AvcNPnMkugQYonXzAspS/Wyzs+PJ7HsDnhL7B96inVCk5Xz+itU0iB3JZXtmHd29
WxPhgwBxwewM2+Gjbbx1T33Us5AJdqCkHYKb4zIMiNLDU5ixppNU9pB0TB7PuLfF
UPWc7iQZdL4nGEc//h2hChkD4h+UQw+EajH8upKlkE+3Xedek7U+5bWEAfljneMH
7lM3lZUWtLzACLYfbsdm6nOashTRL9t5EU/CvPTVpmM+ji0iyBnDMnzD/Qxbv3bZ
dcIrScKKK4y7r8Zzr5P1XsceqYNWCuUH8RCUZm/6ZrpnBTp5TegaNeu0ZtK6hO2U
WjpWImTrBxFZfZcwdeJX+VdmPWtsZy54Gde8KqRX9tIWP8uRawPIcD4WPqZ2vjsF
PePdrKo7Akr2V/SgEXWAZ4QMv3iNQpp49OhT2hHP6ymRBDZP8Ai54T7g063E0ay7
RKbLU+x7UQ/fHs2FeYVAFq3FV8/2K7V7tMBo/mCi8DhQ9CnYeAOUuyeVahm3/dCQ
/ybxMz3Xz6MPb7tfEoA4cRn8h1yb/lpq1KfcIugHSIPBdZb1aPPHzMJxyrOzfZ5W
LlWPDGt2r7OnkTFDvyhOHrBbpKJBNGjd10Zs2MT/TdCop2EHC+7dNHWQ0coY2iDr
4Z7vypjkaZCVaTJa5PgBR/gtSmOJicGdTr47TH2ZvETBQum6Ws9+C+4PL9xs0/mt
MDK1ch2rfZpNHjOY0oynZAHJyDYaplF6QSKR67igK7GNgf0NKGjakMBngLBPwPss
xe8VUAnqxKUzeUsJLq2QL3E7Ko/8zaKohPp2gWcFuQa+4qjEJPou5EFKwpOfdrUJ
dh4ir/32uorXQn99MVsKq+tbylbcYAh+vQJWVoJS1U4Xm8raBxOKbdTVRFuSgvKw
7cloYZVjdjS+rXD9FGTyAqv7mKEevDCZa1DnG6o+15zLrIZIWaWX+Fz2wB6S5Z7y
BPP/m00gQ8Bt+uMUHJ8TM8AL5mGPrOqBSBpmIbLnbJzIBvFlmKsX+ElgT0TNCNGb
x8ZSYPLKlFVTrj9GM8OghBHW6iU1AZOsJQaCQ3DTMO7fyu4YUyTFqfQdz5VnN3V2
LBi6UhLB0IBYsU8CdN7Gi6Vdf01SVrp2Wpu7Au6gHtRBORgXOcfYDAidcfi/wfJm
FuSADaddUZZFME+dauORy2W96xykIhmIhwjIAMvXmM9YUteVyfHlbrOwA2j1IWwU
qWmciKMi/Fq4Zp3h3+ivHq0gfUIGU5xOoFWbyP71ECm/aU1tXwlcnZANmuyg1oWv
aNQfaEo8991helTSLa7/GMuLam3rEPkGXTn/qNsN0fmxqrzWQyc2MF/9rPvoB1p3
n9S618f4aaT7QGyGxbOWqm5OuQxPB3knwifrzWmleVzFz3QGFgsd3Z4x+hw9YEhF
O5q/Zu5jY+q9VldwdDTWtdZT+KKn0x9lTuZoEdN9/DhktRsAw/VL2hXPLp8yObxn
mBsVtXozH5hokJ63BftLscWUXuzBCKwsc6l1uYQ6EU0X6WoHoFDKUNzuqP9YroPl
+rxqC+rgACCCtAbliolzXTLqXYdr5WGcSwnF+u7j02u89op98KKjwTIElObHc2Vl
JjpA6VA6GFM2fnVDB5nNKUFPuA7V672ZtM0VrDnbKxTnxdmqI46kE+CKY8LFPS1D
qYvwzxfzCzHp7UfloOVykueqK0Dd6FjAOMhcwYNTs9K2MkQTOF5BlYf5at4MCXdj
jz3W8j34/pTaDEd/dBkgr6iq+VWOpkTSb1zlxW5nscaCizZYkS2cYDZ+XRaj7b2q
hBo14OlH5uUOdtERrkgvOPatdOEkd1X+4Js6/TY16FdUR6jdRXtY/tr3SNF1QSXA
XeVPA9uin/66Q5cYITrBZ9bzeQ4rUTdIRw27cllVrSEroEXcFkcmcxci83pjtJZm
M9WRFzg+p7pv4ShWsRUrqQxVGoQGiohwGF+tSSaTF2c/Xf+C7XktlRmt15sO/u/d
pFwLwbmPuMP9XVA+ZFh5K8TrYck08qRN1lhmqWRLd6qs/3TzxhYuIgtCwJio1czk
hc/73L1PKM/Pk4zv0Ok8p2bsXYxxfIlh7fGECCiJcALkJQPHmnBVFgT4ExSKELE6
lmB9HV0EhFpa+LiUNLsMKjBM/y2i23W/QEw5/Pi4YTOwdWoAc124PPUtvLj9BcjV
NTJkCqryf8lPf4zj3aWjjTj51gLNvNgdA0mIkG5ap4TeNSlTIdsHzB/A0+h7LukQ
ONlL4MSNcBMMkarZW/CID5NsG4lAhwB3pFghmG96jIi9chk/cSfEYmFjiB0GpYui
QaBkvIJdpil4TGaaxYlY6E5PzRWnqfKZ/oE10+X7ZDMDFI4UsaSbtWvdkI0DlGew
UW7/M7zPuJGPGGimLxVMAxBYff4l6u9P7Ge9u16KXkmeGosH7MmA3QCVtQy3cGMS
idpgSH3wjBcF0YZmkoSVghrvrRO6JXF63xop6u4T+FV5C63Cx67x1dn7F/L96Cu7
g4i+UTLJIOvIx645xVodCeOflD4eKFxKXSAqAmp9s9UJrFdeKx+bFt8BX3oi3qpq
aHK61NOL3SycwzyQX2+YrEFJQ5l3vkuZp8SHnomdoH1SmqD47Eox59mgwme0xikw
mrlRjaxQadhZBAx3+qnbiPxMurced83oivPKe0awSKGA5z40FXXy25ufs529zGlP
rJE9d1gnSdEljaYDRzbg4o2dzJo9IT06hDBmS1yAT6KHWnhxEIEJFE+F7Z8vWWF4
KVARyNLjDBSrQPtKUgxu937ORZBzvlStgKCyY+qzT46dxKh0UpOND2c5g3zNtPdZ
Czu/JYl26sbkQ3Dtp3gIWhDNYmYC36xsw9STU2kniOn++TK3ukcwC7j4e9xGKteq
6L2GV4K38WLKQTKY5dYDrlHmkvhNstrBVs+o6EFn28dZvsWo0ZnEUHLwERdrEJg7
LkjzQMRmKwg6QG0c13RRGvaKt21moW/8pST+jE8Hjdh5YDDk9sFvz9PV46gKVZVP
HpbsOaSO8oAlKQpEdJ8ez2MldNPS8JeYS0ByjAQ1JOoEw/6SzZQ0hORIDymxqJqk
RDjOhmqVU7N9S7mKECWkHEFQ24G3MiJBvWDxoit4rfGogKuNL//IrkDOObkWBCpH
QlFCMl3cCofzwTLrcOmYpI9gxhwPlvJWAUJhiXMiVjDIkEpCosNYBcW64EvG5Mpf
WKCaXGDYbEf3+D8o8FK3m4Ra67NtVnFOEBaAScLJl0R/zBku5wPMQD7JKG5Jmb2m
DTy6fk2dvGvolwriVpsh5y5EFR/c80e60kI60HBOYAKGHUBnXbKSKJVHgt9+GkJI
lqG9MJhZqiotxKNvbP39AcU9bsnunhJ/hvB6JgR40JAOBobMePSYb7gh5v+YLX3g
O5BAD+YDE/8oa7Y8g9cZ71G9Dm66loBSu4iGaP4s0OYz7lfz0VOO2uNp5fAfy746
U1ceseDjVGkrGthqfWivWkAKcXQX9SjG7/PMiWMECeEouqr4Ij/aQcSoUotjGbdS
v8N8PgSdFeEXzCDJQbD+nSO6WDr/DGLZsPzhxoPB9fEcEokSj6UDQbH7rYODchx2
iYl1zYEEEGHlE1Zuw7RM0SAYguGp6pjADuCs577oop9/gPy5ynSZ8SixEVCQl1Md
Fpw47w5hTn8cZdOQMYocdOvGkrV9uizqVexU74/4ELZnb28yYJME1NQSEPHIS5iq
N01l1ioKL8+/u8JESYmSWj16D/vvhptY3E5nfQKWsxCojNWuOINmsFCdr8DLghuA
8BLg1SzKkWNF1ayS8nShlLHSvYfnh9QyRWMRhXlfhA8vlAtNRAKYzh3pmOCnJlRD
y82NQdU86U+Y2IhBSPhhvik6dOnM+Sl6uGGudIs/DonERJgEeJ5qltJwdbjj5a8R
gW5SVZMkpj+2lq/6BZh0mTOWKjj3pMIMYl1PKq85p6nzwmglo0uG0Jl9IEtY9GX7
VA1HICl4hE0k9nSGLyzMUqoL5OG3Ia45FViVSkdykma9T8jv2PiX6pjwPFG0Ssaq
xq8W/YyJbKlDOiEGjXAasEjRI9etuAgCGUWPWeEjb5Iv9ILAK4v1PbSPYgu+LYjG
Vk3ehUA8mrtvgwSTJRQuHYneo3s0NM3NYNVqv4MLG9Tq8UkuxzA5sLNIShSpPwvK
okVi9iX9JD/teU5CXIO03Xl5TLD0LsjZOhH7IRSa3MW3Gt1dp3crrcqRd07Wlu9/
vSrQHlUCcrpFo9ptzBkE6yJajhD3laKgP5u7okbQ25EnV7Xct8D92HM2OF+Sk2Tf
gC6TdvkJCs7kPiLxI6c4DDDrwCuJ9NwjwbppqCrXGYmvnT1eLJnIV/KxaQ66WZ6W
3WhqhQB9GOcuSu7Tczqfa2kdwbJDABkMWwbw2zgmkY4AwrjuNRqTRE5uh4gqu1CY
WnuVj5+yEqGP6XpwN21r3Y6iazY76cCyb+oxFl/99Q6GCdauHzXE0DUIm6vF5mdv
Fi40G7V6hUmBhdyq6uTBOmqP8K4DbNLZeQKsG7ytjslipC7+jOLrI1lbAnquo6dZ
/YsxFs3VXUdF4tCeszihPSP6C5hV1VUW0mio3eh7q1v9meAnSQ3zeD1wah9GY9/0
7ZPRRD+J6fgImSlGzWC3Zkk0vn3h+UJUKvCAu4LSWF2LUYxRmOS2UBM/4/v9dTaV
kwRWC6y0oq/0c35Z7lgCpWLDyrDTrCpOB5bhiRCkyDpRAfoUY9WoanPAWInI8gXw
lfvwQaIaCM56T3QV52I1lsgTQ5cdx5zy2iysh0duL2Ae3EvHFf78XTVrjV43ybWR
jjoo8UrW63iggK6YIKxhZ7vuBRbLq/CryncpeJgEBkrq1zYetp5wwtyX7psBg/X7
2BytRsLCp5e07KjvV1hmuCpCfUIR0/h3psd4PSS0vJari3DfyYJUlAF+YDhAjzMS
1c0LZvaMyhniPU2ZWD0Pgu+7NLa4/HZ+2oEsoa6shnZ9P6l0LVOGx1KkeaHI+wvV
mYifN+wjCMYuhumfR3P3p6uigV66RoTTwaGcLbD0/HAsiaABa9M+pF+0yY+4dQYt
pA9X+wDVgaC+O2JGDXozGAVNOGWFcwxKYHdmwks6dS0jMJw/jUtDyoWfPoodanz9
lIrhTT8XRmWncHd9RNd8hM1saoUxab6gJg8IUQXLrmgVOMNNZqEdB8bRTF21qySI
/7Z2MFChL3lPPKTjCD2UMz1/KFpFimDBABNIhwBCQsHGVuqoieW142nM5UbL8aGQ
aRDwkl8tsKNFOwBFJlfKXor3LWh6nJG8ZAdAUnhe5iqeOTvrfCM4pnqg0ZRp6YWt
gW0klxVlZvcNPuEdnkOl0q3/fkK0oTvNLnGe3PxP8Q3fwsW5FPiw9nLp2WxPFvmd
CYPFAW0iaYZYq+feYbDL/eMcfgZtW5B3fxfv8DKEohQRrDOTA3OxY66c6d9mcsVr
zmfiNwibg3mei6iB0kL1FWMnC+BtjcbL4EbjJs7BmrPdVei/qSdJt59j3PXBC7wx
JQG8GgvuhEWbamGoVUkIcRibAbv759rTjCFyo1ArNJbkeNDQQO0KYeSS6TYpnNrb
w789643KyDIlejW9ZYnfR5kKlKQJHMgtC5Z+VewWeLjGSfEcEkjESiGlfI5zbMvJ
EWPU5ozqU6PjJ7nDL1fpZEv8p13oo0LGjdUB1dJK//mJ5db8rOr2b8IxhOwn4/op
yMEvcXnQv//awA1T3lKrHld7Qm2+lDYj6+3oM2WnghNBNtFzeeSFZ3DSbCWye0H7
S0Te2D5GBj9gBWTnrVeCUBzq02Fqt8KZHwnPf/+WllyKNbDHqXkPojtlX8UE+ztZ
pMjQuyyWjEmP/F7YrLzeTGaa75mWcQhwuTgb51hz1oZS399Um4HWqBNY8IRPm2j+
9pCPbkd7oneucRiB5NcYH8C07i7XVY2nVeHbdkJlABaMdqT4PHPyUhpwgIT7MTTr
SAunc5QuO9wW0ogswfcmopw8fUy8AE0l0l07ULjK9BJNkuI71EU9FKTVr8c5NKPA
9KFrgzLNdAO8Ew/CizhfOjXWtcVu3jtM6b7hwrTPJGZ1qv140UBdHGvJHEENb9Mr
sFG2jHvde9elUuOsOB5xsjO7YeMZbkOwW7Qlp5VqAWw6jUAHqMKzDRRjiUMySB3U
hOTaqch7g+XCxgs4OY4sqvEr4IWJjAtyo794ULNbIZO8Ysx3h72Qz7eM3Hqbx+So
VJ8hmZb7eSg10tLUOjbYZ12aJ5pJAT84DkMU5n3YOzdrV5eJ4kVt+hsfz5V0meBk
VXTcWIgqaOWajbAdEJQWXo4eQ4eEsuNZuE/XBXYeNeVyxI5HXhZfXIOUzq/n7p7n
KXcd4EjTqOVeg1WqywmLhpBoWAqlKc/juhJvjCtoNGVWmQhn2ImjQ5W8zQHO7p3h
Se90MmashmRYUaHNpr86raS4PJZ6i2IsLDAaW/8ems03ruye+r6N7lVvKu0q36zn
lMIyhg99/04ttc4BR5wZdAYrfhPH3IvEA9AyhT96DalL6KfSbFlJbZYZO9K5mMYc
hKPoeAKEIWAcg4GdSCpCCW2aApuk1S3VwhIPjXNDUU8Geipa8v8+BvFPgUqhqRcR
l6grOJtataQH20VJmt4rE+VP6ewInwGcFYdTTpaBXQyIdPmlMG2vJ9BbK0/kn3vg
qT/fiv48iizDbuEKIzCa8XbdQPX27MNmmGchN4Cx7Tijm0q+6i3i5ElpEo1JUlYH
YTI0EqLv5BBgb7uGfxALWeX59Fl2autW5qr/vsnAeNIHu1ZkJnz47qqs/dSu058d
Woh783eZBt0uXuspNBVHDHyLclMbh7Y6W3SKYm8FHCeWOhElw4YXsyRRv+Yaes/r
EplsLFSDzs3kiusQa8UKsEEIwut3+6Iku3ZMsot30sLA+Fu5lmpz+nsv+C5q1nnJ
ikfmWPyh8jkGYvUZMmTgp4SARzPeSkDj5OR/fywg9tfEwtbzGq5otE7aHp54ju5g
TXw3M8+8vwuDx8cNe1o+GMtqlezBlQsa8a1PF15B0DXFp2bnWIph7wOQ8dypKXOf
AitSKeMghmHlA2qa/H3POiwp0/UhzaYcm6AeG1vjqaq72Vd76wDYJXxjGd+g2wFM
t6th73ZfoMWyhMC1KsE37FrymeaNju4BtUobB/4hOCxIf/n0zFrTZLXJigq5biC/
MWREV0vrcHkIuZ2RPSfMjau3wAGDnDX+MPGZWbZj/06f8ZFyE81rSks6HUHxycST
F4dUuN2g//h1qd5S4Pn6DlW5fz+dTIcLsztX65Tp8atFJnzJspc19EdvmRYBJUxO
VaA35pzZ16PuiNwFmMeKkCdK+FLvzCA3ENQohN3SK0BHZTnF421WXoGfNa+3I5ZO
VKFGz4lenNPE5dVI/B8VPfT0Rd6smQxBODxyCsAnGa717n2psWOY2IE5hbVbuZdu
woQBb6eYc6e2fS7XenMWFC8cT/cwYgfS9cKy70VHGKIETv4PDUVEsKly07LSTVHe
6gzGzzF0EFJja117Uq1STgpfgIU1mpFB/Duvh/Q6pQByy+rTciToAVRzItkcN2It
Uyg8KRyCuSgXUiz/XiQIViOHymnavELtj8m9VORtL8SUnHskXsVKOCffeeLQ6QoN
p35Y/MZ6WvhNCo7wcs7Qkcr8TL9PXgWfsLN0S6wUpfiAu9Ay6x4hXYmy8hBFDH/0
RixWtKqEpB0jPDgWHv/4jb+CsfotaTMqjaHPxtXfCCFUnlFkZf7iBJvHhkEL2e+q
Hz/VcYMlSGMMTUKYhU06ox9vH0w74brLe6gQmpdFIDnVKtXm8HzDnS75rwanNmtT
RMakWPhXzBEVvvbxiypeGQFvR7VvIYvtE+IG5NYg8K9QAZIpBYYJ7FIyR0NllPK/
qEbQvKik6TLdWPhdrhCFf+PsuKvWrB65ADPRU8fPb+M7tAf96YcumG+exmZWAdri
wJiq9bxQbxjxKla21+awV+B5wBbuqZuFtIWEM2KR9OG+C7TibHJn56la6b4abXjT
Kzq3ifBhfguv+VM6QznuWzJZYvDkQNfJgJ0S0lQ70sBXP5bvogVLY9bnEXM56OgS
Bhp7mAkZ3mP3ppq+WYfvuIBENjnmVmdZtUx3ZaxKFjP/D0lJ0hSr62nskHRhTDJW
e5OtEmubHo42pD+lju4aO5No9nDvEomqHKwZXFimrU5WfqGd27vs5Q9hvYD7XtJG
iy0ZCChNxmt5E4qyqIvD2pWRtz2hgSqmZ9UqVnXGwlSt5EiFN25+6W6YZY2/pJsk
+ajrl8avtAxxQKu1/ih96W1sj6Si18Wf3QW/MIzE1YMjFKaKaFk89G6J7S8z4qdZ
PnE6i2ERj8X8WFOpcvO1npungXROS0iY15bd/XRmEoMitpfyUItgnv0ZpoBUWHQf
/2QR8FOm7j3jX+RlQnB7le/r8HYrr9YVbzCTPjbAKwHpWn9Jh2gKmiq6t6BnnvZB
v00k+2+VflQocfjA3faJIDSpC+NEngF3wTMY0nlR7H4eyp3nQ41VcGRf1zWIzzhn
ZUFuE36DtdBt71Y+D7TPPpbRZbAsduPsKegJcMlAj9gOprHUYqKvGuh9ieUppjlp
9mtNTJTXFPnAupgoMHrKj2WLfaoSu4CF2au25y0qdQh0Oh4PBgXvJC3nQDgc+XUm
FeUKoQ3qr9vf2RvJH764TRsv/DAfVGL779SmfySot3fD25czFvx37p8BDNvgUN/p
pu+lykUIzPba1Hb50gXAJvWG2O+isC5e9Vcb2HSvo16dG7EgBSruWLWPgaExq+6H
mvMYDEYi6ONTfm6I0O0/zbCCn5nNLyNIYsITBmc0Bx6bfQlEs6ft9ZPWcEJ+5CfA
V7JlZRKKxT0KaAGRjrHgukOC7aM+q846+Rr1W4vV+bwRAfVBAzGz04JQl+Q98AHJ
zNRWnJpQx2iUKdp5+LmQ9ZAk9feyv1Pi4VdqlTzTvTV6KueyeyvHL1YGhOGnn7HR
`protect end_protected