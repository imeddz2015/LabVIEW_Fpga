`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 2896 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/9huKRhRMtvnNqb3Z+UU7TahEoHV+T8U3P3ufru7l1O
3DlgtZzb9QxCbOjthp9+wDkjygH0eUfDrEl1ovhZG62230OIN9JS2cj2BcoIjFfk
PVytt4KqwGZo6TLDNyYlht+nBHyQvdGf4XHiO/pNpDUv+4PL0QHlhnO24GuzamV9
m8n+/s/vjCMZR5qfUNj6MkP2BsxHmvV9EhOU2c8IEXMLWm7w8zImiUJi/gONmHE1
r6fcelkh/9IJ5Ndm9dpcN6emc11xG9O9I5r2oMPZrIoX4SPPPPt5oxI3FQTQFQdf
7mt9/WXaBF1u9JqaFkTBtbHLMrdx6rvjLZMBJ5jumN9oXG8LAsASYkkmEjFXs2qA
SGsnenaf87e0BhlLhB1OZslnH1Nd78DbWL8YcCYgwHi2N1vkcHXkJjzSwWTDZOFn
svDj5cNFJ5ho3Jhm+K0M3eoKfZh192lzJNDtnt/HRzAUDhQZmAaGIuTXUrBMSwYZ
ct5S2IkBrF4jGQVYPb6tG4Rlegqbe+NKG0+biPg0+OS/yv2LWpbwjxvYCIOu7ujy
bYAyx0DjZntkX0P2Cg9FG5KIxVb4g67b8QlStOMU4aNzUNVbN9MNLJg2rN+m5Ldv
ET2ekHwjZ2Fyq0WDHNU9arNjhcarSmbr0ksZ0ieGDgkqhZEgBNQ7auwu8lYY9ixF
5I95jFjFI9hSlsyq/xuiXRKIJ+YpqNArm3npxKbeWHzG54BQtJhxKKywlDVwIjOs
wLPUN9dZeiA8BYqTCeWeUFgB3LNa/Cf377sVBEUxJ5vmljjlS35bVf0ar3AElQRa
w0Bmp4fN3dgEa6oXXUNsuA8OogOwvq8jGBpGIdPZZF16OUzickD3e3l9Gh4Y+4gy
sgy2p20p6WSLGtKda2bfxMZkxsNsm30N1t6CnUtfEtXHkNSXFnZ74LEsuFpmqwiZ
s9kaOAz6v4fWvuKkVE572k8paCpIDFM0cXQqhqJrVpFCVL+tK0weIia0t8ejDWp5
KFQPYbaCQDQMlEnlnOfkXWBIFWVJgGhGxC7KzBUiY2Maj02C9bT/1qOcFpQf7Kty
yL5m2pNHwFyHu+orAqZousJtksLlW6FC3pB2kqQy6/zePkeYbuFqYC4B4L/WY/b0
yn722SwSZLrQVspEaqRU6QosPtbdvAGeP8o9J5TPx56mMJatI0CnjX8iDXUKkpU2
e+v03VeFu1ZVELVRzxtW4I7+ZYoa+zPHsovxfYCHJ6DoPHREPxMFveIbdq0SUuwr
aLnTKDIE7RPZflqRkT7lZY6Xnhuc4Oj+DSacdHdTHBtAsaCpz/A2y9W0x+9hwVnG
OPoCb2GRPrK4CrpiZYl4pNOlpvXvrtiYlyEn3jKF2DmRMcLMQUvLh7sWaeWd5XXS
QMD1/7S7NXRCMTqGMT6dJ8ViYKMNbmu14vVesy93gKSwmJUc++YKULEpMotXvJDb
bpF/84VDe47ubyIMQHHg7MtKDSk6XwgaREFr3gc0cN+YDeLuTrg6Tqc6tJgsf06B
DsLzNIU7pzztlflCp3qISOMLpAS3Kq0KckG/pUyF8hMFy7ysd7C4namFoOc/ct+6
3u9ALLqXlvkZHzYPEoFVQpddFAjCoUbowgAeMJT3fUbniwF6Dn2zufAgzcoYFM2t
1gRaPTtc0CzyxxA3holS8aPHZTvdKPF1M6JC3Tf5DE3+ZrzypJ2qLGH3DcQigFc2
+kXloJYMKhcZgu8GU3lCLRajEe2pDqB99v1eFh4Lo3B0XSden/lMZKkHnyxHwsSd
cLaHDySQLB5hs0fmjCBePHPKsm63dweDVSSQ0L5IDk01YNh1IGD9NG93D+TjL2ta
VSYq9TbYqKkttHysxWnMCrHpzCSMVcRFII8rcMDlFIIPn7xGJtfds53X/CH85Byt
WtynRLNbVoKVTTkSCBQXH+21up28lFP0EYThrp5/WQrfz5wauBH5dRMOMrpVpI4w
Ap+U5C27RE6cRdqtvvurM39gL/HmrtEAUUGCrcml4If8iBPUhgahGMmusrYYdFrC
TVSXm87Dy4QihONBt9pNT07/+pziEifN+Zewyes3UHZQvRkqqyjvoKO+6jC8mnAl
7nEQOzk6qFER0EQ1Rxa8kR0o/6XCV36ib/qFSrLwbvmPSv9PwqNcQ7DFmNMqkDFN
FmLk43KXV9JiNSF3bneTXsdI5iGMJD8DKpjiUpXB1dVZfrGdp0C2RJb5I5ijcU+f
GqxeLBo97t0rI9IwaAQNKtzdgkR4BI7epvG0nauxLWw7J5V4fX0NYp1YTPXka7DN
kY5zV1L15yZIdQXBfD/+37wp4bsp4pFU8KQdANaJJFkvsvOoajJhNmOUpP3/7kUJ
RJsZTcNhTXlipn23A+nuQOpXqT9qXi9Pwl2/peEU8bXXBZ6+kVFZosXzPy+Htafq
4nojwZ+1wak9zvC7D58GCQdaGMLptihAuusdq23BRg8Ku0wVlkea8NAGtvskbSUP
KDrWuhbur7tki7J5+LJzl1BVSQF6zr5jQix/5sCLVB2vrCjjArP1oJmtmG9bq4Jl
5/OZeBrDHEEexLmD0fZ74JNlxSpInMcra9LxIbImrPAc0FVFvUYbZgLjyxxfTKpH
ngLhjQQCyAxb0Qae7IWV+jK10y6B2NqIHO/fnUpNaHNkz6O2BKN3bVdxXJueVEp1
MoDJQstE+sB6Bu2b+bareSjwIWItNEZEvOn8Hcgki0slocY+aC26+qNgkvQB96zg
6aCB17TKjjq9CHsU/xuTDDvjZr+ISawc1LaAP0yMwiLeAG5c0nfm1lWHFelPgzYq
pVt14uf6TqCRJs6QnuQJ4i+PVM+Ur04LFN2ZGL5X+i4uXJkUADMmaLRyjFstorDN
kG/gvS6hxdlrsvNsx4ftgycIb8qSP/ScZU4Fy3F+vRyNrYN3pGVBwwpbI0XhzCTC
liMDGp06UwK0MYSPnYgSivJe8keywdaMggKjCtfcsw4VRZ1/WxQzxFye10cOOpMc
ULKzSaW6aXrDL1VlN9/El6tk5NI5vPNGj9eCWdtDZQFfQMNV6usgXLtWvPnlIV7f
95oO/+Zd2rHKYg4o+RKxGHc2iaNFMhkHPa/g7VJNgnRX7FxvQqsQXpxlOvmw2aoA
eARBPuK+8lFRe8B6+d3j8DFPXZeRL/CkQBV/9W6TWhHF2dn4A7q1VVYrQIrb7xsw
YWPcDKQ24UsF4aJndzX7m3hK/1uY1x3D+vjXz4gkMYGBNlWkzXo39k8fSvUzjtto
PHSPG8H2tsCXLDzfmcldbWTw+Umh1Y/3bX5OFkJtYFClQsYJLQUG361XS9RSiS4m
m/JKWIo2+qe0LCBNi/4nnx9j3MQROBNJ9HBlzm79rE3AWKvi4oc3oGe/wgkbz4VX
WsuPBDGU8ZOIhemh0LsBQZL1zkGroK6aqRlZ8VmgwXGViISGLIMcxOBX20a97hNN
PUszFIDxxxCE1PLP6DnOOcHRsE0KW0ZFez1Y0lVYw9YZjy5c9I5t9N5xMkSkS6Kr
nKtH72EE0rtZXkf4paRyBjveSRP/uY5eBzFB0ot/Mmr3mrDPyZk/pPNu5tc1Qpro
hFTJJNIe24NeXo/N62P/B/kmN8sORweZ8lw/QuWg2p4xzRWlqxfdrUsBdfCHbMIv
iWHo3OqeCyLl92M+fSay/snrXityzex5RF/CrzteUklhDME3k+bMeQ8SPyLlcVMi
lfm4wlceWI6tYlW8hxDRGHyXmytNyAkekM/wUvpr7NTRBUGKKL6/sxF9SrKqJqhS
6PeOd3Ovug3shylCYGbnzJsdthLdxCZTu+DkajUa5WO3jy8Q28LKhOZBypZbgK0T
xNRDLwsdKOWB4blwFH2KlQ==
`protect end_protected