`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 45568 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/9huKRhRMtvnNqb3Z+UU7TahEoHV+T8U3P3ufru7l1O
3DlgtZzb9QxCbOjthp9+wDkjygH0eUfDrEl1ovhZG63HSud+dch267pl+0WTUzhj
jS/LM8GCCvZIbBczAEJS/HWaOVGBtR+IsznRHY0KUwANbQeMKsDPgushE4h1JxH8
8U/vKIpnfupZ7hjeVG4avBIrohx5ODeBUoOrHoqf8NhA9NgAxN05Z3Q9QX7gQ7uW
DUoCrJMYvTMt0YkqEiz1P0/s828rEQkZ23LkTWH+257PBlWfRSq7ryLeUViPF+pz
lc86qkt0wvDfuW5W0/v4qvQFr8SiP1ekjQyEVsACQc6BFGOUbzSdpMepOSPNjnsV
rZz9cqS11dvNp8hLKv9tiesyghwuGx/mkxxceS2h61m1PFQuRwrxlhlT8cC8Qg2R
29paM6g+AI6jH48Gm7c//aPc6pPwZaD7zSJ3brVrj6vxuu+uGXgCdyknB91AaAqB
ZzkQ2KqNfgg3oXYXV7bMi11m5wSNDJ/BwDvrVOTyeGjuC+eWitv3OrrL9GfQb2/r
XaReVWHa6U2yMEcn31p6Kc5TDY+xuAio/AzhYCyjdECqyT/ANsyTE1LvchnXcyfF
De5uYgT54cBgsnjVNyJ2vNbgWW5Bdo8LsiSvy9VR/Syg9kojZzMcO3Btx51f8dOo
Vae7ZDBdwaBSdsK5ahpMfbxWFYowadbfZjek7MAA/+NjOP4dP0Bh5ZK8WtKIRc8b
C+wiEJJfYGF2M6AEG0n8YqwyaXCzNwW2LAvkG3Ucr7Me+ZgsBLKw8r91IznUH4z/
EyzSaz1G8WCFgSubbHRR0CXwJIZVeHAf+nKpMi45sIke92rhqqQA1Z0VxzP5/ORo
m84tvdHVG4aI5mSED/yri048TrSYneMnzqCoW4U3Q0iCstupG7/DR0WWkczHleFT
unM4OWIjlRlTT+y1dl4yIhXg9XozBwr+Ye7a7bL7/D5Z+7u8dUdNBpw8HmJVhVCL
A0UoLbBgevQBB6QcazkiRG1fr6wTMOz0HMNyhOCvzMRqYMlYwzCw1pe4K093pZcl
QQe5tA6hM4hIsZPED+Z/bK5hhvnQlHxBeaz66p/yCo5jV9a1nm4/Hg1R7F8pTop+
UvI5XAxbfR4IcZxj5it1x5lSyb5AL0paEgiF3+WJgqYevh7N36iMXfmTrco7A7xg
FeK+1JW3Il487zGc6tJuDCmebO9YUYsgcFL/sqqJ1tpmZ3tsQ8MBvLJcqAmhW/wW
17uymwPGIhYDKo4IC9y/+SEvieBPK2Z5NogenUs7oLPCco10lJY+p1E5AKFGACM6
qkfcRW6qIUw4333cvyXo+Sp0/qthwKTMhwOXJG9UmjVoHBSjXoRYLKQwc6KzbLI+
c89FCeHb4EIoWVmo/AevnjBLtixf7BRsrsWoxKniMk1meSJIWtcB1i+riOtdZcv3
u3qCG8aHu9t0TXoa/k6wLJFLV+Cr9jT3mUp7hi32pZNkYBVn0GbIVB3SC2YDB5aW
R+crXgqXEMP5eKmNRpJO7KauxwuhNIZMgxk9Ig38ilvE5FcN7TqRa/ACjmVqJZC2
ox5NshMFN3RxwczMFFaHuFUBcM+yrydlVSaBKHc/KzqUZXjPUQ0P4K3jGyvr+/uG
HzF+RlWMQIXsUtRhwms3SpC2gi+LPtopgdFJJkgeV47AqWAocvbrMTdnbfcwyynX
sxXtPoavOTVT1eI9NuildUfq5mAKaI3+bhBMMS8LbwaIIazzXlsAgqe3+F6linpb
nFq1ag7Kl+cgGOashIq7+y3vMJ3I90CMOvoPZ6ytpR4V2dZ+LB08fBLjHGWZknIF
b9OAz5i5VNIFLZR4CUto8ZdABp3Rk4e461l48Po/XC54IeTjqKN8HxUNx6kGdivi
I7lrjD0/zT/Vy21zIxdSDB0eNKcp093S2ftoy5or5PCzC/VRO8PpUOp9x16CQq9R
VWA/ijr1A16qG8KL8j5vud7XBGcQk39uqxGRwksAJhey+CtfZ2n0F+wr7Hl5MPGM
k1lWltKUp0SkfvpWvwxaxgRneoQhdAkBLFtL0BEW4qJUFjJHJgPMqHgBzXjccMGv
QtMX0M/FgwS9kru/KIc8dBi3nQVWdUOuP9doviO0zUfT3viSbXXDDscoek5Ax7sl
p8M9CmtluxmuZjtXvenswxBlonnJytG5/7J4TdvJvO75lNBcweGnad8NuizFn8/E
DOyMdZuMxDXoYuh09QS29K2ONE1w4d0w/eI8h5s18fmBA9KLdeBITs0VwqmUx8kF
Kvb8H2RfWFFSnfS4GOCI70nLzpZJs/SzWbqtC0AOMzjszd3JcMQhTggMcKztiDHZ
w3l92EvCMAA4fLzXR0K6IfV44MuOeX08SY8KEjpoWtD2X83kjKOpJXC+U+qe6L4I
aWuGVyWsQ7LOwbdmuWDpahqQdpjbBC45dUU+vtGpxVL2eQ4RBaGIUEfM8XdF4JYR
4HBk5/znPzDqUt6/YDI0Uam6pXXqJ/q9knPZHswQkIVY/vCwDa/wtFs122u/XeF5
H20MDdOHuU9PjmlMss21jXjrPLoxdamh5tmc/h9ytLXTdY3sIO5ZKYOBOf+BG7ML
KJFGI4CQxkbVSOJcdGD0tZ51NfT9KYqK3e9/mH1K+w7zlEfkJaqk8wSrZdB0m+4H
crMa3gRYUAWwIH26LheLCh18DYENKImV5I7sMsx9bF6keLzX494GXgEpuLH8tUKo
zOXZ+7Duu+iVYQDA4EzcFBGGbRPXx5/Q0Hv3ZTn9LJWyfpC4nTFe2X7qfVvW7UVC
6v1Y6MXAlQO04+p4mekTSp9kw0O6ZzBN+UmsZ1vipOCftqOQmNCif4yZgOPAD+ne
Q8TiDs3A4R7OkDABLShAodZnw/Oxd32+EeRZ6X+kgTc4On3nJzC7neu+kTWfAA/d
3iowdLYUQnB6KW6/6hkC5EPT9PfccpOZqTVK7b3vzBHk2mCRRRErT1EQ50FToTg2
2D3wlehJB5nf2DnqroaG53efgUBk5Z2WWmjkrVUZrz1EXSoR5eSdHc84Wwr8Emto
NRLblTsAUZ36HeR7reAZkBZPXHLyTZPkBfMd2G0xkP+1ljoBe8KjJPyEPwsu1JLg
V6mBLIkJ/ZVJi2GvPP7aBFFDnGSrguybmSeTNVCMZrwWLcvvvRwhd+321xNqLdvq
9SXF2nzn7dSQHliBGJg8K4uSLjMLgKVcHeaEbnNyNFfLLunI/E1vtdeuC/l4Cgop
4oezHZ1fECxMwBhwNatLeFJuMp5anA99Xhc0GWBmsMphLupBUPXTM6fkXHjcSj6C
3zkAJ+gTSIlnGosgEv+oefg2UhfrbSJDQ4W64RPIzzr/4Ka2kq5ixu/i2brTEev0
csXOgxdt9bA1HYabSJ2SvYF1SO3RTddf4RrMWpxjixloy1cKfvRLu3TOiDQdBSqi
j5hBT54MSrq8I/lJ6M8LQH0YTAUK/sLLPERQaz73z81h6rZNMcyN1GU86wytK0H7
uGz/arE9aeJ2rFEz4AjluH9/Jo3TVTVIPWppz07WXJxB1Ei8g6YhDUBwSJsNoRgH
SHUG/jpz50Q23IYvTFbhSepbWK2PGLkp01eRC2Vm376YvdfspUybJef+jXm367Po
lyBcRNVbbY17Ffu+JKd+EoP77GHeuNtj6VhWlBnt/1ZmmBjQI5WvF3ysv+tipD4A
bfh63rtTVE3OaqaUNwqoiWBDtHGbvLjDZRp0JRoQk1E8gMdhBFYMZ+TFLzpEFdLe
6m/75MwlfQKmljK9AfRfBlHGdnq0jKGOa05ZzBzgNPbh+7Y5JAJg5cXmIXPAlTyp
+mzh+p+81oLBkUOzFiibAF0SJlK8YB7cRsfmiKbX5yK+A6WzTy3TZ4C5t3l21V/c
SMyLrYpUlPvjx40XuWG4zWf/bkUN6mohMfZOLJcjeCO0akxXZgZggbGm3GF+KAPP
VSYpshY1uVe/VUWzaxxRD0gCZQBl+hRCJY02XpHlvjFQ0yChzgOlgmg6hHi1Em8j
+xJbCoZC11iCqOivTEkGjKFiIF46JU8O6qZfn4oBWEZNEmjGohyU1MFi3VDXpBii
iZNdlLeB10CD8RGAxu3LLw1wbBUpDq5S6+opUKpO6x/fMKvyoDhiXjekEq+AA4qf
G68jk/WIGJvgH4Q8290z6GhoHCCgpiaVKShI5jpweczYqA8OImhtsLd6CmZru0GK
xFkNB51+7E+l8WsIC4RQFJSooz/vvLCzqADuqaYUL1OyDFUgawJRPvo4joSF3rZs
7BLsWLzW7khoK9vaZUI3XaxHzYK5Bgfy7PHMdstfsGwsRBoKb/omtBymJqpxrlDS
s+0HDRfhaNdMaLxbj4WZMcH/3tk2hxXeB19ANt9O4MQsUQP3q/jydrY7Ccp6tjF5
RlL7Jv7oLnPwcxh0b9zkS3jTv/EmQflOqI/0NcnrSUzpMqew3XDjORzP2jVlrf80
8H2s+UrdBIarA7+bA1z6/6HfpWWAqzuLwd/7cQX4SuX7zut8gTN0R1jTemo0M9Ap
45PdJqSAsbgueT2BXFnPjIseNvDYEJBemX+yh8KsSsHCWhfNdHJbpd58//jIz0/3
HL71hMyCyosiWS4u/eDxBMDVql2Wej89LnNRAI7S7eT+BAdVTwhRVE9E2BRf6FUN
CUbfYAhvBtxRc6VWuYZUpLniSthTu/KrsUQFGF7QEBaw5lrNtHXdEh9Hgew1Yz6h
EUko/u4zrZeaeYV85qyPSeCfsayiZ0UasJqHRfa7nEXQ4JOxrUZg1ZK0VhWzCObQ
DZryvZ6t7jXWBLmPn0j5EnUes7Aaazb7LhLr9DxSCAI6lLhP1wLSxtg4zrImiocC
C79wWAOk6od3iQFcJ/0PKHH7XJFZk9VBTaqyl9cAunReHeV1rRkfASFX6YfmYgNv
QDlyi2F4yasg77UIIHjn7ASQYjAu7AuNaY2r7X5z7eJ2gQZJHpE4ypwgZwS/vvfL
gl4Oqfn33yBeuF6LtgvTsPFB99JTlKZ/9kwLm5qyrKMuktl8ehST/PUog8fjH4gY
jp174T9LgZbnW6e/hsX9C7WeoDxuVr4sdDJCKbPQAek4tQKb0Jf9mdBgky9cBS7k
puFbCYqjOtZLUyzEPpv+lPnjoz0R20QIPozpTlbpjrW+EXqkRenNYTcCVEP58NFO
oaVA0IAVV1ujPTn0C8HngIr25+7NFEHnACrRh3ykI/Z4AyV6PrWU0oApSgcTF8ao
6wseTBj8KK5W3Ro0KcSuYkTmG7ESqx4Hu0QxCYAaV9IMongW61x/jzb60HTU2rAO
ez2Ta9VOcEb3ROLFJTbzLuDZ3X6/K/9xOKjWdacVNXTkKhSSm2ZaW2temBqDGreK
+mx0gkySQxMhgBYE+laXmnaCeWMeFwYBTgvf3h4IpNNLYuqzDH4BiwvhtXnRdO6V
EfwbpLFBSumaJr2OBPl3cal456YZt9DdRNDTSvyAD7a3dYqzVO5A4XFX3dXSX4Jh
NumHM+V2MdRycLEcf++v200QUBF/oOe1upsNXFG+IkozH/q5ONNLIlJ5lOoC2Vdz
dDvyIVurJv174NBg+blXLm5z3JBmVuiqDUXE+SH6pnTf49CwAVprhyTEvRTFfEoh
bWmZ0lkMRKJA0raPEO2r3W5BCy12CgR8jiaahm1eMfezyqAKcEtDcy1YWJAtfi4d
kBsYMbT5w95v/zYmuCM337/eLVmdxPNXnU9pazQakxudTnnvoFKTbPApHvij45Le
/h/0yLTK3eYqDimYNCZl1ls3L7cB+TwDDaIv2HNQ7oZjC4yJaqdQSRE25Q+aYt4o
mCLM5sHTK8iCKJ1skYO6DHsyKJ6VFNx9gGw15uM0yxXkW+f3AsgXck6VVmVM9yxr
JHh2i9+PwuYqLxFoB1vlfvzZcEgFSHJEfz5W5fGMeDuZw6NXZtds7jJgx95aOpk9
dkyofiaYxbIhismgvpg0R1pslKwmSmLL2KHQowIUrZaQp2OWGF4ydG/T7tRZH7u0
Al2ohXNza9Ra6EjMMBvkjb5QBFlGRPe0T3TaN9WzUDWWAY82OcnH5CPQvF1ToqYO
VJ+DNG91UmAlD03zFgvak0SzBb8rNffJ8OFsLL93hYoEdKYSB+0dBp9rK0pY1wza
sSKG9Z2x4/MBB1iiIrX/TPWFn7Y8hpWHOtym/9XDWYH4ylD0cHg6S/rZTxdFe7hB
9nLGfLD24lj+x7VFrIm4waNpj4W/7dDAiyd6++JPXHaQqdUoE1hhLL+fgEnh21gK
27RmI8vhuEu0Oz6Mn3NYNyT6dT5nkMztcAZVRX+jz9nOJSylen425rbX1zQJQEUw
SnIE4b8tdI2Fz54oI/Qzo8oFHQZyS7mXLQZD5KYJzhNpjudx6tbHCarJS56+ufQ9
GDStaWXA4PU4Z7ZUy4Rhy6szRqsKl9p+rL7PTZlWxVWPNf1eZF101ZiY7XTIiHLO
ZSlZP81L1Vc8g1x/9DL5wSzQ09/RjN3yWw70EUM4p/S0vrZUsvW5TPSIaKW8jUx/
JWdMiKmDvKg2/YtoBMhBo4WyAnqDifhufBuWWncAiDA0ssdsV+0yAtDzPJ0xcaBl
oFlWVsh7D9WJ8P/1drP9cm0MvN2gwwjqpiu8OpOxuYCTrTDgi89xOwQjM0emVA7v
+P7ZEE4Tx9nNo8qeRqi7EueT8qJ4iwZgmubgtRQ20zqK6/NYPmaj2UFqwp101C33
B5xRV0MJELtdifwghDbeIKfhUv7AHGtdeZoP6PcM5dJWrkyb1aHY/r5Y33ZLz1tr
8+ph2NpSBghpVf1H/uXkBeiOkFpzPIcMBM5AlZWCZ5lkZWlDWGlganreQJoTDTgj
dINKYOt07B6yq0pi45lWuiHwWmRfcsKw6enXGGZEfaVFH5HxByuFb6W4BQg8Zuhi
znWPDZXJyPsSu5XObyD/VuOwIOxa+J3PW/bbwx7NGe/oqQb+unSXYgw7qLsqM8rC
z5YP0QohjvO48IvlqE7vU50fkz4InxMZRnsJe21/Dyf5IWWvkSV2nH/AyEeKzoYh
N7aAncOQWin2wYAVjLo6C2CVU6p9wODHEMqPFG59zevToldJVHieMq1vB2ZpfLJi
jrAouKnr7c7uW4iiFU9gz7h5SK65frQ6ZZgZd0JfajmlbzusuChNQFxs8qG5jY6R
DgtFyApeWduk4jzHKew4uYNXuN88UAGguaj8/3HEdgv1TqguafxW8faTYs74QhVA
d3z1yIvgV3gMeaducF7w8RQnUQRDEJyBPnqCcKnAjCa1+Bdml/FcKfBEkHLEpv3Y
UmkpefCAgxdZyvHE3S+IvcHJptrD87gK4nVp6Vjj99VF45sZ5iXoJJ1TLKKa2p47
rjxKL9vTNKO8W0azX/8/+4K2pVcRvoAI0nMAS9G4yy2d9v/Tmn1U32GmPkNSi9MG
lf9n0B0tsMaZ+EjHZThopgwZ9dRjJ30WGJEvt7pBoosoeLP5h2KSLkhUiMhpsD6C
ZaSWEm37WmGAY9xMG+mlCLS2RPMBwz1hSHa+9Me3sZoxl7kUB3KzV+omfKCcvGCX
0zxHOv9STSFq8Fj3cOO12Zww1I2sG44DS8eljuqvvCJ8Ow3kgl+rTyt9G3qXKXiq
7KRiFbzV7NsFvSAAjm6CL+fpUYN/z4v/Lvd2mRTeOnANN5IKdi6R4YBCeFmmYQah
k9zusyx+kHLc9n3qPSwiAG0Rwl5j8a9Ueoy3N9o481oI4Xxi/EavpAjWw7ILvKRp
klMSUpQvK6Hgz2NMek0Vh6o7JhfTz5cGuYEzungG4BaYz/KX19qHZ9p63SYWINlu
KM3JymlAlDWpOQHZP4cMGxwL5mnLYEAA8uixWjRqNdHo+wW1NE5/Xp2Et6CCw7Np
kUcThbYlKEEwNtXpZGIT3Gux4KXKTbGTJmkTGMV6IDMoTiUQdiLk9tLsSMPx6BjL
qrk6ar8vjl6ndU26QBeQxezzTQbB6CgxSAR8sVg0OaXSGfc9ozpwrPZo+nbv2Gju
M4ZL0RieVsdg1Jl+X+827XWN+enzKjO7cHnjE11uECyShRkK55wPJdM7AqFZD3uA
YRB7B5fPu6k1dcNQ0p4NQGTRzxj1R8Po5i4MjbvPszHzqf1MJ7ajgqNC07UcvyEu
9oDlAMjUFobzOQXqc2YNSD9rHGyUHYapes1hk5cRnYGtz74NAWssTtdqkBDBJ5u6
KROw9Nv2uj90kdL3XoE3+EhaZkwBZoSnEnnw3pdIjisBmgU5s9VDAzTR8DxIA613
z9aoEOzllCpFWJhLI7JZQ9b4P2Fkq4jGYRM3UQ7zUklxA+UIkuCo7IeE5Bn88KaU
anbB9vbCM+u/ijLXAlinwqAHOA1YA8/LW9GP06zxm/ME/kRN8nSIum8iiBZnYVj7
xKt95YzJDObv5qwGQD6bwg61hS+E/xekfesV48M0QzCVYxaQ0pX8Lm8idQjzvJTN
mE2UtEmGe3/m1Lq3maLmDrBY2r2+uUjnMg/nE4hI3HbUlHZ4CcDDE1pTvPqa2zch
8OyMcojTDfqK14bDWIYaRqkFo06RgbUYrED/SlLv1+8m6JtsbEN7Dad0Y/80VZuE
Q/pW+EHOgljrxfdVRPsnB9Axed/ydKYRfWwNpt3mrD/HUtm1sGM+JKMAt2xRvX2o
6VserYJaZFhDZHAQldM+kCHrbVwFaLCcGJ+zRisR1bhAylr46qqpqKyeUqHSTQJZ
DpRc5RPQUVqQAMVJPu+dNqcHZtd9/lXOHx6zEaBYaw6hmm50yyvEf2g+DtaK5KxC
Fwlqmy3FJfaEM8OvcWgbW3pPHz0bmR3q3lTRxzAfpQrcdObVeLSOptJr5B3YLybf
avOxBHHjT8k6SRTs8aQ9CjG+Oatb4i5LjHpQ9zdRcQ9nkjX6V4D3h+hnQzkANwY7
DssIiTo9urge9Sz36Ke9kxP34sHUuxFD0H2xupa+EOM8eKUXga8sp67ckSEtToDF
1hLSyXL6iRYABfGollrf0+8ltU+0TlRzmpODj7r1FNxqRqA7j2vrXJ/WVv7fF+0Z
xew4VAIYkolEu1NTC76Y8ru88WamYlWp/MzamHWtVOff/od6dAIaBwqcxWihWkjm
5BdFWxSxcVFh1O7cyKBXNkPep055mhbOYckYmOoScckZOoJtK3VQEPdgl0A4f5ir
pkqk4jbWghlOA/VySotGvh60DriIRMrPt1mTHjlSbIUv3XGL5hJbb7gEFbtyJAE9
i4djDJydLXAi3UVRjO11mMwd5lp42dkuV+tx996/n/BcWjTHijDN4BjcJXoCAJi+
VvxYueFbgtvaD1dqIddLErnrgC1yp1Dx8/68WFmAzQsBGyLE9vRBbQZ20WBe+RL1
qUmCDpOCpkLEQ93alyhomgpX0iJ/+vyod5Op5ji9Rw7sWWnwj9vx/ccIgGJ4kams
rt0xAABoW/P5KW7Jre1DHICIrAmK0onNuoj0EiR9/ewO1acBBl5GLO5eFlvohGsO
Ij9yc6M5q9eojTvC7I97Un3mZMb4NU0RsbOVQejiOSsF7XzGCEZzccbk37IR5S8D
5dIL50fy2IM2M34IsDOasOCRBm69nw1Wgi+V9X3eiMHUzBv/Qld5tSBJxJSXEjGz
uEin4dju6D0SDHfwlmnK3ft7yF6DOC9JleL14Y0RQGqQOgY1PzoyvWhCYDvdzyzy
zSFSUSdICuWqjNAJtjRIDMkN79ZfPrVDLQ5AKnddcfHJG/mbTGhTYAcMeSut82HF
t0tFu0ZkiKJQJWCmzKKDJP/nq2DUl4mnZsJHT5Ak1tFtViHk43cpeFmETQuK17z3
TcBzKkB5GJwf868o1QYadXpdYXFLYrohJcqpTeHg4FMYLT1P8/WEGXAGkvC8VmXz
k+Ds1LBBkYii6GxWjI+Naiia4aB5SSTGCUdp3/U4vhFdCKo+hMKzRYE0oGu+8hIL
7riUijxXgw+o/R89SGoeIa/LAybeV3cVD1JAyYzpOEksavSrmIgQTyV7KMDfl6fs
3eYwKrpjL56sLyXBLmASXb1M/kZ8VMj/JbK4p3MnjQ47f5/3rujRltimDjRDVtKH
vf7dMSPM07H2D7HLTroa4mqVbq4W1rT+Vb/cdZ3jURqOBHE2dtMkE/Dot6EgHHXg
xoviK0gD4RXEMiycIBapt19VdQxUO6cPnQrEigE94+h3w6oAh/6sabB4UZzeeRpx
n6fuA6Mv410BplPrCjvfsm4xuWHSjnYVtBildmQjbUcEaTssDnXVKOgUXJimMvQV
hRvwd/DfODIpThDZvgEmOMf7YRyrYt0YxieqlViV8BRSaJ/CQqisDOYNblEKt1BF
1H2/9Sj0j6dBo/CwOqTrcSmeQiUqEWTQvH/o+bSiX2mmcqrBkXoGcIuaQ6ZEaXgE
dAVR6ztlLgGvVvtQNTbPAj9DwKGVIyOr/JT+0ApI4G0ooabmHEHwC/wZnqwG0SVc
ZwWdi4B+ntbj9TrXQ5NVG7Jul4xvR6PXKKSFpcwwVLs2KUIByvK1Tb5Sy0Tky/WS
uudxIn+nVjIQHduCZ+lW41bn5ZQDmwf/KTYBRwn3tXeWBEk4ztxjfY6SLvvQlgSM
p2O6ugjfjIc16Xyog0bRwxyZY2iF+kNGG5G6g2BigVqEwQD+Jq8WwoREeTUikYRO
CEIMymCBnOGwp/tO/B/XYLWCyJGYtd3X9sLMS5PD6rx0TQpNuqLBLVsLoK/VxPJ7
gM/WNcn1npITJfuPkrmnMg2kWblzrnNeRCgemzhFhGZ72yNu5cS+0cJgt1wTW1Gf
RVSuF2ncF8fpWZopkgT2zXqarOCcmuOG+g3e2pXRAtyeU8X4UJrp8dRGu17WUZCi
sDilcEO/8Gy8GVTZn7suatugx35qtLGCFwyV0N5PozO8BGFx9rsrF0f1Es/CKVmH
Vb7YY+wvYlafdlSorzfTQEeFjeToFBqvcmF6aqgOC3c1gRiSHhKnZL8ydcqv5ywj
nEfnKn02L8emd/I880SCUSrKlDC3mB1b7AffwjgIsrsh6xslSBnHJlwv0M7kfDXk
pzPLJr3R2SfozCpwQFQpQVOjpZZCR29AdHKC8hlL198dDRQnnEoVUEGKbP7enajE
OhqvLb2y3wNkUxo5M4XRiNyuvONIxSW+WptV86/qyfVjdzEY2Srg4BoqjDjC6DaV
xtWNRaCyFCj53eKi/0Ho6duIMWUi0EBQT3zeU7JWmbInS5nfcwwdFZe87NPGYl0S
m1UrWAnRs7x+pUOP/88qUgy3C89hQu6pJUxa2uDndvJd0e+dA9tQt4qRSaE04YSQ
JkwFk8K4Q9TOSH5NLBFd7wp0HV376uLvX4Yi2GZew/4rDXnrJphSd+pgdNRVfjH7
hit2yreFbkReScfkKFs0rUYJVFzAlvnIL+XCvPApvzOfK/SF7zb/Y+Cvr94s15DB
mkLX87k6oa0IZZZ4EViClfpHoEPwPnBoWuVtT/ojxbhFFJ98cKhebN5wC1A5+Q6G
D/rN3usXLqS2xz5VWaJcY1wgJKUOr2SvbgDGYuNrGkr9bAOHF1EOV3/cH+Tur+7Q
lgqulqRHjr9r5pqmrVstaOxsPHh9L9q9VXq1lPGcVgmOy09z1OyLTEwShnDrVq2B
aJOkwlX/dT8B/bLlqu8CQ4mCPylp+X8UqOI/Jjxyp0h8hJewco8vCNfmx51k/hI0
vSiME+82PeUy3CSL9whp/fwX9diRsOiyguk6Wf5wWnbNOZ2+AhcbwA8ogeIlDpyP
8kAoULlcSc+JgKNH7S+B7N9Ul56V3SFyXlmPs9rRj26BMd9ihQzk6UbQBSj/wMje
a8WotF8MgCgwADE5CDCmchcgTBwN1brc6dUS1T7Jw3oKBP5YZg7XGv8WqGQ0hDwT
ynELXdEj2SBM8dikrK7ZovzN4zvjCQfg2QUUr7jvDsCAdeB8Nm250YA+eWwgHtxj
oTTetnmeVoHgaWBjnN4Vs0juPWp6UamkygEOuskfQS6ZJsZdHpep8Jxn61kj+Fyb
eQR1yTJTmR0C43zS2/AZZcx+bAdoQ2VYF1GjHgHT8Fn6pZXU9Kcp0r3vxGhYwara
O8BuICbDYuRGzetwdY48tsqmfeawY7/GxYjUuD3N7O+JZPN0Tov+ln/sns5UIlbf
SvOMwy/LFAZ/2tU2QTS1UD5jm9+BZfyfPujVotTcIuovbCKfGcb/6wsPcLbrzy+t
QcJrVQCBShrZK8m872PnV146DScHLFLY0xJ7LQZeYHfGQh16Xp4fy789DJSQ9X9G
N4bveXqZSgxX5j2mxKmfBXYE2EAoc7reHz1aQHH/l5SOBi32iIYo8oiD1EheDzPD
6reSzpn83cOphm9fVO4Jvk9NK0jX/JS5TsxJkHbFqx5AQEAMGUkzZ41xYk5hAO/G
swkeb3gBPG/lnHDKTy6xyxyWVkMvvVXDTeukW3nrA1cgHQzWsd2BiDyBWrPicSyl
6fgev56+SlIvTrA82tt6ofA7PKfJ0WaceCznpMwvC5by0PfvRpnagbuV3lAM0oDS
GSk5YJEaUXdF6XnfLUogDDFP+4EIMr0v7K4KPdR+wwZwcDlfQ448jA9pEyOt4zAi
08xTmHFyMx6MoGFp8Aj+2buFNeP+5529UxaXTwhzKsEKWo6OSbmqxNK8FAJiFo3s
53X+1IdLoQJN6YKwCu+YbJ8r1NFeOTJH0WhqwWIkZA30p8aWliZIGiAHfRahRJTh
Ww6Wjnx88V1IMKuqZbJCM/wbvkDE9sAeLvBkkm/N2txOjAzEh8xp9xTqHrx6i9Qo
igDvbso/cL+K1MIaFVhxzHkkCcjeTmg2rClI14C9UAq/rbdtpJmlKipbIMM+EeSV
qDk9X2nnZmtv9ijGr0k94oJqxlxkp7ncePOCwiM/lIj6/RJ6LEUZn55tgYSmoETw
sNvUomARqbrhBPoGzlzC5oLjOJ7fWADLbcyTS9oXlrQFmOwLEZDY3eXOn4S2CfMC
X/wKb/7HPAyv1AlE+0g3qXqE/O0mdR30879kofJV5RK8gt+rx8cOKbeQa5CKHrdS
cVmdO9WaI9aQJ8X80CvI94WacqlC40b1bh3b0Zm2aRD7tMdrevjWuKpv2Pgzjlxn
TOcFT6r1/o2HPFTtTdQi61TvtKPm78llFgFaI0O0OsUr4uXovcrR6El1IWC5kOSJ
OyskZHEoLIh4sCc3n4Mz0UyvQTy5q3fXv1mm/9xtcXLPRq64GUkmTNqiORWn9l8M
t+it9sSbUTlQ6rL620lM47s4M0UwY13lCkyCPtBMVGs1Dn5xWkqG20jHUgrZRWKI
29Ax1zZCxPD4eQaxqYjBcZH+/4ZdeFKC0Xp1Zc2esBD2Yi24H8wwxsB9eBCfMk4Y
pDQgbOFVck7b1V7ypXMrM/N4DQHxGnmEIcuF/L+h1RcGnoBuXB+ItnIvillrpz5w
7xQk6H3Yr71D3SYp/Xym0DPZNvODm5fUA+xAsBl9zTJPd9n8qC9NwvPLxJF9XttW
bAHm306/vXOLsC3CqLPxmnwYc4Tx9THGoTcZ2evnWuhFgbk3ovMSUvVN/+U4ab6y
B715aJ1hZPNf9WhqhiN+SeRr2QlSKYM8Ag2aRsoa/qNr9wkmSt0e7Zc2h8qGNI6c
X7WuvS7yTQ5ui6/dNWtL9S4kZ53so2oCrPjKrgKYTEJyHeAB33AoXoQvtjYP6fBX
u2tQyKG21CaZVXhvQx8m6HjV6sNcIaU0b2g+wbDzm1rmjWEYCWYBezp8SjCE3+pZ
pyzhOe9ZJwFmEhVFCIw+GXwOaC5MRx9/yP8sMSAq6qsSPNgE2OgVQbM1nWiiYs6R
aAusTb1T6suf2o0UFsYWITS2D+FQJVsGhvJEsqYF7owKBS3VMjIk07kBkhFIVLZs
FK4KFuQF2yrFxhpvMYxCjCDPddtxg45oy8+CI+HuqANQ5Zc1jki9U/mOGObXDk2C
8bg/Uq9e6LihivtgpJuuFr9KeyrLIhsZoDWWbThxe8AVTwF5LRa0REYAL0aKOj7N
ikJCb3ar+ZxNO622us8uQo5tVF98HxAdtQ0CV5WqcYyIZLHkgrkDX/GiSVLY5QkB
V4xwuJUe5oHfJ3tVKplE1dZd8+3p4F39rGQi1Dpqjhhdt6B3DUC0v8DyoVgeQp/l
Tr86jugIW6w4wrrHpYZKJhtYqe2veXc2RvqJAb9daTDCFXF25syR8ykm64I5kRhh
48YH1pLzYXpqdy8LOU4FhfqatqMGxDJk+tme3Ru0kCuNFXq2x/tX1xSHF153ClWd
k9I5QjfjNxjgc07xRZhu8b+VQlRpFO2hdcJqgwQYiMXMT6IxOEuQ8+SxaM+O9T1/
Tnizk/Z7d+ua+WGkP89+X6GZjRLfwL/vBiM3woOvND5ajnbbLTpzqi/Ymzk6sj2X
KH5aLe8sxh+bwnNnwWOdpSqNMJsLnMcFfkEd/DIpw0mPOGVpkwNRmxYHhzWr0w4G
Y+bXLGsUQHEYPpLHdO0SMRgqR21LrtFJuD4NTsLOoB/VyYIYHg85inhOSn903CNa
ANTt6QeYtZP0c0vUr0bDqxdTW8LPPuT1c0wuKsNylQ6mK82cmtbAasq0qNuaaxin
9pjMNbOY+GyCxVCJcfPlp+VSc3RMRXOOeAKoVVcDPRktiOeFEd9jbxAz/gKhvBSo
HB0vcFsZbwiRqT7+t3XtIfb8Q3z75fOEic1zW9MUpX54TvSbPXQ4pXKmmitTKfr8
xWdXyud70/4LhPyyWgLXksTr7cuq9wLUMidzx4ITL9QVRRbvExEBfF5p0N/asj+z
gLlvbJHLV0rG74xcJfLt6IC/T14ftmkqVA8F1jJpGJzO6IGBZJuXu+ydYsgJT/IA
1ozkvNT4/b1OtGiOlcmzekps7/9D5U/oLHVq6CO+FJGnc9TQ2AwErCeCfcyhFnQ3
Qx+NezMfLjNTpOGFsDd9ti3fRO7IrcvmKhapWjHuX2kShQ/VBVBvQt0HzBndVrTc
KEUyNqqHN3g7YBfkw508T4wnTN6mA3inn5QnIaiAhLlWklbraBylNYT2tdULrYme
hrt/FJ57Xym3+ndi7jFqBwZcQ1+X+8xQq6X2iQ9EFkGj9JUAGjNQ4pij5Y7a7tJa
9WCBUK+H6d2UVXa/Po6vp2dC9PRzdVdj+sC+nuDJeAp48h6xIyDGue7ySl/5cTWl
UOtUKGZzu6qzyENDN3BLPF3/O1Hrmh2pKCk55FpEPsPRQPUyz2u3IFCsZHI6twYf
cEpv1Haur+c9Y/3Jc5zuybGBcYhA0G+K2bioiKuHYGFNQFj9Bwy/tw1Rn+dnQwQ5
15aRDrreP0XUVafA+ayyRWkeLvTDZXadIVb/CcaMhtb38cVU3YTxFXJS0v8BNKbK
nljFg+fckz6hoSdoHf/rGUEFIsOUL8+NPBXyKfT3O1RQJuX9Qd72H0nYBSP3P2EU
zYHkcYujCo58yAjU/+ymRq6tp6YPad0lBk3mvmKHSDd/6GR+S0jyO2bn/g1M2rmD
xYV0cnxz9Ka4FkGxb1A4KB5EUBbSuJvtCAuIHs3jsmJVNPD2NJ32vFK4E/JNhtu2
rxAQ/QOXhjtAZ1lQCH8qfslmXZ4vGNssVuV461q8PVRCE48DybT8T2hs3QnsGbG0
P63iZ2gpo4YAx9uexlt/tV6tm6j47h3sYSqP1nSWuL7lV3b7FkFJSfZVjK6nUhcr
ebJgJPvdYDpKWvLquJQghUiQhqo1euHfTl+kzAGLxejfzQBnD3L1w1s0X+dZzRTE
tr4Qx4StFl/KCQJCc3lK1iWEkOcOIB3f2gOFeFHbVpO3KZDKQEBcmas0/1mk5M+P
HLnAidwPpLC66ZzalrHEs+mfkoESFvt+hSXCCIjFsrIsq+HVvWZ2FQ+KUm/S2uK3
l6bKUia8sJW5gK74yDxSCKfJvqxqA1TzA/Yy6p9CMQ2GNAGNTNL20rUTwon8NZQU
Lxmf024nvLANeNn8yw1cO/6bPfEXA6mi/3LIRYG0Sa/pkeAOPBVpR2QeigLHoZW5
uBcdh5Y53YvXzv002/IDcLMc4bLfVsxkSbpSRMkfkcyHaeI5qqOXglndzsauWMey
gJ3LxAu9KVHAKavIt2DYwfFTBlIKzqaaGAPtwlfqMILJN6MqC/Ru9OoS6arQKJc4
HnKIqJRxJm6W5eaGCNAHIPlX0S7lfjmvQi69X9+Ms6ueCqUjdkvTRRSCDFDbN5D+
uWG6N94yNHESeifBT8A+UACanu8rQvjKEWXYHZ//OOfAZ2QPrqFBr75avIuJutF8
MGOutQjEmqzCqbU9xVfsF6xNQBR8HW/VCbPdf4vxXxDo4yC4QVgxkaxPC6A5s69K
c4vhL8V/ZMxEFA7cHBJpFXsWES1YebLm7KpcSnrgUQJIJdtshKxy6obgaffhCpl5
QFgY76vHWS8WPlo/8Gcqgjz3iPoKYWngKN6+3zAru5z8yw8OKC9gAO35+xZI78H1
RiTy/DLd/PDS4fnLOzmc7sr8D2vL6ng0VGl3UU/EPZ438wRy4letxjs1KhN9SqxA
3tFtDZs3q2rsR617Px5Znp2KBw6eOn8lVzqmGxfpnAnqjFl1o609tDiBvMY3G5Pp
2+Zng1hMmuj7at7Ec3UP6JErceHwKaveLDNnJH6rQpY8lOO6CAN5z5FA+PUKaVMM
5jXFGVFpqtI0ADJutjBXBpe9vYL7apvOZJMksQ/ygBSiGcpzKcKCP1VdVn116BUK
u/CNd/w1PKqF9uN4W1ZfCQE8qypY49gS9dxsTp/AtbPlhRFvbb0zerW+DLJAqy3+
JWXAfu3kwBy4OorXEyVOTy13YFRMQY+1zt8fpammWG8GhHt/WvX4mZXPDlcCw2kh
k17Lv5I2OADAbTrd1ewZjqpUnAKzA01mPjtlNlTxbfwhI8UNTcLzZ86hBo3L4X3s
/PgnBYR/nX2O/9PpLReS9D7Vf3yTosBbC9Qn82wTyoftv0XIgcklY41DYr9mr3vP
BqxuY2dXOAcoxAYeIBtVqgX9UfTOeLnjlIBZ8wN2wVs44sokzEBR1i/XK7wigOzA
EEDajKGqAH0xRmOuq8iwguO8Scxs2XGT8wNk3kUOFfvxKpMLAsl6N/Bug2dQqsfO
D+Ipbxs4hBoQFhtrb56eTVuhb/CrnZzyK6EKtVgUcWzDabDFwTAnGo4eoczC+5co
hqRSGPaFHhX99HOyLLH3oewDrUWUlXhNeuenLG54WxsbuFw/h7bkvbXeV56BiZso
VC//fRqQpB5fLcT1L+szzdi4eh7LFrEjV6M/f/WiqvRly6Bt3qWtBj1Fruc+fmmG
mnZQMjX2gU9N4H7FlD6oECVrVlo6hWsBEmcykONJLZkqGIOQUE3mA72CjjX5WCAb
MxNhSE4Sur3ZvK5KIvM0ZKQkaUPAkzeG5LbY7YMn8qd0vv0TrJZUVbK6ZuXZlZ8l
J31eoIJXD1nPVwuPf9LTq3S3VM2luA7Q77ufjTJMveAvZiMK+xlQxTK2+Fj/YLPg
F9VacvSCKvSfsL1r4oD5hST9D/Fav3uRP8+yrwD/ktjFqdK35+iPnInCs2hJKass
tvVom5v9t0RZ2Ves645kBC6ZyCK0GuTajSSnbKNpECGtUTMkNxcx0Mj6UCc4tliA
CWdbGhiqHY4S4nVf+8hxpo/fU/Prui9lzUyGH4wuZ0LcBhm4aEkWjNsRoZfsEPmW
w5fDTWQKZbiflVADQoZ6GeQpaAvXEI+esyvO+fPH3bdZtfG5u9hhipfPuhLNLmzO
Vuo/avBJRTRV5EIYeczLg/e6IyiP0g3RQUIzuupv4ZEuw+jA1NoKPfYcYeCmJFvs
QVa5L+caRS001tRNueT5z6/YDxY8rTHrC6rJN8oL6yKghmH8RmlSUCKoSBy633Xh
NTBgKWBt+Ic8uoPO0mkU0APvQen7jbcXGsBomB1ozak9QA9G6KyBLR3ueUrAxFfb
REr3BvB5swnm6jw6kIRqGKZYzUYpy8CWhYRbXw9JdLb8XJDU58yjxwC/3Td6MH9G
WijazAeThURFyWVqEF+WYdVLaStAZnmVR6L29CnUpJ1ajndq/wEqNARP3sQD2sz5
l9h1/4wwX/Qk1IJfRJiXhyW8ylW9lLpl2ni4DRIhScyuwstMK3Ctq0+HePkyX+zg
tKkvxZsPY/i5/xrRLasCaYcZMUy5+OmAel1pmIhlCa2N7vjsVen++OgENzJbGNa2
GCkdesR+4SjavnXN6fUzhFkl2YzQd8bD9x9bz7XFXOnE0dni2fAyftuJNlGMaHVy
FmRgst3uZtJexZT1KhZBU1gew4pMfbP6vovyQnbBAir4NW4kwbqX41yyl08M2LRJ
LAj/UzmRoahBC4BoPsr1RSmF7RG1BeV4BEs3nRiz1d5sqUf3dpa33JojrBD6f+L/
S2w6nnNZFLVXTcZF27Jqd70Oxb/BWVxyG/ooyU6glQNEIdFaD8ImIPHP+7L+8xj8
MmUihRdj0H0wmYZlV1GBkatm23/fRstyD5nRwRsFynGy3TA/o2IaTE3ExiHQ3h4h
vE5WyuWv4b7vKIhrLjuLXdwrcTx+qiI6HzHdiaG5M22qTymx92vUqMTvQj7rVsgI
XKv0grewiqYd0BJ2QIUFsaHsTQFggdc2oRtgt2J7PUMZgNeoev4AUG7kM8hXX2pT
mo1Km1DuBqem1OBq7u96ko4UBAxOLzM6EO0cJKOwfz7cRUo17WxfxCAYoFoH4QtX
knNnkRFPLXQRtmtYF52nF7tB/GLDq2ASLh3F3A6CH/18ctY+rIgvhGIV/Wd4kwa9
8vOEI25IzX7UTVIYtxsZlGJYXzMRcZ/yD8fzFj2IyRq0+NwSbNjFaOpAC2AbzDAS
e7RzNTAtqo2B3SYs4TrcSMu9jI8iR3xYwk5wK8gXAgUcolYzifHeCRH7MIygfI4d
QH0jY2b47gHX7P6aF1Uk0we+8fYdUKnHu+NRYnQI/9GraGOgTafk7ad9/SMSCc4i
fvOqGTlyzFc2rLNJ3tpZY2EOMgl+aM0jqmC52LiLxDwTqQ1MI6BhPaaKMyw5oIcE
wKeGSySTKIasZRmdu7Vb+ijobResiE8B0Jqj8Fz/bmhp/UISFQrxg5hShI7AVY0U
8M4prs4q2PmHmEJ46AG3LugOknqANf3wCPcfrCFfsoa/XNuM8IZuxvCfSOqw5OKZ
ljlocm0R8cywqZAJ2dMhhiCyEp5sV9vPi/jiNY0lvQNQZKcauvelHnQILrFGPQ47
GHhza+t2NaRQmZmrZ3ugD4ZMWLD60U+adJzG4ZXo+DwzQFzFjgz4tgV0okG5X+f6
fbO7FKRgEiwNtSDwGnxMsZcFc8G3beqXUWQUzA+ZpgNY0uV26n3GEV2AI8LC00SM
sXmpDSct9NLmsDfmLi8Dvn010LSsLXfEJsHq4n+y/ffQKWELHD+KqU4Cv/nSJCPc
dZdqfgz5Qii6jU03EseJ1Yyp8DiFbA7BOlHYNX+YpXiZxE/J/o9lP2A+cNpW0s72
dOsrMWDDsiEUFvIacXr6WmN3IK6NokL0VcmL1pkgQuq2JCMeMmK/Na4kEer3D2fN
8+s8KPM+9MZOCYRfL6coFbY7LFjygofylEMKJd+3ZXC+IMT927bFQBjsK4FHO5XK
hFUTpMJf1bUwGx5bBAdi02zETIYABCORyYyN08T50ApeGXjlFgev/PdkCd58iO5n
azdkf6zeQ94l6b298yoc6lNLOY2SxZLHUw+ILaPWe0jhP+//20ev0UzsMVo4Wr9i
CBJN4kMvLv4eg+6M6ZGbJ1/NAxeYP5MujGSV+ssgxG+MKIG4Q0Asbj881gV79avx
7booYxY5vGSz3svaqmWpCHgLiOSljoZZPee3M2ukJE5W6TJdiUqZliBF+mWx+esc
DVVg1A8a4IWbpgTpfgaPXcfNJCOwJK9I/73kD3W6is9yYiXFXEGub4clsmTog6wE
u00ZLdS1FEMhl5jZg/yZQbrq2XNthoRNZblqUHVNsGI+QtlCLCd6Ilx9KdF/wTA0
y8bwFCIFf9ThBj1djp6TiEgBUrGFPnwuQl4H5prv8VW+xjzvOrbtQBVT1bCFF3YU
VHetKN0dqiabQLb+VefR3msNfDU17HMBzCVbLYcyzfxl6Z8u+7WUzKL9tYJdWZvU
AQ/kty+OKGeNzzGknKfKJr+kIt2cgBlAGt7/N5gtg8iAEItbY7nPdwKyDFK+6mWO
UVDrcSrpidR2tgs6RvcldnOAyGzULQsiNk0po+WthHAPK7UPxFzaqKPn3+OAI3ml
U8uq3jLab/Nat/F3O/WTLNKvJz2E5hHvO4g9zo3ip9sRGiByLfLpDAurW+gUTJC1
/3lcgrU2dkYVr5poV6Ioz2UYOTdW5Ohm5SD1QT57hPRMCfFCUlF1p/fENanTlg0n
dkmQoY69zHtwQX41jx//Osk07/jyP/vbaMFysctHdNMuMkCuEYzlYzDHRk3grjY+
Up345FkZJHoTl1Fmonq9srGsBSk7tjZ/n7fYHjR6JGbrVBdcepdO2EuZHkPEt/9F
J0MkuwTJTwDJ4RT2SmO0jKxHM3Dl2KJCGZzhKsJ7drwRq74bOnqP0QB1ze9VNn52
h7bBU5aXx0Jjjx9nxUgoITcz2PGsVz5R1GkAa+nzbr4jHlTFhKYeAnStMSF8/dW0
i59x8BUg2RyCU+H5aunVbzQ7iY5XRo9lIo8owtogSIeoPI0J1OcttLY5GVEdvAlR
FCyd5C/7O218KJNifHKDADgzL+mk8bgjjOoReMJwAqC2FAGXYAvhSYcwWuKzgUD/
mfXrII5M5L/NdqGb5DKf5iUbAueIGRTj+48NGyU8HiPDSRWFOBHK+tpXwgo6Kf+E
0JEwI8y/DhSEu9PaFrMpQNr5yV7yFt8FYUWNbdDSQkV5WNOYCXPD4d91wieNsm29
oy+75EnYH/v3yFv7HU4WUA3YL/dzTvmvnS8C8XttyhCf5ufDdydVtzCSLzgLYrwH
FT1HQme9BowWIkMbfXBx7ZgXJJLTwj5kzVUwzhYJas6sKStyYf1elmglST0wcuok
QUjP24JqnCP+0h+0l7MRXC2dWfrz40iiVaTmuMNvlkPnXfTCebizfV2B9yz7EcEu
fe4rBJl3+L8ELtP6jevCdqWTyBmqkNtfUwxMKitppL39c0zemLmdWwKVWkJLpVKO
jxeWkHyo1u7AU6bZZTaueV3DXSwHeVkzUvCOIb044r2AxOwyhzlTJ2KO1Dz73x+4
uowrSYqZ1RW3uawrGFIpMtOu+41Is147eObF7DfFZwsUv0qEMXvGCzVGjwSdivMi
/oBxjvr2MHdJoZUA8MjXBBRlXyC95SuR5tD+ItXM3OHQhdJNhYSPBHoJ1tQ/8vf0
lcHW3gSzv5EG599tlyE5Xhvb3+xCuxcOtsssDKYNNtkJABWILK1GDO2d0QR9XGFE
c5TlxoIYW+8Sht5BR7wsJptphHKvGcN/4csCIL851c2Y1vDLGb2LwUau8K8u6zAy
jF2XyCMWjukIjKCbbTeBqxc22bgswWQI68cBnRm/ps5xesooidzsvyw2c1MxyUc5
5jknqVZWIDTrpmUpJelNTAGgFsl3LDtrflzMbBSFBaGXgwWMlSxcLgRu5+l/L7g0
oyxHGiEy35Jr8H/8m00eYMS3a6Eo7HDf0qnbcJCOGgmD+EMmfZoWofjUq3v/bJsB
99OfLyA4gIlN1aiUtC+5AA342/1Ok4QXalfmGeD7oY852hvnCGeiFeUCZv8TZeVs
cYLBvb7F9OMGVn+Sysb7TQV7i36m8laPFPNfk5AQ/Qu+9dbF/O7AWNNEsHxbBKLd
9FsKnVBqAudmUleuJYCLbM77pI7BDNHENOVOSV307TiTZ8+VnntKLpe0R00gSHPk
YTOwm96JLCJ6Z9cjDnUJWIl8n116i+gQRT0mHPaqnxTTU927IqsonCANvPwCl5L8
DFRF+mZ1U2ApWUzJK/MnXn+k7LKSV+VgYl6uW4WF+wswEjEWfYISR7qj0hUl4zVP
6HOKW+2BgfWOLUeaBZFF5rNESMJrWO0h+r0JoFVglE4fje8jOzYRC9O+r3zrwCNE
Ir4imKLey3uVu+VpmgrRgnFQohDEiSMw46VwfpXSljl6e+wdvtGbqPtAczpMhtxS
VaMjYFyFeY7oVlI/GhXi2EvDC7T7julBlmo9v1yd4XOGmUQHMnf/dyij/6LCt16S
X3bkAdcrmehdxv2PG7h3c7YWtuH/W8V3Szjle/vXi+1RMR03fWAh97fesjQcoyug
KhG40Ey6L02Fv75cyH+rRRsHfn1zetoWBEpEGm+RJx1miWPtJ7DVPJjgZXcvNyuN
WMNnS42TmQpv8JD3VqwG/sicX/QFyAu461WdHKnbeTNkNXjnef4Hua5+ITlAeLFE
dj8XhwPIthgla5i41fx0UipKWy6xqpAklVFHYge8fVeNgvy9HR5qd8WSsSlL5Dxh
wpqs1udwKOckbdGLhP5JmCjqgnwphI9hH805PI8aDayFKzmrT1cG8XtUrLofDmXq
rSTRmjNT0brnlWGn4gSp5vI1FMyZ3GUk32657Tf0uvXYHj9YrbTHraC2UycO8r24
4LNloujNadMQq9eFdr+g0ArtyfubXEwcO3Eo8YP3PPjs0ROIphMEaz2K2y0/ynWV
zmAL2JuuKUY6w4G/PfIw6wp6X/mwdy7+1xUzzI/uBkKSMo7S8iyahlr5UJGl4EZ5
17WBWI8YlDpxtm69q2atXpJxZg7Hdi3pkc8/f2ZzGQanDIf9suA/uPljpTsts26b
zQs/Zvv4/9f1QK6I9jpH7Ss0THXf+kUs75IkaTH+qDUNPrwC+NurGVnW1Wyzc0cJ
sLjqnIb86cs/gy61+o/d/4SrbMNY7exB2IiHWXDHRcJ8XcTXsfH6KQtr0NeG5/Ji
ghJY4SLZbtRCcutcBS67hdJ7fhhZxdSRUHys4JaznNIhxxAqSOwVS510IN3Bq04g
RP/W5ognCfciI5WBWMxrRxBN9ise+CR1GIIbA1gyjuVi72T0RvCnLQ2WOsNrKW70
y2Y8DW0rbsG1cfJZFOGJlDwitlLrGi9wdZhepSRYSDjz8uYNpJ4v32EVoP6ss3OU
J0C1L3KtUXbTgjyKsnrMaEtv+D46SXnAhbKaCu5cZqPjjIulIetaP/IXRKpa6/+P
ThPZge/FLqdPQEv/GSuJkZo6sufStg1/y5JWcsTBJbfJJ67vfRoMQQg+jm58CvTi
GBHx0bnli08jrwN7a6k8XXdG6QXmygTQs7SbZ6BbBFCvU+Sgl9n76XqZfnGUijka
G6Rd3TJgeZrapvlFVRwtw04PrOAmzC9WJy8RqmwlMmUirmfDdfYqx5QjLGfsuDIf
y/MS9cuVrB6RjMsDNyV5a21IthTZcsXK0ejzNnnB4ncqsyxITLtrHhHbkHsrj4OW
+N9OQNRBZH+gsE5mhq8Vzrteuu07msAB1gRZKhRX2Lu7J+XsSvoA71FvsboW7y92
7vZ7wMIXq4mbcGg38mH5dv6PGRGNWThrWnlzs303jKoCFZ6ruRg6JWKpZt6bMfsT
lnYJx0jJ95Bur0zJHsefrqAvvKcSJGvtNR2ZLsMRipLG2T5DkAVQQ2ELdjyVmrK3
tvqZrWosxiF4BmLd8MFYTeJC66p5R3tulu9IBbDictPD51jklOCsalX1dhU5F9N1
IDSW+jRXyTFozFcXZojAUmBZLKytHqS7TJ2e5lU6MatRIB9PmtO1Gu+KHj+7aL3P
DBDO59z1ndGSUE31tyOd2Gi60/JyVhaFWPWikT4oMAzk2MWCtOUL1dp4c8LGcMYC
iuCpgUJIr3Ahl5U6KHonbA0eZShkiuHBvRu0ztsWOMht41uJNvmpplUec/FHEg8B
HxStpGf4R465SReGASIbx0Ytsl+GtGv3u7+BtdrEawzWfifSJ0bqZpeL+V05diW4
soMcISg3GUjnW6cnd7Bi6Qhj526xW+1KipkW+4y99fHAt/T01jhUqldy21n08yTf
ctHAKaNKChIu3U982Ry64g8owuSWCnS5wy9qrqCVo2Wq7Gd9OeMrbkAaf00PrklI
NHrTRhXp7YS+SsfL58KfEwyQg9ZnH+t9PIF4xg/6UteoRkzD/dkifN/0GTRoXEss
bswH8O8Qvdi7Xf15aSN2I/vMX76vqQrJH94q6AiMcpF6KVJRod0cGCAjwEa9DaWy
rbuQNxtgKPoplwiOtThCr2QqvbCKsLxxSNGxHvJFHcxNchcx2vvh72hH1mKbsYZD
i/S/zJdY1G3YlARfD/5MF7XoUINL8cSj4QGoZYxZhg8SV8tcbrLijJ72Rzbko9dY
dOeuc0C+y9mcLLu22cOWSxDQx7yTsyOUZFBJVffIgIoKD1e6/urXGRjJuP8NBrG1
HyJ1xUTCr3u9a1g0YP3+dalo8b0p8vQoP9v0Hr0O6+LYQlxz6tkuOCh2H5qs9pdw
fzS5VlVym7RnQIFcESzJOIaQ9yPSV7QPX6staoXdRa6SD+n5QEXXGzZwMFCbDO18
6PSZb7FrZBAOVqKl16TgEcSor1FX50elhHlofYdhVYVlkq9iRl9GslZQP2LoaEfl
4EX1WoD5EY+jj36Mool6crBCmYJiDqyGsgxAq5mGoT9pN+ZMq37nUshkLvU6TgzL
zhyWqXOnkaOO4XWcuWimizb/G613MtM/0rOyExSOuPQ686OrShAZUMupeByUpUei
uoAi9YI24NN2yZbBsrI8DVW5ykgmjc+3M+phKQYX8o8sOUFCMTov+0D62XwHUbFC
nPQuCxy5ABzveJeesgLZ2jfXl93ot2mdCbSHFrRmn2RwWDHZq+YMFgPktBp/t7ji
mpJ8d8hQSD0UfH+9VspAI9U+P+O6MzDEqf/A1Y2ZXsi3KosDAe9XA34kAuvcf7K/
6kmSKwYm20Vv2AsWFhChYR9zYq6xDZtI+siHSi64EmQgYElAndBZUmM6QMn86eKW
yE72vu6wE5Vfwb8p+tltj1bGPr0fRAMILLH07tYBM30I/vYbQsiqEi/htx+9F4N1
zEUzQ6g53t3DX923Imj8s6io80jekId18n17GZk2aEgZyalik4hbjcIYS7utKTZS
pI5LKifCR8l20nzuzvxYZagChjOOs/UzdHyHczhcbcEKmJqa7rJh4nmhHlTT3z0j
zTrCaU10nQCQ4x3gD9FeisK54NuAqaT6O9mZ70AaS58crNoFy8PKeJ+ybB/+wcBV
hN48JcCdtrPRN4+1n5tkC657X0IvdvfhPs5Xpm3T/Z/LAd+HbcPCAhHZfx+h6Xnq
uG826/LB3zMZtwhdz1QE5mJk2xJ5RU3J2pNJ7nN71Abhm+b4tEZmwkVXvzDnrtTR
iI1SWXJNgokVZVQXg5VLStreJnOR5UTYnNIrP/3Le7qifcHZJGLclCDtuKZtTNyB
x4fHrHUXn60HdYofpMze1+QIvlL7uUQKVIGqA665AbbiZMLyjlMwrceuam6lkFSp
KStfhhym/GhfYUtVO60I35ACe9xfzRWUxw21HywST/g3Z7Mu/EISicIpK7AhRByl
nl8vrSTGpXJBmTTHBLtdmXImd2ENxhYmHKTxMN0BL3QuuxlFIDP9p9f2Lmxi5K1V
yIjg+/+OJIg0AHjK4D2phj9Sm7dPgjglNbkoghpkMluOggp8DigsQgAsEaKOwyf4
/c7Uz458kx2pVGdkSH36Xr/QbBfuQVVsiESOHge3PDnS8KdO1JM/DgfdZH7VXsl8
AmtSEFxWsTSYzm+6ZOf05mjAieRyzHKb46CRcHmHPB5g9Z0goiBuRMPKw+KH+UBq
iJmzTjsuIOa25UYY+F6vCp7KiT8iKWzgVtvSWCpdy5vkjWESm6WSztGLXUByt4E0
pB5nU0j3LBo4G6IKbXy/2lXbN+p9K4/QPZP558/H/RQJnxLVajzSnVc9o4Nep4si
A8p72RCg7LEWK0oxizGb6nT+x6OllG8mE/7pzqVppFcZSEIG+TqRARsrxLvytNMA
4vxPmUujvhIdzLx4LzEzN1PNZqLA7pH2S4E62jpAJbacpXhbO6WRGj8VUbxIhZ2q
XrrYfm+AKNvMQny677wgHqE/Jnr9/ALwxdUCMlJcI+P2MQSVdHZio4T1s6raO1Tp
W/zApX4ZhZUT4f1AJHr5fLCMfCRiShgDOIIOSQwrQWcykbMZ+NiPM81EAqZYgAPy
PPzmMAFIX3Tp00Twoe7rk3fO40VqwypNqa2wuRW4ASlrUhsQ4uxRWHG/ORnInZpM
C6TqEYRKvIH2yVIxjDMw1yy+/IiP/EzznLdQuFjnYJ2dlCPSZ+w1C9Nx7A+B8AJI
ycZu2+UD/JvZrFWeP4SwijUedaKVOuDr38VKXbDqvsHMN7dbMUnz5l+cKksadA7S
LQY7gpHa0Mo3hron529cdo9V3lJzaGjcIu655076e4JQ6UjJTiuP8loUZDh25QXM
8nA/jdHZaDYwJ8XwK0EjP5o+L3uMvXzoFyxLXALjrRM3SXcFKq3FGoSO+/R3/a8+
MLBsVeBh8jJ7FsWLSX5d8Vs3cw9K7Lrz2AT35v2TFamznJC0A+66DGYa+OlISTDz
/U4phwuH/G4wibFpy7EZ7VevVDdHDmcm+mzMWuimcXYpbkIxGq1psBtZFsKbvNR5
Cpw6dBzW+Ps4PBFSc5hIst6/83thdpEQ6UnHQqxQyvq1snzn5uIZeTzryN8BPURa
T7JsE1XH6hfMEp2vcVf9gMoB7TNOHVrYVmSNg4ASTEBXdcXXGwV3Jus2kI/FuaHn
/ruBbySKtE2h1ut6ypTZYtojaAfLUFqTiDQT/2DVL47B2AWYr6pn8WXMO2X6moIV
yw8JhQVemlVcfbCRiIAQX99UTjVJ8+Uu3pFisKQ0h6663zk97WCDkZYOKoOXGJXe
wpDHOWDS557aEuud4lA42PPN4mBR01pzWNs0SO3JDEY9rZ3Gmg9sWSSFL5Ip7e85
JeATuDhwc6KENb6J86cuYL4FpXYgSW4rMx4Mrvw7vXTbAzHRydTnfDUYotXa6Sdw
F+E90P8sHgOcrHshZXTgwfOkGRcYEHDfWIJp31w76IblSDkhvAiVJ2HzPCrxI1gW
bbSU7RCXgfQnwtYX/G0NrM+Oiw1gj15ihZNHJ2OK6fglZVu8YhHnVRY6l7Gqxtgs
vva/r5ONCf56ONtmW5kQ26iY/Hf4QIw6KGruSnwMur51wMMhxEURaKwlBVCAEm9r
WffbdV87ca3W5ePQgK1ODdiBWEZ+f6st2oFOsIbAXYxcuIfs4ngF0p/XDIExivn1
ymSU1U2/0WxPlxyHEJXBPu3umVp2+pTc7kYWkrXbjQzyuKv2lM5fDuQ9/o877PAu
UpJB0cVB/vtVYv3+EkMm4m1WvaASbjAHN8aY7VZbWC/XiNE1iRjFTwbQvXTvGf4f
YgEcpRq68EW2yTZv27LEgZH+OOX66FdlNbNXsvgVccWnUDOGEX6W0sqcUjdDvWlV
VEum1krTLqpjpp4snCIF5/cBVc9YF5l+jRQZpcJ7Nodtc6cnRMFCJcQ/QDtXPb3Y
OVAIYKPL1tlR1yy5h86DZULLcIzt6Je8a9n8QipgXGerG623GQWQBLUXv3Wb9zir
h3qdyOUGDWmV0/j0NspC3wtQ8mbAbUVDMGw8gPGsZlhnHy0dmqzN5Jp9I9xpecJs
UO1KM2+d+BvbLCaspVEBo7cjSo/G63XcTUx9I2ynpfht8zcG54A0R98NrenwESYe
dexhcsY6mFx/V8lRUPwqAN6nBgOTsdehryL1zf8K2G08Y2Ov66SJVmO/zpt+ahPx
4uabLOhrDDnepkWJ6+rOz2ZJu48ICp26ejx+pUQtigE7Q8n1qj07uQjh6DpZ9HJC
V4TsdWOG8h3ETvLblY7tDBvoPWbaiL+dgQyQ4gTJpe8pxcAvJdZZNWmbXFg1UfL/
2Kvn3aXYJImVIfYfClO8NxSEFih9rCFaqvDPKAywi9xcUHKS3Yi1nR/K6wvo066i
e/3Hoc1J0thInj/08FwOFsmtDWpN0zFvEt9yRsMREtFZ56c0qvmE9iXFrJcJe0Dk
Clu6rCvs/IWncwAyaPLgdx3kBlJBTnp5apPAwwY5Lmo3ScR1jwv4DC3ZiIBwivOy
ooz5JTFDWYucARpoJus5/h72RHZFYt77Qd6aufCbs/0HgYv7vJlwWerrYmAjkTBX
2tKntHDKzdAF5Ej2VBTVicSttn/9MUtvn1H/IT+9YPUgh3+IUq8tc2M4/KJHsH1v
mSMbMulS/7YsftzbO5zmtbePpQwrOLvf2gO6sN0YmJ5BU9/O66qbfeULp0cxOyif
pzKNY46EallamzFaoDxxkNYlYdxjr+OvXdsJkBzVs1NmBBIJi21n3GNNWDoXXge/
aEOZIfGsLwkpOysG6ImA+Tf7i8xR3K9aaK29S3FEX7tKOemS9HyB83SpiZTYgjFK
2na1M4lVX/8k9G0jdshk2WCqlejQMkgo7aN3nhlTyDC+ztmHhHO7uhIflAjYTV61
kItozs8LWEoAFV7V4pfY49cKvKpPAhxKG1VZuqHM/x1qqpFIeic506UBIQENcp0I
gpjylFpQ9I5jInmfEGR9YNPq127vxYF0BfX8/cNxDty5ChCtda3fUHeEsLYxpszc
AYGPwbF3SwtqRCqMDLcgiig7Y2cjEWrYI3gr96Y+Wigj+AHw+E7xo7NNNHiwHgmr
84/ZvP93DEqRAE05CFTrdzaz++CR5a74ooSCwp0+l0aWvvb/Wxwg4/PoDBX110ec
Xr09nPG4SVws3334zrI1nfIq/rnLXFoD31lsAuvfcrUoxgdqbAfGdyAMzUNY+TvA
b5u2e3j+0fmiEVV9Hr6lY6CDU/ef6aw4LhmOED6R2Y0t1TqHiwbWg+0QguM9ifdv
/DRxAqKEU+sqXk4YqK/9v+BC3S5DnygQGNmgn6iMGHTTnkJ+Uvjv+Pem4y2p/jGH
7S35T23w5VKrqFGFcIX4hhMAPFssHjgfou9/Oq/i15/bFpA8SRLnfmckyXbedLaN
OtmEyglMFEgE056Ig1njg4tJkfVogzmHgoJplpjwSEMdd9nXOQCX+mU3FUn49iAU
WX/w2mnxR/nXUPKte/BO3VVq5LiQraMUFVd8h6khleOvRGF0tZYmLKMaTOS1dNFj
n9WY90tyroZXMnbWvr9tTPPdfBEm6gibUDAYcKbos9APtfhrBEBn14WZM5oJuUIf
dDdirS9QoqaA44jLSVdgOiybFJliA3TbmpnRtIiBzTP9CsIxoBHhbJVgPrxwpxxg
Aw7v8he7NBzRfilBMAXHaq+27FVLZHFZqvLaJVK6qfrKb20hYu1rxwSHkJR7ZXFk
kfsdF7IVEKzOat/o89fVj1ZoS6DgnJWXdI3vzPs8GPKPyTwiLQDG8M8K6G9J0R91
oSmyIo5y/57Dis72nHEAnZbUYhZEEgDTMgP+ypkwDPA5DRvyXocqGXuWMDxDCCy4
mXNL+3CHLqghBY5KkiF44eBm8ICDtsfji4NLIlLnLpyrKb91n8DTwmX7nOEAquhL
MKmFFSirR/FwjC9bHJNfs1G+4tc1EgxvOn47QfV6C3hpctjxnhHxlTCWWCAKipJK
ms1LTQ7gmHH63PJYHahDm7O63eLpYImQrFia1qRZ09ZDvQCtHjRSUVtFLDFuedgn
H+f2/r9/l0iwRGkCkb6hsvtAki89J5jfgutXjore+JLk5Erz7aUkSQKb/wZTHi3/
dR8sqiZivwXOxXfZ8C9lt0sFxf8r/NLvF3Qqg0mqOp8T6YE6a7NPlRYH2GCQIXJg
/o9HtQ1aLvnB44hVfhFuclqC3T2yGESpr3XlZTojZT1/BvjimfA76SYHH56u3Ibx
5TlL2nlDVyl/SdoXWyJAHkYJOfTkrlNw4dCFMIq/cLD1n5IRG9SAjpXGt3N+ZRsO
vzvPc5OBpRJe0onM4xdZ+WsAoJ1JnHwhENj4PIkwYsfX8Lka0sQK9GLSzesC6Lmd
Rl/0SbOdIcQy7/BoDgAEc9d8XTw2qRmoUzAsooTAc8juPrIAsnDaQkSiXv29DssX
e/P/KD/mdpDToUk1+ZLHuY9NfHNiRpjwXYMno+ei03hfOiGU1z9HI4YITWlUHj6q
3+BoDscfnQLsu0eRnT4eZMjk7R6s99kYbvgRFOA8RgJBblgiAsX1Ep9nMlXvhWlo
u7zpGe0V0TM0ZMjGnTWXDDXwP15NrZLTMKP5IBkXoRF1djIXJomhe6ZXwOqOmT67
Tths6Fah51TtDeoaVo9aBV8QvAWPGmav23P3XWIOYsZnWwE4B+tVWMa/AmHP479S
V78pyHTJWU879jNWXV9hSTQNfMePBeSHgcs4R4y6O7Au8jXp7tyA0opuLZUdtP31
EO3FmAoXQowBR0+6Qdw6ATW24A/wnjqzNLdlZuBTPROS/gGilVzIAPZX/n2n3KHo
EZW5UWVqXuiXz3KPTMORpz1mQKwQ6yuIW0rWSUs2RYR0cw03NwL6B2fA/BqUs1xf
ZEXzi2fFhN0UAYdGPX7UqmGj5Y60m9Ocr041SrBGLJBc+wqGZnSHZmZ+epnltV8I
mwpums4P3/kOhQ57fgajp+iZTmZzYh/01mlLZ3a63qZQuvTyyqCJJEGzFZtVQiBR
OGaWWv4lJCpx3TNCZ+skbPVpv9A/N2uqa7K2f8tYCYbbzf70/1tUfa4epYBXBqCx
GoeMNm/jnLGAUxWT9oewG6FrL8HDessvIppY5GI8Qom6hp19iByAD2XvG9Gi9zhv
/MkC1k1kdb5Jt5aZ/e7BPOaj3AOgzs52V9cdXBXGKxdDP6/X1j8QWel8lv0fEJgR
bYlgjUzZeL1a/+1Ds2ikCMBxrdABkUSW+TSvPkyeI3S5jcPfrCrQ340aPaoj3ZxH
JzqjC0ksJE9P7cdxOuYCaYkGKzr6+HktCHwMf45CL7YMQgE18EnFEyEHi60PGyi5
+2sApULUsyxeGc/N+ECsoauyiZ7EwCtbvj7amXemnVElGi+s7A1aEkwX3gJjlVYZ
WaGdyCfR7Z2ks2qsQg9a22WYoYL2r/wyFnDGsHVzQ0B9yAIoaVMxqnTWXEmLsd0s
Ea0SU+feno2tETnHT6oL37aPAhi3+wEnBuH2iJ5P+fb7d1qnVrgDKznCqt6kLCJx
jiFcWGojv0yXhWmZw/bm87TlYwbIdo94LiDn4dplYMHlDre/qmhxE0k8l6bMbbzc
yO35NKjZgX6pumxqBQLWfYpGuJGzRbZGnlLyYx3jFrlqlwxkqnKueVLnDGnQ8Fq5
Mo7TMyUcYx49NT5F5iMtb8mTo/e16q9BU8nVnqBaFXaKin6x5WJFDuNm8dTJApul
j9MC8jZZ7j2arV6qj6qef5a+aaDIa0+l1qvEImTPiy88JtAShcp9S0U37pEZomCO
kIQBLkbyvQWbXLEq2zkIwRLKxiylAjCqUr+X552/eo3veeJTFoN6MB6DAubOvshU
FIigl8s4JFmUGf28RWlwE/DsT9fmGxOwvUnNpl8Zd7J5pVVem5mJWELivCZcF9pd
+Jhl8Tt3ZAkIWBpg0wxfz8Fbq7z3V9DNsXGMIF4e4cx41Cza6yIcaypL98KkXRBS
G5aukTTen8cvPqb6G2b0uTuaz3FYIVhLB1MECGHq46j/BLXURRUNXfhB0v6n36Ub
ODoRxuLWTMaEienwUp1VJhw0cpfeTaXVQkRGYF1Z83urKmT/YhBZznSKuCNsXPDa
aNxWn21DG4amD0F7JFbFJlvLY4urOi4BkmI+wzzHPy/slEPEXLra9598si96d+bC
EkhDNOXhd3XgKPwds5CWT3g/nQeCiFJ56DYSXXRMYu90qXuaPra8Ux0cvB/Echa+
++gTbj1ugGRJgpH23KVcFG2caNBtaewQC62y8MUAAeKsnphzGO9dCB+y1Jft0MKm
P8jRi/Bpag9wKnACqBt/mAmHunVO/lMCbqnCaylmtxCypuIBrV4vbSnnUMA+U2B/
DeXW4oEGmS6eHAY0GIUTUGRQP4RLUHC1kby8IpGvvZraLaUeUmWXlvfwr285ORus
VhjldlUkP4X3fDbqKE792b9Ds8FaSW1UYEJxJ3DR4dWR5tANBKHc1qMu0uaPR2b4
ov1HPlaF7gw2OrnP5XUua0ictf8J+FjiOryYB+28qt9DB6YGCO/c3CTvQW9LsvVv
BuFBHOCqOJTGO/DcsnbnF/EWE52JZ8NF5Lq119uuPyg1JBbIBBJC6czpOuf83Rpe
irzVQP3Jg2js+z0j5iHTgHZHedNVhlPuvjyZ/bLZPuVKegPiAugLN0CyGmzDM73R
IgmCCs++DfMJc4wN+k8R/895/6ikxnQDQWhdzu1LUiA7D9QgbMpyLkoJm9E1pidN
vLepemJMEYQhe3hpwJfvusdMafSK4iEOfJqFS4UfULEQ2csRbTV0d+HBFGlcByJK
JvVhOOuQHB9/PWF0qQo/4xIi+eC2SkozvfwaaLSrOifaqMbLxEhLDT66/qHO2W5P
TpodHWKtYMaT5bkAvwb8PJptDit14M/oSC8xFFGm9UfCfiWtaDyPZDXB/uGnacJm
Cz1ETsZQHkkDEeKcUkzV5rN0DXUDch4SyCSwKXEWEQYlOKJlkdeuaWINsNXVUwbQ
rAb/JpJRyjHnmh9WU3USaY/HAPL76gNFC9nOaP6aqfW5uRN8va8Kz0DfGcYc5WBv
hFDu+x4ZZ2SUTEHaOTaGc+eypVboW3ktlw1ij/r8VLOXtj7uGjBOkzzWNVmuyS0k
NTMDp4CHqhm15QAkZmFss6/HKCfeTXr9XODaRtzBgG+nJarTOrxIvtVz329idvCa
yPRdyDomJ/sZpEj1HsEtS9ufqBldurPKt2f0/DzYt//ZYgSlctHAdcXuuJzC0C5u
sDpItAmSAOCex8Smio6YmZZdXaENTBELDFSAyCuMrASHPA7K6I59KqzbxHanP8pt
6pHc2TDcMbc2xSg+axRfnyyiHZDXcqD7tKFfV3G76omBGYPITLOb2zk4ZxCTAxd8
OJwtH/3HNL34+2lr8TSD/VLEQsu+hVt66ZJOuTWyA7cHeoAVNU1pX1nwWQj50d3M
B2dv34MfdMoTfhpRLCEFmySo39UUFavfyvLRY/I0goxTwvY8uvPhlyiyHS1MfRvU
DSiej1C8Dn9roa53XwiF2WhA4Lz4k6dnE4feR/D78o/3LXUEOG8wPi4NR0nI4wLA
tVPSkBQXT/NXXLN/p/j7o+6FqxFV3eJACaz3XszeasjNIJxWvz0c6PFzN5ORpVXX
SoB6/GO+8QnCoddmWZqjJa0mXPwGJzW7S4sgzQH75eIha5yG3mGKQOP4umNtpvjN
uBlBpQrIon4DYyOUGOBHL97mW05NI+okj2cYZBxXqfvogGO5XSP525sHKSrAWw7m
JFMJCP9TRQEo13QnHHqHNhWjWrrTXys+qwgddx8pPhXMQh7pLqniHQsJaqjZFwJA
LcmqHi6lQuUqv7cJ1O0dyEj7fI8A6FqWNeTwd2IbW9K8kY/hr0uJhH8+obp0v893
k+aZ0dUdjCnAkw0L0pkdPEPYWrn6JjndWFRqqVXMsNihrbno97fd7Wvapt0l+Mvw
oNbVq0YN1idDjNyJ9FD5MQ9GCvFLB0fE5FWLsOjOs4/Oe88ZZtYS7/xC9S6DG2JD
ucrCNS/Blz6pTRYZ+47Ch1sOXxWrN025LvkPDJ/szcSeGTeFRwr5s/9lheeBowWe
M2qw/0fMUF3ZESUOFyYxD2hol4i2Y/fRFdNz2XaZaZ6WseDjL3CBoyyfnBX0Hury
nVmdvJxtbnddBKXHTep0WQqx1J7rhyCjPLikOokJKkISVzpTxJwKb2JrPA3gaPZA
VMaL+BhOvyr/v68VOqHt9APOTeyxzwwpILRbK5yv+rgFQMO3JmB3G24joiA1R+ly
czTzSUzS21kTAE0Pr2NlHpVIE0wgnqA5iV1596LBHDpFh+fSOiQa02owVlux6Nqt
IFmqHuaovX7ArD/rhrDRZq8/OBcblIvO0SWf9GRXTTT1BeWkk4ZK8lGGuiQjv/ul
jVoxx32/OxnRjAWK6VMtZ0/Fb51nE6M8JZAuEoprO3vezv7acTspP4c/Q/799jMK
fvrJKtpJiLuT9Ov2b0V+0oZ61NtXK8kGYs14C4JHqJVhi+PxU5DkqNST9WEJW9Tj
D1xI7oYzPcuAcPDNUYkjdEjK3ll+e8adblsp51FwYqoQYxAMnI3i9cP6T4yTU50V
+lJiELAoOtDNNbdAvIVLt+EeX8BIaxqtcqnfb2BMT1EAqX1zL8m6LQEPeLH8m2GM
EAdzHMJRgAwrhdhy38fDauMG/YOSIGAxcZRh0LkJlvGB8pH4RKq1xEtQf0uYHmwX
caCgnHQ3NOijOhn1NgQNLQHOo6CXBcRSLA3PuFtBDICufmzof6m8C0sIL1hRRfuQ
8a32HADtsStacMyqp/qp86q3AFsBbccVv4gnMNtkQq/gEm8lKp9YKYbPeXqiWeS7
+Q5BwidF5SXBb2rovXCmIBNkQWL4hqFL9G4i3wD8Crnpyf77P2fJDn+y0cq9rba8
TzpD/8spj8YBQ0PjWeW4jL1+sJaZeiJGr46//6diEWi+xfMqxXv0hxSgY47fK5/o
ZIKga6A0kpQ6OErlccLafftxGcg7pALarhd16OYXvA3jL3NFTrWpblLKTUx06SmF
OtEJtgPat0yfywMVLsC+AHYjvKvM32QSyHtccwXQ3mJyVOFpXIAr3qodY4S9E5e8
PrxYAak/bMAZbCJSH99z0Te/vxPFjw4yb5/OV8HWyRe19hp/ohuqRSKSyVJC9mDK
xyz80ud97BRGmHTlyYIhB7ceDC+2Yrn2utMajSUuj3yWK8w55fz5mcHQ6Gwch3+8
wrp3WLjF06PXwqaNBGEu0k/qdd0udXy96ydPvZLuS4LB0/Y3Wce5nlk8n3QqpmVp
rEww7oS6GQdmg9fB0C+3yfNik10bvQzyDOdvhXPWqkS1t4V5E0UImncEcpNYhVty
01iX4eNyqJEgak+VWqY0BW+SXFNr/xZU/oh+OxF4y3WzxPgxCIg6XlFGokb4FgdR
zG0NJnkuYSl0QjX+dYQwoPsbr0pjKuwFvAqx/lKPy/u6ez19RacpXYtYNSCXvJTQ
+5sddhMXFL1vNu452KOiw0wXlbGnexnVFYUGYcxHzpGIapKgEHy5FE1rIFrCJFgJ
0nHpVIxzVHkQjqRWATSUmzRGnTAMUgvOm/393bSemcOiujYzpd3qPLHsrP8XkG8i
9NM2OjclBJJFiqJaSVDeV0LVlvEr1LWT4HwAjttPt6v9I42mxad+3ISLmF7lVmro
wzz+jaHpkbXCrMPVjS/OeDfGrsa14VjdFT/zt9l0qMBBBwyxixOoIGSa+Md125Mw
YLdnntQ19B9xh0LldQj1xIrHOz67p5OSZjFl3DJvLtzaxo/BkKV3+SpWU0dQGQWm
uTa+40yXNcWtgYMoSt1ffReXxXNB7jlc636RHvtLNquvLLIcuvVKT8HlfjUNax3G
qk89BZSTiVS4eoMnp+tisYwuL8obEXGE9BvI/YsQShZGUj//vtpof4HFKc2U+Ml5
Ru8LCftU3mDR3OSWbxMoAOqw6uoRb6CT47DB9mAZtshG1ZkD8rrarE6decSklYPM
3vrny9wlqO0KSynXOh3HeM9KtH5TPqK38oq1URY54WHN0jwhej+/kTkNmVrHFDrI
WbWNj/0ISmv8OT9LN7h/6AtiCgWT2zlWAqwVbfrRSYe6xT5GgcIqAEoP7u5XXf75
LyfEWTYLMDvYMrQKg/IikmWO+FJ5trfC5ZGe46ZEUpfUnc/mFTQhVse51ao2MgJW
tvrRG/abhQ+x6OfBuDso3rxuJLAsHlgdgp2KJmMlTEcnBJj36IonLFyDIDUoJe9m
51deLtU9+Sa3sNXee+lqaccVG68udfwyk8xMFZZpaqRLLUCZIfJAkOFzf+QxCse8
1oVMc+hRLpL2r9vld942c+4KNZ1lLBOVuurGaco9zVNi5waZKZsN3Ev5iRXEP/CM
ti+QsO7N74ISQimKFmJdyHSGvIHR4pShuKugfxZlLT6hnZVVvZKf0S6kOuOE68Gp
lQmakIXl5QtOLH3Cn069F3KjlgjjEWioQx9i4ozbRrGR2cqdoSw+aw5uO0l+pHWR
FGpfrP/fKbTP5NpoiJ6OLHSBy2jOPtWDAVCsNMTkauNeHgNkaHInFD4rRa3J4Iuk
c4yKkP4vqKiV0Sw72xG2VLb1rdtwBlKQKiFKA4mODUOWqtIYdsbme1lGvwjYIvTM
S3nC76zhoTd2Lyvwy1oY9jv0s0p8E7OzwU0+1rFHZmZxm2hWNy/4pmB7z7yrX9MR
3h8f5FUec4zjuAxgJIo+7nx6hfpfgLI5u+gDinAae3sHXEj2WRPOCKGDotNFypEQ
+Mc0X4oV3Ypfdg3w1cco3KLNn2O80M2BnvaM+4W+ntTzpBsXXXJbJEhp/oCw+xRk
NFQIIO53W/OQn9mlVIR7KiYsNOllIc9zffpulBWV3oRUTjhaSFsnTJhkc0ne6P0U
usF7tjfljfELo1+f1/21kHdYefdH+zJ4eaJGVEayWmoLsNZiKnBlFpTK+y9Iu1bY
khyPIwpWTSHOJRCrXEjOQ9wRKtmVScSwBbM4nI0AmcoGvj/2TWMWe93aHJGDC/ec
vxrGFgMlL8PzIaoJcsdfOiNCIXCAPjkakRn0StlCHaFeEItc5HmyzlzdnNXmFv5g
kQZGPmZM/E384lARxo2rDYQebuwsxemHjRskPe6xacatwjR11AlMSd4XfC9OFXMY
2R5rQpAnEMtNxi6SDRKxPQ+u/E5wxd/rR4nL5tPxUo5OZGrIb1oKUD7ONZavNdna
566fmdmr28kCX/k+pUthhTnSDE0WutR1NdbD1mZYfrPbK67L+gliSEuqvbXJ3/BO
AKVyTWtqhMhlDpno8jRue4e9CmxO7FDzqwqxgZmjYL0XyW2D35rDrn1mYEH3awGh
UNJHQUPuERB5YpLcIhcwJFt7GURIVfKR8sImWUo0yYtmaXbI1Er5JdZ6HTmCT4/v
lLtcAdlVIOKx03XXL9f2BOG12sxjwKDCdqureLeiuXAeWbsDYGWtXpGXfKElTmpw
hgYpc29sY/RkpmLbV5v5uuWQ8XSviTPMYoCKpF8n3Z1E4zhMi3FJ32ZiGjrzY8R5
DTqlOrSb4dPNBuY3UVX2K9luEIGbzdqzIh+5vsb8lojRnIVvz9EuwIQsfC/hLDui
zVUn/i/0UC+QKERJT59KC5k0bJKdhVphlZOOY3juK2RSVXxZimBhVCD/ItMbjf7X
zXf06KB6fxMLEa7rGcKBaxh6BAHoa996M5nRtMywqaPX8LoQ9A+CnZZUEFibaFUr
kxBB4hRnoKc8JdIH7DtFVrJYC0URlLY5iYpg27vieWsBF27J/QbJv6Al1y8shuDu
vqE1bxBRLeYjFZCxHVZerAVARq717vY7cSeHeWiV3s+bk47uKJzq9I1RcXhy1Y4y
zUBM6sFtKSa/sFZt/irioFCwfgLnz0VcuMLwJRGxzEpSiUaeDHpP3OZPfFMW6buA
JHJwYIEP/xCpb7qSDWFVVMVtaMdseZDs3b+bKJBM/XpFgnSr+DioYYZCb94Zo4IJ
29qXe4t5PYwSrPPe+RfFpOACj47ttMttpXsHIvnWogqcWDpxAejLD373PPTgWqlC
OIr8T+nCwgf4K/Hha42LMeeUOA3yQsQyMKsnXYPWv8xjcMFgWP/2R0KSP9KO4LlS
tkaiRCHl3bIA5/RFQgpWRhAwVdYDz8MUXtiS6fT8MfSp9koB+Kq0PV+IbUS8iggR
/EpwQZKOoQ7e3SXppcze6LOBUpUYdtWVpvY0EbAPoehpbjiXbwBfYhnQV7LVLfO4
Deb3YY5wuss9MBKxpplxS7NlncTO6a2/kHcaL9GHPi5uat3RKXCMPcyNxJ2hWvSy
vH9NOGKEbilDPpQfPmH1D1+b+M3ZEvgBpYmrMm0Nf6ejbDG0CCvhL0s+7wdQPiWq
naOCxWch5tqO/TI5HkqQB5CSQA4jcIn++ovGF/486em1TkFJNKl0fUHHFn5CWlOm
UjF/MYalQjtdRAWbvIW+J29Xp5DeFZLtyAOASmbQcKADPmm4IDAIAci4r5gPiYZv
jd+N6NWQ8nW6H6qfa8UKp1aDZeyULhxNntjmXlv/43zqLNs7vF5+BmbLQgJy3AX6
nD+AHyk+PxVHoZByxqdeXdfdz0yLLLubnIGSBcxyrpHZnsZqZf0pgYGRrSJhKg+/
6mhGdU5HRE4eOpIZv6aVvXtazfNTdjQMEewERf8kufgApP9NGx+USLAUtQbvki4/
di4+pSJMr4MMwPpa2FzQQyMBbCI7Kv8rP6Ce5KeNTM4HeVC8VQpe15ctZ6Grkyaj
VIDH+ZC5qQzfxIA0qD9BY1LCal6NlRFdELNuVy3Jw5DgLQQoD4Vt9ozhC3aofQ/R
xU+DmMhCixaa9HcR5XBlizJ9PFFb8nb+M+hBFb7iKHkun2eWB/Mai8tXiZH1sVLr
L4viS3JIzTKJErmKF7h3ONHx5G0xeDdnF6IbWfaPg2ND2x747xR8/JjTHiVMqeB1
GrYLbD80k8lC/4XCj5Xt0EOGnh/rugaCaoXuZyZL9yuKbxUHMNYqpIVcxe03tsT3
hEqMSWyjeHMKRCdXz34WyJCmlo7ay5waZ0I86/ttkCMD/Y1pKh+tev++kJsHENHj
6+P8/p0uynP3wMgPQSyAJB9kh9lK46TEqWSRkaZ2kpu9jzsv+DL6OxDhIsgCJiDI
a8jeIenr3/5tnA9w2Gykd3kuKnzb8ohKhGGkPjJb+LkxZo3x6Zxm8ppaAQIhY9rJ
5YyPlZQy8qlnKyhdc5HltSlqmv7Jd8CS0ct5HBqqcS0lpzV9gUkVwwIVtNpx8rgV
hIjQpuX66OWwC7vWeUjQFr54C+KapcJTCCC6aYtwi+Avft0VNOGIbzej9c5jPT5q
azK3u1NNwuNSJ5bNDnlIvPeMYe623Cyk65HEfPjYNW322p/bfk7/34FnZ7pwVmEd
yOSWQxCnp5ej3HlDxAmNeTYyQR5IsBeIvAn0P+lUU9nD1roZHQimxap5RUa/gpUS
wRpMRkaIML4BvEUs07xsrJD+niviIxfw6RJu1DqMrP/utagg96EoYa5NQ8aBAIX0
O1eo7VG/Fbk7VN++lz5bIsJ7IheSi8oSTXc2POtBflj+XYQgvLea5tKTqwQC+a1l
o10uFRH/LNGr9JNbvf14kEz4BUJST1D1yk3O5CvYxfjHRGtKJauX03UOj8eMaH8q
YzvzWFHD33MtcNLSS/2YicJim1PjzwI0r7ekwmK8n/K16jMhc4gdHd3WFm2ljkx7
Oh6ng7dvKl5f/jVUaTzYJJaEDtB1y0erfKY7bcgaHEi1CDQLWlDcjRX/unk6SAoa
tHbnbktm2iV5sk1ceRd8SuCYH6YKJe/7o9BCSd7fghbSwk/jUOd6AlTctz30Klji
qsA8QBSmkSk7R0XddQ7N1lYyunlpQfr+2ahkCSXxn3flHEG7j208MCO9n09SQ5K1
/fTRvvl6+iXsKFueLQAYJPZezaim+3GvajOJXS0PL2NU07ihB7BtvIOwWf5ldzMT
seLZNK/Zoz4DyDCpFtjX/U+T73O25Xf0yP1AoJ+er0tuWrt/NEbd52Opznu6dTmV
gzVyyuC1u39wH/EyMKJNdsN4IUlaNo7fXa82C16CKr7sIT6cULnpTyjJUB/zEdpW
/88zgR9niR4Q/PFmdO0xIq75RjpPDyNSfS+kRYIldUmlpaoFqF6Cn4E+yBc+ccft
WvHvK6uSTfX5yTKCsL3DuLyFzrVNwyzRAZ7fVD2NUklGZqY/HdNdTrR8I6QwvYn6
xDGXGpeorqsCJpOzTfGg7Og8TLQxXTyBlASBUvwwsKK1O6L2wzgV0XhGbxSZoPao
A2SCB0dif6fEtoRmM3JyhvwDZXVNVWqKc7KLtSk81TWUImGOt29TlJdWva6STicW
BDYeO6usVCIYndEBV7Zn6apl5ZJgItaRabG1qgHepCYeRGFx8KDD5bcFfvoGrPeB
11gquH/n3O7nahOCSwMeQQx/+Q3Cu5hf+zYwOjaZu92mgzQntltqms3nzcVfj85H
MEHhOfQbt4kEXlKUFeGfaXP5b4p12StJXs9O9rDgcNFnj51Rlc3CkY2tKpyadxfg
gurEkUtceX2+9IaMiOwjqFjIG7qWsyecwRmOSHHSYSqfXqK3ut2h6WpRgV9jZ6Mo
PsCm1k8gG06qCvX3yxy2Yhc49l++S1Y0/9vSrSvhry9M67uvmge2QF6hU6ktVrUK
C3K+mMdnK4HgxqK//jgWba95cpI5MztmEShEK/9UhQ0Yk+RRO7os9H0INI0cvV5m
wzjgXFi4u7Njf74MesQdhrkwbmgN7WCphWsrPDAa73O6nDOd4CI+dxElaVbxvJ4X
zQwh624Wd8rWIknIWWUFW9AYPWXjTPODNa8g6cyrlzeTVW1CgiAo5jgclJt6nXCe
4A22NblmZnjWOd8MoVLaGp+QEJThi8fIGFlQk5TO16LZN3wpRYCr7PosA7WkB3yQ
3l5XnlcQUyOs19G5UMN+48hmQuVQsRGgrj+MVEWCa5YnaRE2VRCpFMvVQJ3jxNzQ
hxq1fp+ZuN0D75a/iWVzok9V508JUn+5xp2X0v+79F3GDiPk0p68CHvWtmrBaGDi
Ihv82m14/mqCtVbAWJqHbT1BcOSBZKBtREBMGvk3sGUHpuA/9W8bnlO9HcNR7+K9
oaO4sWJYrKIaAnbgKWKhJR/RA+CjDh0NlznFqeLzKpIzLvJg/3waVDE+6kh348iu
MRJhHsfUTCSaTEjJCgufJgbIxsGKK9frOdgA96I1p/ZzGp+nyBvaBUzPl2GrW/38
gR8UXDFcn2RzOlsJl3cgIhcTE06qW70ghUHRMjcmoqDC9i0uIn9hR8iAtToyGZT3
Hi7v1juyzyRyrnOOVFto4ryfnx3VhE/bBvyfNqmcVgR2+NldjqUcIYrluosGF5kx
j1ScvGapa0FV6dGDEmjW5pIilBWvOUbzYrph8CwSEdfz+q5YrrB7Byf3T/6BLZOF
x9b35iwYCnaN1OgvVuoN45HKGBS61WDiBevBUNjwKt8S1ew34DDdLrOhEXmdQ4Qa
Gq5cp3K9P2ava6+YvhIU1PsETFhxpbzmiYTOUFDNNDtx97B7UL3vpbyiP0HFH4rI
Ag9VM8DXG7yKIPun4vW3F5/5i08HsB9EbiAYpLrswPE3V1s5Ioz64rgjLbYNUfRu
+EY5ExVxgnq9wFb6mLwyLn+ijzhyYVrvbCKBwwxxgToVQPeeRxiVZ8+cUuCVT3U1
MpSYp69bA9cBW8KhDTMePppOPl/9gm2R6n9ZoEvCF/d54XJZavex599H8XWwTl/P
mxWYhXS9Tdh+hqAOPmbiWJ//XVQ8h0GTTilhVnuMr8uMTMnCNiq9pnPADMz4D1OP
6yE4D7cyy2DVR8BPwYtU9DTLV+Gp8kzjw+EVaOvMFdQRhaDPPd/cabpjes7FP+Dt
Hexp3FGCprTdJbPUkH+cFvU9ihd0T1h3cpeXu0polCUyTF68JPH10AqIBNRvug/x
x2dJd4iKbfmCeAinC5ZhmBh5HjuA10SnosozSR//PKXxcru0NgGKSqmdWa1QgsIv
/OiWxm6YIl/YXY2YZzscpiqe4NPiyYSBoK3qu45XmCwqJYuN1GJTZCQ1jfrggyFO
S3KAPBQkdgwYyd5SY/ECaJRrX5sns7lYQ9iWoaTSienM6lru2J3JCW5Bb7VGNklA
yVNGtnIHPIjXs54ZZhpGj7esTcUQMxooI9FkNqXqWOZ3Z6pCmdUDGg4a2Lcz65Dc
mbE9H5W0Vks5G+VqkbJ7LlqxWcjb9rhCed1RsCpEsp09MYmtTpSMYBDakvfmf4Hq
FHmisDN3HYu9uOPeRVtm4v5f3heAuTlk7kMz59XiFKi3ZuxonVED03ZB6hHylzpZ
IlmWZKnAg/0TmUHVgbClimS4vlVP8LyeI75HIb9omgCIAGKzm7/TBKqRf6jltHro
ImrOOtUGgoBlNlQ7Vf16+sRb3qmhA9pkPgiSUaGtqGstC0RhnFcraY//IpFU+Em2
d+IRWo3/1TC9uXAvmbtrMIiuSxHJloMihQnX6yc4i9+GgNGG4eCCCWas+PCwQBry
yXjPZZOvrxNMy1j6VVv+grM6ZfiKLcyr5yHV1OVoyZSpn5cUbAFpxKh5+xJ+Idwu
MDSKWziKSE1lQmVD3iTypYVZOO6o5iZm7G9lC1nvHXBCZrpeTbMO9AT3prt7EpJS
b0fmWWiBOpENrnqpKKfvtl/Ykn1hUsrpD2w+ES9kbJOBV6OgINhcMkkWc0FGaR6P
zKcioVaawpGwhhg4wkwQ3RcII2a+OooQ2c6qDZBnMykMAQgEF4uViFs6IPLTmV8x
XDihCn9mag67WMkdms/rnSqEzcIHvgPsrAufXm7HSwDgKIs1fN6tWrW+pOJX5uij
OqrKHnz4felMIOm368F8PNuHVuJpLNs0R/ugW+XhCFGLGCYimMypvDKnILAhrxJd
Kb6aNSErzfwttdMQD8ZZ4rRE6usLLMCB9XnBiPDCZnU2L9t+AC7zCVmNFKP5zpDJ
0GOT5XLK/ZgapUCq9JtXIyKw9uKbCrcVM7YGH1EA5w8sbd+qCOX2GIEkGlA2Rxdq
Q6bjVaUW5iZdCsIzUKflrc3W2gWLxorNZKA3DS7UAdHpW7N5Sx6X/AZToQj3x4iD
whvv7OmNUwHm2OFUhGao0kSuMslras4Od2kNO5Nq+uskhEzguQXD7thQhs2ZFqp+
90bBMsLKTkzhKqSjYV0Wn/Zw1BSaZueRDHZ2kpYb/rp6+CU9TjD2lsYzGU45GDRr
nFUsFU8UZQ3tAgGhYYouR3r8Mc0ys9Hd9lzfkH2Eojicy7tAV/MhGQ/TX3b1h0Z2
Yz+RQYQJbCXMDU58P8clVgiXQ85J3bDLqmwDHZ1jNo6u1UOiOAVpD2ERE8uan5SM
Uox45Oq0rLsmUk+6o4zS5p6DlLJddTCmbZDEv4dYta4V7rDn+wINO6nKLerzLNAe
bAwrBX6S+zxrq4/PkC7ey+jhc13qIayBFXrun04e8cOThpPWKoXDqz+oTCnvZv6p
tv8lTi4nSlhxmyumuCUoXL/4+mTJOVctW2itC2Bm1cYc8O4tpps+0XtjwqKh//+A
JfZnFNrLyyXdfdoXJuBDmSeaZe85nAdy8CPRGo4VJTDdiNtgn1/ZdU0kR4j8uwYB
unk0Y0GatHptbySA4YUnvPpouvD/ywH6AAXNIJ02ZFdb/jGFTabYkOb68dZbXqM1
MbAm9Lz6nhUOl/j1QExGDDU7fknGnMtYb67hTwEhjiAkgWRUKYbpn2e9iZNI0lTi
cI4BHugk4rQZk509ESihCDZieilEbgEzNBPYs125fLmdAIsRDAsUjWuEcsfwH88H
2FVk7cTXk1wekNraxvee41EhjYdMz4A7wyKgb7g8XVZ2VMlE1ZAOv3/CMArgj9oU
2z2wBgIMZEUzrbwvgsUMs3k+M1fgV3YVT15l7B8i4lAgW0vTys6i74GHKfAs2SjD
Yfhbau4a3CXUIf7ldJMdCXyUXS4GGgNqOSAfPwDQDdKfNJBQA/2NFKmvmF2R7yxP
Vh8l2QuTaXd1BrZDWf8YZaVoVgIqeadnieJsFBfbJtIbD8rkEsCze3TLpbKAocjv
16VM4oGRQ161FVSaBdZaZtf0ZFNJ1dct9+C56v/Npc00kEbXp7FTFxKAytmh+DGT
rVlw8+B9tuDvSbbcnfdTDo+/ME46bR86OWpHKxkmDYvVz2pUErmh51tcwlCi25d0
ilxRIHgtealitMXZud8HQaDdc/u0CizeUNOmhfqAbJPBYka/2sVzMMT0ozPPgKkE
4kNgOXODXkHJyw9/pUqsLt1ZGd/Dux8ohiiB3EKZ077tODWB7/i2SheHxc4B+arD
ZKXv8Mw/6ZkIVP0lhcxAfT6YNq7bn0qPEy7GIBgm0zh3oIjzc2GEQGLEMDHCUbUb
XOJ73sVfG4KqzhEgQXVMibWZ7Rly4MTkYNZSddU4aHNRvBuIW+GpdJlBoC0hF4bc
RimsXpC+eJ7zhjR/a9XWZ8y7jyVjK/DgomQW/PeC05X21oaqSROEw9kiQ9HvGNxG
3qZFVnDOKRYxVNQcp/Ex5d0ak7Zu0xBqM/oBWgC3W1tQMs/Zc8mCBRw+eIW+IqJU
JJtWfgstRjp+diw0IlbCHLn0F25y3gOHCpHDEKZdy1AtTMQc9omMCLhR7hrvqLN6
bhslu+m+gNdafMkylewsNHY3ggj3QLdNirLg080CnajB3HLnQt53AfbCGr8Sxsis
aIZ0v9KB/fOPEgvREQ3OP71sYCRtu5FCDKawX743a1GJlgpxcn4rBiZP89d5OfMQ
T1JjPY7BqFdGFwdEC87KniAzYCR7zZiSKE6W9dCEo/afmcI6zbFRhMFzF4uo3thU
AbDefo1rR15mRHB//mJCLw3VH3iXXbklzehM++NV7jrjHao4kJSxlHFe4rKpE4s6
L7M6SIZjwgICsQ3N09XPSCn7y1Cd0YkmxdsKA2ip5SMoUjz+Sh1O7eolJ4hTApR+
z6isXthDH69vhSyDwvcoRJxc7WGEdgGrsYJgzr52qVcXZyhELE6I9zGBQAMORiD6
/VRcbBUcenT22SuDMjVgs0XsZiiXKY0xUN7hkJO1xxt0Adzkk8trOzAmAVVeurid
uthuY4NOGdtL1WDdhKgIXD/C3i+lZJZcYCtHs/MwzKAs54phXG7vKVulE0tP8mPS
oGGhvKYNIpzzEhJeXubSKkIaa+d5iITrndNA2arr6Mp02/f6evcF2kMO1TCbDH5G
GjZ4TMTWOsGy1GIHA6vISXq/+aJpFWBclTE+Zcx4vkt6s8IVojnY2MB7r1Vzw7Wv
bLLL8mRLsqj+uZgfKmugJOB7ttGiWq2GbZ1DSI1mUPo+sJbSBdSE6xwhB3l7GcCP
9rc5DWWdGl2xP9p1ChEsDmj4d5d4kM+kEEPGzZEQaiG4iTfzdDZ3Ahhgmugsg//I
8uMbnZb+ls9LnnHymbNRLifzM1zVhJjsDUCrLMloEJ0WnmMRcw/IsbFeIG1VgZNx
nysA4M/X81+uMFQU0E/r1/3BP19ABrjezwTKXxpVNYGq1D/PFj/HJpzuFSAEAnWu
XnoQHpEucbl07QIz+IQwpCvgrtjXJvg+KuXvEGJ7dv3bG2X+qDl55hVBc3Ms5o9D
sumyGymKTw1+89a7Uuac5FQ8gCE/ZnppcjlhAywxM6/IhOY3dYhb3LGz2Lb4VfIR
qWruRJ76gLp0q2XIvgA6WXKbhnPq9B6pyVHwek2pZdlMuviA3WFKbM985bL6y/WW
HJNUtr0oBOrqEDDJNX2aEss/zfuCh2Y8YvwYMRNqpzs4II75FkkR7cOLHEoYyjvs
VwAC5KNubLOZguxwNqmKgrn/rADKV0zxv1KwTCv9E9GqQ4v34OxvA6C01uTvgmjH
gyDoisnC9/o5RpcypQEdktdUu4TJhA4YtWozg+YBSsSLqV3mRo+/H0fHI5ijdKvV
vTy5rJFeyS+FdLV4GSTCk6qb7SCDpgtAi9TQBrdCD37DrHc9FQ38fXQqza8H0/Jt
eLx9GQ52BZjJAeDy1FED36QP767eO1UR9fhR3NljU4GlphPDzQDRKAjy0uCOwZVW
gKLkq5e/X/3t7/zTeezR6qrIyLljQa99hssc/WMhe1fdWLrgMrr0ZYExk9cKvLjJ
kq5bIruUYPf4AtdeuCv/refi1Fyh4qimDT0UVjQ7InhmzrJXL5O+HXOF0ohn+hak
hF3kqf/sv0af/1PMHT2e22+3QOxxCt89QCq6nO3jJhrH+rYzsWboVDMUeNOEEE7m
DjpDRWLkrkj6NE17QPll8ntby8Vm5OS1ujPlJLoL2C49Ls6AQvAYjw2io4g1GX5X
eqMy3YYkl3QsAmhKiT1yCtsyTIvnQ/VL8mr9UK4pFN9h42LMKME37yIjS9qDfh5K
lXc2GXaq7QrgHbWoquDnTTa5/Q7OTd6yiQLHlyEwl0oqBipRd1AD/i/B7bfcb0M8
qbE2LEnpZ1NO5DG4H6lxIHVXMSZSbuP640ApXnhm8Vc6/56/4zlmiFu8YYfNJiA1
zJi14nGUgJeyAi7tlzghfx/p+on1cAiiL7Jp2nveCqovuzGgEa+REqh2/sNX3TNc
7qFGuMcQJP7hc43kHjuo6gsqNbhMMAYmOqcqwJ/9oNAsM3qvAeQXQdrxCxDphqRN
eiE/nkeUkkVAWTPKnKfxRsNoiGxoFiW4cWaHUhQO9xP30cw7RnNWSFCP94fjpa96
cNQIwoU+WkIKj7a6C/GYjZJQ8vVb00dO21GoFYPdreq9B8wgaYcXK5QePqWy9b0U
Bw6SV24aYBKSeXSxl6nUUlg7efKW5okIddmXR/oRm5DS5EY6im5ba6CGDb7fmAzD
cl+2SBDKV4W2306rmrgGk6XCe2JmceL2nq1JWkj6F4xg5UdlT5X5Mzf1Zhz5A7VK
3VBsACAjvAT8bEZI1gfFp0xzsQpTlAenq/f4oJ/mTYbmjJwrWRt85oHfSscCv8kq
qwwuYW73KzaOJMwR+Amt1Zq4xL1dzQyiICq9pb9+u+TuuB7sB80tRGJnpSSbHW9V
Xx0IeMrFIvrDYXdUZxGhf7b7kLG5/fEH9kI6DV6hCr/izagtllr5TGbwGzlgg6ly
RD6V7mnj7X8zuBw7K+14ucBRMisJBjZ35i6ku9HT8utilrH5uubh1foo6hfINCKT
xRRn5+VIFxj4xJbyv/S4D9st+sqwt8hRXEHTOgmvC1dWzNUT2KV0Ik7QHvzLKAR/
H/7fVB82bHNx6Du6E1Tto1FrkN/ryo32FZdhxPvdodcUrhfndQYp1N9JeD0z/fW2
eV5kKnVmMRRekEzAXeSx6kQRK63lGHI+d9gvS1EhwdyiDephmd2FyFCm8eA+xHIx
RGPOOnbHugx2CbNyrnDA8cYVGdv7fquCDHw03owiOXFAMULcg+PyOU1DN0LzkYip
lixaHn1aWUOjscI9zV4UrsHEfw20onkh7Sf5+xmHEx8LfAA8P5dduMJh7L0Sq4dt
dK8H+ImFutAoboiOBLnHmaqU/wF+vvrUqZiWr+7+JVT4B6OBdUNForHPW5CXbvdR
Gsm6oXHvRfSXdj1hyNNak5uA8njf6tmVo0z6HnkzXQErk75SeIts0+pC7kZxdV/3
O9l4FANAwAw+RptSwo38m1DiaXq6PKP2ukuIQGBqcaOZ4mCtxgOfFZd581ehmAvL
1G+cniWdRHDIOXmj5zcm0SsxB6M/7KOe4rVlcqXSg+SbBIqxooD2v0UjBa3wPVdV
R6nS10WEgD8UQap2HfTxYGapgqbE9xecR2nIBtW8ym3xiSnQ7mBPMrGWBvfsKjvI
/4A+0aZbZQ+xtb2z2GxaahiW2Cv1OJ9YRSYtTr19RkBYxyUHjbXcoZiRlCuwQdYS
OGqsWO113bhMSXnSeP1bS/7RI6T6cfo+D0vXX0xBVDZhDDknkXFiFW1yXVBrz2uC
/XcbUP331/+f5BQc/I1qUJtee8roTqsjjZQDZnJtDlZNIWJj0fgOyZku+KVIdhN8
f64lmUf0YMfmCWex99MO5q3I0BaMk8AOT1mPtSh64QvZJYr3ZzKpPSbHnZrBH542
siQh7QHe07ZCoZJbWkWzgljc9X2YKTcXl4lKaId7QXdRct8KTLUdgTf3KSXmm6DT
PZCoDuvPDZ/amQZ0C4OPohzmRm80d1C/U+4Q7lAk+aF5i6LNf1JweS8MXMHQgepa
vx4LKCmwUOVUr/L6u7dunSUMDRWUBtxIxE5Ene+1Zli+sv1jPyP0Ni3wtgcIy1/3
1n5TbxMbIBZ/TWslRLz6p9oIS6BsVl88WTMF+o0BQleUeHhheQw8aqM20S/8H12M
W438MhAeT5NhieL7kpxZLx1SYy0TrYYL0Zo+TTO+AV6TPP8A3u1QEKbmNAU9iXeI
yTjTV96/YpvIvfgbPHsinxmiSP3De49KOz3o65+FpGNkPNEORSKqZpdyB1BU4GwY
7iDvXS8M6EjT/55JVyGk7pe3MbuxRbf9w+hiGjFBN7veVOswGFwHDfDgAMC8f83w
300hH8f+EqHOe89piFADH/j0wsjUVf1hIxYBnacTV9fHUEy5P2t/W+Y/1L0vCC6R
S4MO42nghN3wYSn+8KiTxZRBOkHyOq/82eCipsVaThvE4OAFal+x85UNSpf7aJ4t
H4VsrimWXQkQUX1qZ205jF+qs0SdSybbNbHMPAlIxeC5FaFxNDg9JXXbKlsBjLVO
yRSazCiJ5s0u2zcP2zZFEUX0tPzAsQ2/061KB7wmVK0Yp86u13/HJ9vcQaRxXURU
XejSrJrnPMbGKcvwwhSRFNBQcqRyzUoSGeS9LGq2PgU92ZIHYbKq7OJTVNLU/MDM
1x3mC4lSmQNGfkiuTbjQR45Wv3LSyI1lKw1Ulkc/GXmQfDEDsJCfn6DGQFbM1a5d
tFTXMGZY4ZBqyE4ClMk4ofo7NiB1qKAo/lfrAxDFh/jfWWeCsm4aVKr0vE+QLmsT
AOrdzh0uG7s20BLXE1I/L2ZaE7T/l7vuLhoaa/IXnUEfQS8j9Ff4MhXcdE783L8y
qiamtGreWMyuGfEfMP6j0fxmOEcVioUFbcSyh81H6KH0MOEuWT5bwjdmgAKswy8L
36V6WOeM2t9qFSQU+XHduiSI6sPU2CmGgUaFe6YfHoTMeJMN2SDL+/6+MkKw7dji
6x3kigQU1YxrsM/N3LXhGnR2tW9NBkD5OfPp3OIAKS0WPRxnpcINA/qnGZsHW1aD
EOp96Bkdiqc8Wq3F2/UMsuYDFOOT4hUr0QfcGwJ8lCKy81UHI2OY/xkWa6Hibhqt
KOkolHlpteojD6+0pyEXeM0MeSJzjsk3gx5NsuWkla9y17eB/9ut4aIph7leqsHT
MRcUMcqhEXYNNvJek9BSPVkaU+B7Qs2x8EM9TtEe7GKNLFM8vZhCeh8RltL8SdxP
F3gUBDo3Qqa7hWre2r64IFegjWDj9EMWttbgz6V++oX5ntuSfvWlEvNH/0G9pLZo
ATyjnO1DBEc3lrvk5TM5ph/g2QdbLbwv4M/BMnHVbfryh6WUwiKJV1cjzxnTs8nu
QTVsbiNLzFAEQ4UBL6dbmKITO4o3U6TvKnIDp2uN2nSiWnyyF0cRKegPGQVurDFR
KCEcl6lDhq1Om1evKWv862owmxaL5L4hL+Sk1Xk6F80uFKZH+zTsebrvEEGs3iJM
aQeDPsSBta31MLifmb6J2ageX2mpbUnm7FlAKy9vgFUcNShg6BWwmk6TC95R4HST
AeQDCoFjiVQ+qFkqCinavC0an8wGkw4IAGROryApktq2JrR4xChibj00RNRXaCWU
AX9362deMCgWlQktYTtE8Ok3XxwpDMoirmVz5FzA7chw4pNTdDcZoelMs9bt/ejj
8IOPMyStuhcKT41LeJiGo/xZTMat/k2jKUsEz4M9EiHW0TzDHwTWFpfZAYY5dLZa
blsw0pjE7B2yCAhT6R0rHN2pMumfhX4y2rbqxPdKHa/osWM6+3VGs+bS4TNVmuU8
29FaoehmsBxZkOT8YwTG03e6/D5xtT33VxxgjsCfxZuDld+/bfl0k2M74p/L8zfX
vHkx+OhOahoAj8bqkSDC6F69aUJ4EMiTgjABFrTDoLB8hLm+Ff2TGReuiHWVh8t9
prIfcJaI1dzyiW3Wggkh1y6pM4YbuieGTzem+5LS0dpmUgHPWC0jm5buIn9LIFeC
ieZhLMCZAMTcZOejmxrC6XFjYpF0FA2vgK9rzmI9shDhNtwPFiU0EMVcWTzj/LDn
qpo219zqQ82CZaKNEWyr7XLkuMPVEawPiktOBqF7tsuUV/++FfXQmoi5RtLMo+VP
QgcO+gZ7RjyK2/69YPaelk6DGcKPJnTsmrtNucICoyoLIp0dfjULFAwchx8a47Bn
HjPcsF3Iv43LBoyBzOqvDtI7fOtwW/QDyJHk2Up045tLfYN9FBtYVBdnYTPWJ20o
0pyQT6WQxYiq5alMFuJ8RsVS4ViP1fiERZHEorRaF6vkFC0IoaLFvSZ9+AtkkhQT
iVXleLaW+ppcFTKijz7VdnSh2OkPjuvQw7akCbrvZxx7XjCXA8fhWA7SkTaTnj4L
T0KEYTxiJuZ8hk4Hej38FLCQouI+NqmVuCS3a6cxlaXWBmS8N27tYJNVcLK9dEWU
1Z0b6XUdSew/2XrweOR+BLM19q/o0n1RkvyBVMahVhHH/GtePA2Ltxb6HiH0Xrlx
SeZ6xX3RcYWkgoVBeiZclf8z/NO5lX3kCuZ6MK8LmlMNFOw+v7bJa5Y1WehqLOYZ
hmh8l3B94+yeaCNCkc0suEWqcxWrKoCXYBx5isTfV4Pq7ACmxsxfpN97fLqOXCPy
uyBRqUKELp7jQLyPrlQ1tQzosUsqpZcq5WuUiZAXx3F1+flLzkCotUuvIyKcfq3K
QCtCZlsl3EP7DDaCkSFVUrHkiCHuDlftwWxfSvh2MaVEv/q+WNAY3iwH6vCqSTWG
zOjEVOEzP0kRsoMIyGa97wCrBhh9npI5u1O5GWhFWn0lAs4wu6KU9UlITYukOACQ
vjxL6wGE7jO4GFtZesypm+rdEMNWEByhSjpkTTM3+HscCFl3cySQLBK6s6UxLj1c
gHQL7BMcIsBoq5k6AItpRkvjvIsXXv6qYf0iiDVM+nlk7T059u4Q4CbLFoOF/Mdq
AkY1RhXeJJyHN+AUd1gwHztnG65Vimm7rwSkuGCykxsHgkNrVChCJ684zrmDteTB
SBfFLY4oKN9DhEFPX5zgodPiCr5KpMydiPWW8y9wN7IFCXz+nsquVQ8Bl5JY5abS
/sMu6qM4ppcxSJi9IOC3j5ImUZKhYw8z9rSd7L2Rf7qohqx8SoDF4zMWyDBZgqyJ
yxx6LZ9dePeeWTqjc+ycuEzKNeuuPjhDvYJ3jMOl2r65hrSC4hHJqPXSNMrKU/OD
uxPj003cqSD0+HiInW/PuNwrpk8xDUP/knGvULUDVEQKrHzFF6H8qXSBPIE8D6aa
ITP8BJtRY1vCTMHSCpMtTCZVk/grVYBJCgejGZl++fMj6rjfrKmTSjCAa5tgb9of
8cdCwIc+KIgapXCsWErzt4N1Tpir36lfQCKi0x4HdgOignO71XvyGCmijQcswVkf
5Q3jAgN88coQpz7X4hbQvm/ZcTXXBI/8fJYpSMcbwBTXOWoF2xwHNFV4eXEhKNAq
4qPhsq2zsOp+GMQfIlXGa3QPE4vWgZIjvo0d1/hjkNhA38GBKNYOeRITw1ZJWBdC
RlLwKUbH2R/vFBP3NBx4wtLTSd0LM6Od4Gr/wn4du/rDMageqPBjcJwtakJxTFxv
3yKvKOmM6SOhZuAYvhgmyF5ms4e8dUhmHw3T9p3kim0hLgmLG81VoyIz+0Y5e8lm
eEHNXWs+JouAvvu3PNF2iahZCd8kdlxyU7s2cvCUAuAh0qbjMncY+v2EqE3VBgJp
D1cEiCHqQwA7ooIn1gfzHl9HIDt+tFf6bDoNRHAtXFaohH/XWDpmsW5pBZs7A46e
hOhXVcqtnIqQVgkjJhPv+xQ8B5cjy7/kIWO7/X/WrVQ57kAQZPe6O7vPELcJY5jO
ulEXIcPDG3HKLQOKxsjJuyAVdaQRMxoAJwcUNQmLzd4HbZTUaDsjvMJ9Id/4P7jO
Ltc+S92Dbzu8zsuc6BMBRT1sVvKfyMeeV+3ncJClseJ2jbPQcrlZ6ZT77E9+tBup
yy3J7U9q4ql/fkO3T1//8aLGwILspydt7+zERd9hJwpC9fjJIDvIaVtPrP+J1BnB
RetsKZYtc5jwd+chs+MtTb+YqRKgxBSvLEDJanaOB33rcYGwj11ManU2c4/9csP5
crOGnX3RmjRQSfxADj5e6fUxRTXn1jmhtK9oi4IJzfX10Yz0ssSgUe/dOEM6WORq
a2j1wnPyLam4X09FpJZeGTbZ+JzUudh5LE1PZ67uSUhvwmz4RGCHOMmD5tbAYKHv
6fTd/pdRfcEktKS3WOTSpAS0jAxUTHzw7uwTP4dcf+q6frimdsXad3LaN3GCqRMo
AhUc4QQvNteDxpOqbI2ZKGiVf36LEMivL17J6VBnEPAOZozdbuMV5xED3n8CPWZO
9+rdvDO7m3BIKAv2XHPRWFv7phmcFXiONPA1CN2+G+XqjVpzFFViRUf4xeClLZhK
D3SZmoGocKsHhOwdSMwZ/JEBzJjE38vGtjW6p7SI0pBR2o10Em7fdVQAZOzbRX4e
uur4HE1OJjiPL+7Y0IdZ8L4JIaQHhowdYxY9hD2R7If232ooiVYc0OPgYMCqiqBK
LDCe/1s+soNTRuMZAKIq1JvYRbG7fukTUSBsx/x3kE4I6kneWRGWs7tzR9yy0k+b
02kF3gomCc2r8AiSzXztcjaEZETJyViidLf/miWmffLtdy4JnLwLZMpYrP6YOI3C
byQwxK6IuSyUmJ3eMnn6Ow0T8/G99oE2igJMbCKG7WsF8EDF9oK3r16DBMq3uose
H3g3/FqeX/jvbSzsm4u0jwYDVGj0onbf2rCCN8A8sENsErM8XdhRCEe59TOmxAIR
A+Pql2cKBgWZwTMTb4JdStmPllvNTH3Z8484BsQ7I2AmSrM7uqA7hUNhqVm9MAYc
RssuEeAgI6KPhdINPJ12Ux4FTv39J4QTSBXuzLTHK9YKPHyoVD1Gfb1ToonYoo2C
Cemr2ZweeU5x8eh0DJ0sYhnG1oxFc5RIn65WigomuCXOcNsHtbgEH0ckjC00sZg0
vDjNlTjx79r+QtP8/+CGR1YUYWKi0Eo0vzPC9zga8ezqQ6Tx5nVxuSCXPAVHSa1s
jJulzrINgFJ9t7rdfYfTColLEtISqhHwRwmZKOgCkz7LHf3XwsAenevoWGK40DFj
xJbCXCEFNu/F7RHIGrwPC97a32cLAptr8I5IJwTZat/GiuSHd/n8fF40HQkw9L3b
G0DcgUY4PehDDafUr5R9qpAl96+aVU2U4IQ+y8FKdAjhoY2pufQIbNnhz1ioUL2R
JBAyFgTCZrpPo4fiFLrT5PWi+cwOGpV8m3BLrz+giHGwNgl8fls4/tB9r9ULOZMy
U+2ZCuAqoc17CzGtl5r5AuLuCpLQNA0p/GxOmk/RY+3ahjRw5B/9PL1aTU5hclC+
0cgprF9vtUWMoyM0AqQY8RQkoWOPScT9wSblcrR/Xjgv4uCVTWS3P2EqGFfbFBDc
hJ3VwC4yv9dhslBVgL945mNavP56iZ4RhCi4z0n3X3bk9eyfJgh3hWkPdaaKMsiD
eJUvQaD4+qsK9tSFxdPuRpRJbr3sHSp/4OC3eLgqrzHh6usgRgWZv4fvdZXojW3Y
KrOk4Y8Xfcn28Xb2IhWtYi+Ek24QmORTELcAbIaW85XZiv6WZ1POEvwqlnEZHRks
U+LmBdu0JMFIE3u2GQoOY65caOdASmuRHtg8OFYYlxEfB2a0+42YkmCUb5P9nCcA
wuSLSjYaGIl1WwvEM79F3svcx6A1997rEzK8/OMVQi84xbVKovN0jQRrLT8qnTH4
f9iIpPKdL2mTtXbz6zagNKDq2x+JhQjf70YMLCNchyt22RxvS8/r76VOzj3eMusA
3B31GX8HHjwVEJVMCAv+DVxII7irX7slApcGNPvvrUIgvC4FiknYqA55GasPGrbg
vS5dO3VlR/8Y/8w9fk9vdAL6USeDFrjxRMgu6d5Mne6lzU95BEgppNUOUbpjBBe9
SuFw44CWz3JmFsXHLm7LXVsow084lg1GJJIpkpNdlQfIlIYMztysTEi1jA2YGBUU
yyVdmPaQfIIja5Efwvgp3jHiE41R6oqH8YBOz6UdOdN6wXl9LfVkMW3AvSzrTVy9
Ju1pfUXDEp7B+e9KDpqTo5vNRe648/+wtnM4zOrmDX6lw7Zs0MCFY6wLRiZvi4Pp
W84sZuU5dAowCf1dib6ArQX2i4fpPLDM/ZSA00bIieP50tm79yGqHw5mA5aUoZbn
yEaeQwCYPaE31694M2JE0/LDK+TsD4eoxRWt5Qz3yN8aWyxMES2epd1ID3GP4ZSy
zW+C/b6CLwJLxP0h9cOvnK7LAFOsU5rG4Fzki/tlbbYjvUorViB9KuUcajQ26oO0
FzQSTU7MhIIxW0RgjLRvKrkzElt2rIS/6jFZNwf5FS9X4iM/MFM7iPex3I8087XL
Ae9wzrbMOovBEGZxgVqnElBGdBqfS7Lxf3JQieDy5zdBImHWpGOxqGqfNnqcIBKp
M10tSxaOKVD8pLvxvJ2pxSOYy+e8Qd2fv1QEqcu8UCO5+kt5t6WsOpByCHoN27W+
mPowD7JSd/Js2OIwZnsOg8TzWkXvu/SEBJALw7hseN32kxaDKlJw+wvxhYvijqW9
t8Grln7SBD2QuPVYsAj/kAGe17ksRGjBix4B8ijqeUtReP1HW0/yP3d1Ga+jW9/H
VmU9auZWF/dd9uuT3uJw0Li45o40b6NN2T3Ls7dprQgwG8mZW/3sfV5RB+EHSm6k
+xzN1BK9ADRR2Z/MTlYk7iqnVC/OiJv0J0PoeBcfS1yyrDMfckMEuqxC6B18mpnR
UevLEIjI2kbvSXcSdJjAfS/AeCfYipi6uNrFT3GuAWTn2RGcj014AlheOKfFNWSw
SZGk8GpSbBfdVrSXW0cmULgkkPIk+pgNQHgNxSKKDqMm5uHbLqsr04JIjXBJoq/a
h2UazvjmaCSIJlCSEr+QL9nGiwmMyUW/revwxmSshObaMRd1nPqNEE/1qH22j73H
MVE/5BHLLEzyQOYYflt668hLfny8tkfU5CRsOS2vOCEi0FwvCW/9Tbo4J2F7Hm6g
AphDS7TRTMwtPokSimddiR8JhjbBiXkXkQ011kc6CTkhdHxatOvEl2jXvJRZtfg6
K208pPKtwxJtJHhSCtpcsrGmPjoJlbUi/pLIANBXGudZKIpi+XjJzzRzowFUF1f5
nIhxDmJGDpwPZj9inHQg9h1r3urW+APoJz1/maUtplTAEERJ/861NmEN7hNRttz8
d+zDsHVIOYJ2eEfgtgZqXBvYpKTgCgrg9tCCjUb4Fd+10No9FfkFqb88I+1PaFEU
lpGR7/FO+8gxoYADGRBui35kUGCVw+KCkmxjdKNNLQzmZEeKmC/ZtATFl5fWMomg
gbuaqk9fyPFaD9ZOIm3cM9j8wdlRhyU+v3yA+MV39oorfA5ywXeOSuvxz3ZHZrqB
ICMNr5pQrsnA1HFg8DRqli9TD/SfPaekzXDl8lieQanEvzyIaJEN1Oq5Obmtl4D2
OPhk1svuV16LSnrzPSoCyM52ImkWcfK06sHuE/Nh8tRm+LYn45BhHIaSvzVcgi6L
6gEA+ixYWJeotP577KnEsl8ZZkgLTWCRJ0GT2/BFwLLYY5rfeWkhv/+rqFSdRL0c
yyIU3RfPYrs+mhNOrkmoS1w4MRLh8xzHN42CJ1RREViYTa/RK8ilXgbvyfyhhycr
TSzgctMJu80BZsb74wlHmHjEDo0qZEyDrls8mq3WUfxNNy9PuVdWTwsZeT0FXwGp
EmZarzSr2NuslpVKeLBPjRWHwzTaqmKs9bjTJvZ30CgtXngKOXHtqFcjvCX3sfqE
Ob7NKuCl1qEgSczfIzFzgszHlkXkZHf1JL8kl6xf7HaWG8CPLVTmLtyHhO55i+H0
uYmOMfAGJPmeQjBMet9OAHkbaAqUcahQHq+nGrzYHOIUYIXYib7+7GKqCg3yJjLt
SBfvw5St2H0BI+1ptQu1yQ53kn21ZdV8NKnfP5ubQIv817LRnGhf6Ryrj3uqjjwm
oIVq4owenOJSB/euSTxR3+Cgme53EpyWblotDz0MqsYbvoxSE7ytj1egsVldL5ru
XqfJqkmxeV1kkBAZB3XFJcA+IAlCO/5KnCBY8al8dJpN7t3veUhB/n3ZmqawSzzj
CahhB2sI/uHZW+1BrnH6v8RaK1JQzS7oI5HeR26f7rzt0XJytLWxpRtAO3hK+Zqe
FaTSZ/8ZH2qNIt0abk2i6kbW8gz45REAxRYoUk6BNJAIAzXj+DAY7FqnjiQKm+nP
rKSgygx4n2AovARXUDWutbaAFyDiBe7F450UZ5B1TF520iFc617mqMgvd4zcdjZ3
bI/WbwdNVQU+DMGviZh+IZaAciDIlckHsLT5+5kcQgNmUhp/WEGLa4JC2618nHJr
Omiotzu2Qg/S+fYMqUKNKCfyivRxFxfENLxRdm8sO3y056BO0wp/i8bvN0aImVqq
XHn3IDAs0ZIGlha01fvNYVRkQPQ/mocWlkrf/DSULsKO4NFBXmz2v7grPprJrml+
Cz3LPjb+EazPnkQ1XZt+uciENRISf2959l1XYtLYg+57xb574t4zDAA4KzeRPABX
0+7na1zaLlIfR0wF1bRr1RKfb1Am/xyVft5s1HmIfmkrzns4VZP8pH4YIZg1IAUY
b1HtwjrRLqowUNj4e02GEj2Y+P5CZD2fK4Yjp/9Rkou2YizpIDQ6pTDs5IHlyUCF
OafXidc7mBqC3yRDagaHvT4VbyGcchw77GwyKFf7E+3/7gm4se2O5qEnquSvSHPE
tvj5A2AeR+c+IQFqc426kjPkx8ibxGQ8XTIQMaoT3uj/cbw1+TvvzhZzkSqrbWDJ
tKoqBjgUSEcmkssIDIUGxWKsUUnwI4sTmYiuzaG5jWeDDTme3ebe3Lt9KYekmGBx
vXijZJB432JU1oGBR6zilAjOfxtDFmEmrI2bBa2JQ1SlZlQaGX6GH31E7dfcsSIB
QTsTnkqln2IM4CrZ6lHjI4nO5RJIHCJMIZ1E7BaeERcp56R3dcynM4Q1UN5OpolN
5CBcmWY/o5hrW7aa5Jsel4TfLUZYTeGv/ndnhlwqJwIErtPyPlsHDvfQ1zHDcEBe
jqf7owLg5nFMZ6dBc1HkAN28LtXj9Jl4a55hqDwQjy4U6FOK4W+wS8XEnvcCbxVX
5FpMOJKb9yolRvAvEbDV6YHOITu565Wf1ux+cZg57+BnPV+BL4MM6iyjgOfeJvvd
ugQX9YQeqnjPEuMT5+GQ1S8tKIk+UftDv+eQxdSHd5YwYgXEoHt0x2cKwD6Ymo+3
9E3MJfugQs+1CGeW92bDABsGNeYuMqSt2bBWrD//K3FhMVaBwQefwFhwytoxmbDv
YSiChBUj5kNqN+VP0MIk/O3CCQLCvqxcrBEpkcUWHYQny20Kuituvbe42YO72XCS
j3oDdZSWojqQGA/8legP6672MuP0SzJ/ZxoOnQO70mDegXyLahDoEsTtpnTeyen1
eg7J5VPp/5s97Ct5/kQB9ITjobx8qcMcyKSDvpUYkU1LhDGS+X+/gL5uElrNQe4F
DCbQKM1QuMYyZKF/AWY7vjlJxuRq5GLqypICVeoAllFbWLd/+pbFhsUi5ZgrmiJ+
q4t2sTiCw5/0LieKJqyTWblFZmrLlUG6zh/2B6eSpKMnzAhHjpE2yjbsijJQaqGM
5dPwTu5BoAbldjdaRagbcrUjPsDtcQWhXVPIy/SeDqNwQHTrna+GBifzwnEdXnlZ
Guf0c3xcEl6iDg/nbihk7jY8TJnYKqW6vDgX6W0RwIpMxuzOhrVaU0JCIrIVGf0I
iuBB5i2WbU7hp/Ti+4cYcAPEW34ia2wvzs6vLUs2WCTBVOkwUVbDhEVe9zlpYgEc
filW90Eq/FJmonnAjUjkNkRMibK78OwGgcP8mM+nboDaq5RSkIOKYn6ytFL/6NBg
2R7/Mm54nnqlMAX/YVWUjEW/PnSzd9DZZcOkkMLv0iWc0ZG1Xugc8Hq7t1QWZAcs
Ao+/z/B1+qWPm8TLxzR27+aeNIH9wu0w8yYduAQP2zW4N85IRi7ar00TLs+HGtgR
Yd8sz2A4gc3tj5lwdeX0TiU9EmbzID9WDByF/8B6hxgsga3cwxNR62HIptgnvQw1
gIweuil3mdTQMT6CRhpE3HJD0z1V/Ar/myCbaqm/QAhC2Hcly0mdnS+b+bQ3w1OY
wnmhYV0/YM8auSZw8ESFylGO3eF/80cKXCFRqAG1f6hWw89rRgYHrF8YzhPn6Sv+
Hf0i7wNEv1YKv82r7nf+x6AayCB/xn/5oqQSL+zDfMgjpcWiDaRlbOkPLSvxOeNb
qFfwoWSETjgbdDAP6v2Gxf63CdcVlImUE29MYo+MxDGvEhQv4VnHpHqLGHwSDPXZ
9Ob9eBh8ndtrg+ZyQ6Z3z0wUUxYCtyT0PSm2hUcgMMDwVMCb+VttuvLFsrbgIVhM
oiawNwEs+kfMtWDDc6SKE0sIwLa/0hePce2TaZnnY4A+h2fXlh508Ur6/9IshA1Y
IFF9xbSYVmycXJ7Uhq3QXGlImC8e7tbWzhNLshUoLLzT+KKeiVmeJetyuBWDlI7B
V0K+adX6Oj5V1P1NU8pQBTMDJxWVvcSbia57gk0jqAKfRHFvlO5juFZKD8ryDTcU
9POPCaXz7uT22ZGF71Xlp0f7W8FwNVCGbAKHtKkJeE1VOMPNjz7DZv0XKs1KsNSk
om5G4FzOjhy+GVL3HNM6UtcKxO0VcBdyHP1du+SQPiyQ7x5adq1IheVokqFDADRj
J/tcPz/poJmI1rWaobaNWzX291rlJD3ZhPlN2NLW8Cb7rUgU6vf1Gp6LG++sH+EW
UBiKtn7Tk1/LR5pr++fmjjX2QbOzaMWCY3JLSPNCKs3DphsGbfYNOyQ8RTLVMy8g
1tuZ9Z9xLdXqyNxbNNph+Zusd3GfNZGyq/NQGD+n82wEQxnmYP7ZWAO07RT2CCEX
fAyqYzPs7ySPftM6DGlkldpQU3ChgjCXbqtr00IipjY9y3/wB7X4+ZW4SY1NJ13H
CgKkzrYraMMc80z1BfCID71FwQdqoSOz3Rvr+uNnctVllROtf2Mg7VPgRpliXKmI
N6wlWbDqK6tGfwe+Q/CHc/CEc6EN+4LzJopshEIEVhpI49+x3ElJ4zhBS8RN0ccU
R8q/TdP7Agkpadg/6apIBQjQlo2wRiGLAYytdNdHmymJ1k241PS/CL2/PBapQes5
5w8H5J7I6316nOlEMT055qNsxT0Z51XfdlFGptwSGNM8yFNSs38n5zFkJrL5kqJY
/sG+GgnGB1fOkJwklh1U5EHT/TkPaw8+x4JDPVt35ihtGZPYTiXNc4UznnQBgmND
CcH2N/tTFEb3J+YPscdTBUhflOSH5XxZB84e6RsRxeOl7Pt6GSVOdqGRkD1h5J48
n+q4oJLPhAJL8raV6pBIttJ316slBK+2hCYrLCCtFnklhVPqF2v0ahqFs80g5Z8g
TmpGxBe/XpRyYbZGEbdrU462LUFdIAGVgZahnAGghil9HHoQABE6qOs3qiwy8qaC
emWFp68NGYSqUkoFNg+FR4zKULEd0O+6IYeZCeVVvexNZZEDa64lS8G0Zb0DuwmW
ukqEtxkWmoRxP4ZUXLXeRjMu0v19WlVupVYZRsnypmYxP8ia/UlpKkEaNO6SxwHW
SXZmDd7vE5ovVUV2SGeDIcoinDPHR1rTUcjppJSYQH77s4xk+hHAC0t8rzitGmCO
Cwew8HHHIut16H5c7WOW7B8+wMkP+7chuEAurz+A2PkQMtV9K6mPnHUQ4djY3xY8
XpGq14Jmm8eFMN7hoEBieq23/rp7dtncwVHklGlSYJ5HTiOqck8NIdYWOi90fTOn
d3AGrAMg27WxYx52dg4OXO+zBq1zIfgtejFyWkfvD5NhMcP0sSG0HVn3WpVV0hf6
6QKTFEjSYKyWbz8ymC4UHs4CrHZmgrMG//9gHh5wgOXzZiMtAm5SE6AfBTzRz4S4
+Xe+UApKBIlkhAqJ+4BS5fxLObV1Iu1ZPf+BKDTb8Tbw4jhinDvPxfXp9/GvHuzl
cWOAMArZs+AtgDjvw9ZhZiSU4tD3Q7WOPWj9GWGTX2q4fATS7o9D6fKkwefXe5S9
a+YdhOtGzO4aeLzJSK3D1wcavFQFpPjxmhHyumuBc7Bc44hO6OBYJtWae78CL1/C
ajzbi0RL4RdOVVYwWFuh5TY2HxK2l5rYmsFAbDUPewCLcBRP+8TL0qeDHEunYafu
S72hCtFMPwMdubY4pwuphmECXl4gnYkjEO6qBPwe+SD5p8hEQKi9vCEDBunwwxs3
3Jn8H+J62A9pAr6iyr4EgSKNNDBtntLVruj+rW/kOoiSpQPxYiGLKlEFxbliJYxY
QMk+kdgIgcT/LmgoujhGNlyzHRbo8RMHzgoxwofNQ4NhXjZQkccbxiCeDlQog6Qh
ZbvLLTT57q8OjUqR5BGePl4GVTMiZwI1YlxkMwLSLfku4bAXBgjEi54I8rJdjxer
ZYJWw17Ak/T9cNy2UdtuvYZvsCp0fHKsGUpFaLqAV21Eua0TE+AX4oeLtGylzHG3
xDTYdLDdXRy3Oxtz1L6K0y2ph24eAZhhBtuHhmECoYm2ZqDydKc9Ijk6xovg1Snv
w01SiM4IMOcC6hs4F0UKetu+LO61vfU7+wVTdbiQWtK0ca0fsjf07wgIdsMfCwbR
+NzgPseunkRCN3iwa/RT7H+Gp520jYDpAtxUMJlAxTcDAUm5i9Up1v5kMfcx+p2d
FP249dXf1w4rno6H+98DUuFzozXIXfCQGeuK80gubpaxWaG4Myce8/HxO14IH+yk
FRC2Ic0KAU63Cp0mYgAlFW+RzFwz37OD3nptGHYEOcJXuhJfcLdCF5LQ580AjOBB
awAjbbvACZf6/oqyiA+u1a0wcA6XWkbCdHqvaAHdrM2+8rP0gJG+sZvwCzjeyuMg
0Wvy58CXvjl9tyZ97u2QKxkKCXp4k6eA3h0K8oHCNC3qAcN/Lr6rhqS4PFHfOmb6
1tGJOvNYspUdYIZwUmAvim/RdZUdy8+eyOWl9GeDezqOhBrpEvZ425r3nudDUTOP
xHphdToSXVPGtxZqhdc5n8Ae2HWuupJdb7ejfdCcy+gpJCFLuQZ8j0Voqn21e5g2
zyIZXULWsz764r21U7yaJQ==
`protect end_protected