`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 2496 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/9huKRhRMtvnNqb3Z+UU7TahEoHV+T8U3P3ufru7l1O
3DlgtZzb9QxCbOjthp9+wDkjygH0eUfDrEl1ovhZG63IrPVD9PvydVccdM+Ptq7M
c8obqSvZ1L0go3f4z2t1ihWAMvx+4+5HE9YGR+VaLvl6R31JH28cwmKb0AOJII0b
ON1VuKnQAZy2+aT0X6A1dDod+N4xJ/dWTbmPn6OI/FDnDF9DAKJo9yZ/wQzQWvCj
dvWbN+2tKbppsQ9EzOp0MrlorOxmSbP0wauWWoAh30XPCEXmsoNQIUIZZAMTuD8c
9jWbCMp/U7JuaO1gIvmo1nTvIPBPEZrVKEe3EAx6uiyKqhfCr7+LBlgCtb4gytyb
G3FEzbm6tDZ+hNPZK4W5/8bTJ2/ZT97KQrx9Kn6J3cHwwKQkG6F7iXccbU6Z1yhP
LCLI5waX+GLK9RISmxgpi4XQa1EA4WmoGeB5q6QnVBS5nVmlEMGXSt/FiXwSBxj2
kKan+R9X0xhZZLDPzyxQwZhH7INkF5Hoh1gisnh6+XdpyDnvljZXc1jsDDRX1VYH
Us72+p9qz+xvjNB0KSig6Pm2m52wXNKbpdV1J7V7s67YXrn0VJQ8DCwUi9b6eWKz
MlIh5hNblajpoBL8ASrW5U76hZpHS1Xc6PAbj2rZIZw3rVV+3D11kMqlMfJNLiTU
Qdbg518w8zLcjlx4XK9d7z5jZH08Bt+7elVsNrpzSPxkLzbG+q9HfjpFphyDqGUM
W1J7bfMxR1Wk59xfWmAzs/BqXRBVWG3pr8AhveqC38j/fVP/oV7mJJd6ZMILP9B8
q0kExeFSwnJxlC/LSBFV0l8+JZmfhRAjmS4oCmtQjd0AdahDZhLcL22husjAFOAH
nYCkbOMnpZ7skD6IM6aq8pmiP4IuEDvtY6IaDxgP/h5Z59LupCju0+ou5dLaogzL
/KBtkRj6nBFKJSRH5k5+jkQ7K2THo1zbu3xU1l4cgzbr2xUeauD2Isbz936onMBl
/ENWoFCHGIW2pf3oIx4ktHU6orrVPrqT+ZD5w/RvS9p0rA3SftL1oMtxp3aK5VmG
JQVzGQ+7JvXgZneRHp8Ivo19Ll+WdFumedbxXqWwA1Jdn2vioxELnFNVnCXagtIN
vrh2Z6qdvtMPwvKY+SeM3LrxhU83pJUxkt+wyxk/lI2zijraAETDQHecMXLvy++h
a8Q0CErLB0pZQif3kkBDi7QpkdyRcUfQ8Ccd4/BcZ3W6ArPMKNBvhzMysk4ECLzl
NtNolNbJU8XGOcSSrR888hqa47G6nEK1q5XkPSM0EgeMBxlnY2iIJdYOpJJDPmXf
zcSKfQGHPWv/QinCRVDN9nSGoYR35HeTd4qxNooVTdUWVbn6heGErEUZgI8sEAf6
kJHGdLMnnF1adbgHZFtei41CmhvkGItG1xdfIRBAGRyR+Ivz/Q6hkqTseIhJ94gc
p9m/FwONelotVC9OmsB8w54h4z9q+jsihCZe0LM25LWiJNzq+MxDH8Dysc9OxSKy
RfFCf0l4oJayESxf6SFNfpnWXkcn5CuA/5lHYKxzHcQTD7wYSJpyB88PH2bhaHX6
WxxBxQGCs91Si6D/ByqfAXQyo/ZfYg4JrfJeySVYZcOFr46Zkgl0xvCskOt8ucou
DkBglzoelgPL96VJSM9NGk4Ge033GRDRz4dk2nLQYuNzvuzSaQfUpdyX/ZJEbCLc
JBcL2CvqhzOy6i2fQBAEQ+JD0bt4eHO1CSWsyF3Ph2T2wfsdX71v1ThbWg3gJS8v
jVCwVJlkMb5GS25eqd5cegiW8I221tZL9r3B1zMfHvykJqcHZbZd/0d1p+RvVsmz
rUEg4dkxASI0V3EDmyGYDjbf2n0tzFvmLQmmuAOkWyvUflw86mWpefB0CjsdtrWz
STB/2uDbhf+/J/FmfCVOyPu8yRgxPenr94ZdG1TJph1IoSjIIb2+1WXl1Oerf6xA
0J1MWLBLdwirFhqqB1XNTB+UjuXtNchIJdP94s/2Ww9Dcp8YGpVfZy6ewKGUn9/I
ogpZPyKXoUH2/+Drcne/naPi07lS9iJvRL1afaBODLAIIJ2zO/3XsLUtxqJPVltR
/4BPcxUwjtimc74vHcnnhunKbEm4VVqQAVfGSawhpV8DJk047Y/6OGEyjD0BPvY2
NvEObNKYpgcw0r6GOvllyi6DOIi1biVdocZeYgWRzYEubVus08IyyqF+qlbNedhm
1ZOZk5fxYA/oYt2NPHFiaR0u2MlhNEZ3B4J1HdXA9Z5TEpc3vpQyG1suF/0HDVEs
2BmUt0/9fofUBZhLiReMStxEAwB57l2VZwf0Gn3zlidKdib/t4K9RYN7k1hyzThX
hrokYlbVXlDm6ybZetRcI7x3aP/lmzXMeUYaWynNsIG33yAHpPLvTf96bikkjvA5
tybGQ+bNy0tNndZqho8NEXSiH4TAfu3BObsRT+YYj6jfJgtSmxm780/Zu12+AL4q
s0v0RyELCqhh5E6ZqHYyqM8uyUIVp04oxVb4AP4D7964pzsm8AEjARcp0Xvt4VdW
H1LpFLpnVnpUYVr/fizvOM0RI2yJAkmYr/bHS1c4q+Qg0AcIrDT8Qh9MLTSzqvFl
J3BqmtIRbPdeSGbZgfH7l7YC3GeWNeSCYV/0rpOoSRK0o+DS6Fa1mk/xBAFsK92Z
Uo6ZxIYM1B/t2k54uXc7UuYarl4q0Sov5HUXy5214CsUl+bJptwUZCX5MzwRFHtU
SPJFNQIO5DW3fpsZCbZ4tH9mneiaRlqPR/cjW73hzOp1zWaFMex06LthaWmvFISB
sKjXomYlDyJvjEZh/q1niiHJAV4/0sykYJQydxGRA4ogWBKi2V726gba/2MXHD4j
2rkcI+INsSZFuSr53DdTyYsKSzUomP6A9rvDShXrgWogFpBqFkgEHfxhiuPGRmIQ
T2mrUXOdZkrjPJ31uk+pRUBFc72A7rThSeCWzz+GfIHybMliRBicIDWsgG+Z7A1q
5MEipHKG/bizvi0Y4P5o25gZSOpMtYCKKeYc411jmx4GW0yJOqUHFGiYxy/ai1zI
WCpqlpr4il7fElzrsMe/Hl51KWmmI/YCWGloCazm8f0LLM1h/jDE6CYmnqvI7JeX
k1gGaSTh6ralFrEzKQnBFb5q4+eueucA/Gvtx7ov9iCXqoFR6zfBppCI8YzesFNi
9tel1SyDTGywJuyVJdpFQYx1eQf96aec3wRdzWGY7N1weQvTTqJEmP9nhJ4qdSjB
8uxcXLtKzELU3kqhyrYC1paAPFdR6qCE40BhNjzhGzipLIBke1W95qKgKSlxF+rG
`protect end_protected