`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 2912 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/9huKRhRMtvnNqb3Z+UU7TahEoHV+T8U3P3ufru7l1O
3DlgtZzb9QxCbOjthp9+wDkjygH0eUfDrEl1ovhZG61jbSdF+mr+/cHo/rem9aGz
obPE73nJajb+N5FRI0Yb21ZgLybmAcog7QCMgp/jxp9tJMYFZejazV8rBH5pCl+K
Gqdfirtp9+dVxiBFqLdOf/5ZefU1Zyj5UdkEbJsnbCxzLP9kXrG6UO4zp4E80ptQ
97OaKuC3+qVLPn0kbBko4rCs/kX9Cv8yvSJx7gFbcmX+sMpCFzxhjRKNoeYTBi8F
kYTNjYDtRNR/qCXUp7ZwVLXDOi27mPcke3AEEkfxQSuMpDaEWv7R7L3y9g1dvNGu
IyX/64kgpVsL6ks/lTCNIFhqpvAaoKYh9bnct7Eqlr+p8bwYiYw3rkj52IG26JQ5
ZNHNFdikIrcpf+D3xNRvAnspgwMG4r1OgC8xwNA4VQXOqAmPEC8lKVAX2DCj21Xe
iLlNDhijGcU0zJzytZso8hZ7zSvCOpZGETCvpNsxEKRmJlCPvwvr0fxyY8KInj4/
1aC7ziN+j9eHt92UsUBWtTX1Mazl1FeqsNqdiBbpsA/w/xyl0ReT+rSpP9wvsXbL
IruDDpMU66o3Kb08Lq37tQ0ExHfcnZ0IvuCSynia/bpmKO+Bjs0k6ZOc1OLT5AIA
mob2Qn+H+aJlIHcxakVdmISaaNcVxyi0pp2AwIEooy4fFdOtxC2mUy7Y7YRbOM35
8IOLF3UhbD+0cF2N+1jzyBr7UHSTOyhgykGzXbLuOKrs14LfeAwXFymETwrilezh
8WbLzONz4anXpPoogMm8m1HUtcTsRLXuJFgu9K3oHME/vCFhDdLHVUe60Njm35dd
BYaLBYtSAQ0zGh6txgUxtx1OZTol4E793AEhJ9l8AfIA+XzMIt7eoiba4sOq3378
gvXQ5sBrzvWD6IJI/nm+Uie1ksfusyxHFOFyQg83WgqPg7c3xKXLxLBLDPI8zZIK
AX+TPcR+xknOlli66qUGYN8Cd4S95drZ0+vyoLBjts2Mayhdw9Q3so1igJG+Dqbm
Dvs4X6lSPsJ73XE9lhFO25IixO6iPRMEzRsBo9jpwDxz8OiUAmcilRTSx+vno6Qt
JbG3v0CfvAITS8U0oqi+wf6tjGEhb+4WZ5hSysjeH+2EWZ3LeLY/Aix4zWM9dIkp
s49yHhKujlQ4j4Sz8ydFKn16iEaMe4oopFa6jYJhsg5SxLNPRc/ukCnpkFneemhz
ZBSLoRYPybDGgL8prqNgpxD0HiQT4zt3kl8GGWzlEMFI4rjZfow0oMRjNe+YTM4z
3D7igIL4hl0tT9eCAv12iR99dKvV7SYEGsDKibEmA3SqgSWd5pnMK5KyNnK8VKS8
28AWMcfWuh0gdi5Y1x8N+lKQQXuoyYepz0DCOu4k4+ndRp/hWrFHfvxA00yHhWLI
j/ikNv1A/tKYQYYHp8Ien5X7eRYWMlNJIpm4yd36bVHGF3+F2ncwbcnJSnUnTrYw
fOqdAXTl61pow4KLFqYW1QycxHA0qD/u7CETOcllNYHQXgivihnVfGNisbnXHmf8
Ma3yPQyXshHjLE9DdVcQu59TQlNPYB4t/J8jnj/tHY8hQVGsWU9+Q6csID91sOHO
6bYuJRDbtjN/zLMNhGotO1uSSSHPvgdDJhiM2Beu7xKLEUZMI2tX++7ase7FV3yK
6h2nHhUzSxaNv53veGka+OFGQmaCT6qspL/+TtpC1rAFxkeEFQP/DB5g6zeb2242
vTe3KIFsw9TSORKn2PMEQymcsVX5WzwE9kE9UUYBSWv8jGNbHX8Gip7Y+vnXBKVi
WMtABlviFnUb3JeaeadbUmqxYVCsCk4MBskXJmm0Ck30Yx/fC+8dSaSdinsea50M
zAffSW8weqPeAPqcQnO76YLXfjsyK1hlUlF62DvZSge0F9qOtVgJC9d6z1yBipD1
J4fobeHGAz4fzwK/jgDAu+8xxG6+eeCT3lnjpwRNQLHcFdpLdfJg4sr2CVJWGmjh
0gtWxdOF7+bad10yy/uYQVE1r/BUMzlrMouF3iI/U/nTRSj/U7FSNQjXsW6Zn+HQ
PcM+FvxkKu16zdd5LjouyEI+PbnWLuOWTgwD+x2X1Wz8kS7o7RtEgHbAnRHMLHE0
AY7NZW+/QHT84phtbHTTCR0y1kBLp4fZ5m+NIXhJbFHr/LGngZXjt9NnjR2dyx2n
keWgnlsrK93LRdcGez/YuY7af78C79pu/Tg8jvcngwd7VAnmb6yt7wPWJBY/8bXH
4JWaV+S6W+M15v3ofjLLgFpnM9uxvGJ3kzeRy4Uwv+hCT7W8B8c99vuEwF1PZ9pt
edTxJ2tUufLKqII4unvhdl878TdxQht8qJOIfhgcrOW253bTeryiHrQ1Kk+gbIuE
Ezq/anOW7qSzaTwude0/yVF3PRnlgzQXgJFgORBAZ0ud36pzCtiBknBLWqLTK5Xj
TydEQ9C+6g6MfMITWc8azXSpUdjXtOeAx0q4Rz5/OAg/zv/JqIyq9ezthYyV/Q4J
3q1rYQuGnL6zIcaW2XB4HYrbpB8CrDdIsEpzvwbgbO5J9gjGbaOUnPVc7LKapNIQ
pAuA14BcL3lNEUKpQXxYRmP1/M0m4G4rN+E9PNHfxzrNlKr/f/X7PrFUkYedk0XT
SDBrT8Hz0dak+Dna0CUVToIZdq1BWxeB5SIQsurgguWQSnRIx2vQTFRKRfiAz+yc
6BbVB5fzFRniiAAQ0o7jh0wZducpDMux/4Df3Hduu1WcLwG6tONnj4yV4JGQpmYb
BEktOX6zpFI9GzdVXtDM+9V46Bmqm/1IfKKKmlJ/7JeZ4yPazqTupE1UmREKrZzs
34bDsZwKY7RPkKvxqI6d8v1cmdbeE+EF1Hh0HiDsk475IcXu2XhgbHnnNRHLGrGo
k1wn8sjw/LfhlwRBCHJ9FQQLC6gsFtqTtYd25SEY7FkFXP0o+rNQuBEIkcGMm+wd
LPHd83u5GfZf+kq2nrA2GpZGt2EM3tQsJUCL+cpZh+5DFo1CYFy5sGDFde8mVSjV
hWihLLFHsurTbZs7gwABu4J1yI7w8J69PbeY9hMv0jCsZPv26Ngu1Vg+6fwZkur5
9x0odwQqNoARvQp5FViPz6yG11y2BwGJ8jBwggYp1mqo6oAdlXVLJnZkH3XvZllM
J9o6r7ww4D42rDQTgArntiAL5sUF++/yzGAmdLIjKSbSxEsDH72DTa1f8QfthvdJ
FuDArA77/P+6gkx3kLK1qg2isDBQkVA1yaCGB+VgKdnDUxT/5OyE1Ux6QfoT+wd9
3Spbf4iKwYmLxx18S98oAnyIMtTQs/wgalLzas9uJeHAu1mB1EuRq0DW47tYyqlb
pS+4y4zz2NZO9DX7XfPuFJsozhoJRvtsV6S5yGo5WGDblumZurcQhFXK85MP52W1
WA7mZKDAqgI9ZfjbyzjrbEKl2bhPlnaQWGPAYRgyrPOXl+/NqWvjh1Gc5gnGqMqZ
ujwjxpJLi2fx0Z9GGsQ5SfUH5K05TtuCqCVDWrYH2kr1TKEMrV46cE0O+a4J681V
LB8CXj4gGS7aNIiA55Jx7LqbcRlhbhF6GO3UFm+5Utg3uyKNMvL44fQmNBn5Bn8s
3MoDHnph3sqdnh31RF0x7Ghs+L1DVCYXUVUW+oJXBcDnTtKOGjfcQLKHlLaJJq/T
WB4zIC+LxWKyf+EPWP4GvA7UksnGdguWgrFXCR8ugefVTxdHY5CxTAsqPh7Us/S1
DAuAvckJjtQJGqB36GSOpApp856MK4CXSzhoB27KTPDCfqOJQGA3W7/Z7//TXHS/
dERwcMwH0g2hBDfNFQF8+EB/fhFwvjQ/8et/WV0xViQ=
`protect end_protected