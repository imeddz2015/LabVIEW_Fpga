`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 57136 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/9huKRhRMtvnNqb3Z+UU7TahEoHV+T8U3P3ufru7l1O
3DlgtZzb9QxCbOjthp9+wDkjygH0eUfDrEl1ovhZG620gPX///imeIN817GMKyl/
KQr6k8KuqWjJdubusSA1BYkTQ9SGJmiomvTEif7lFp1UNVBp7VtrDEvPAecjoTtl
fgKSS8czeC2p4dUD9yCuyXLIYlh5UDsm7AyqqIADVqS5BdcYul0rmiZI8Nztz8XL
O7B08QYXhGZTxEEZG7d4iCDNzX0w+i6SWi9/fDuWHq65rNh1I8HHmz2Wg2S0Dv+8
Ckw9A3FxQWAWKGpoq7G8zp3ac53/ZAW+vHqqR/+Ow+RodnMYn6icpQTyjJnRsx9V
86V22w97W10oVQ6u8qCUgaPEN5r/HXcfw0NGC8gqG75/h9A79iSWW2cTnR3V2Q3H
c4QutqbkXPo5v831m8i7Po5JHTdr4c2D9PbN+IGfOlJjP6yCm9NwYR8p+c7ZkM0L
V1VK6b6AXyUSYULSpKrcwed13xf8eqiOW8JEuo6Y0Wjv73pO/ZpGQWmak3paHmkC
rSoAfrJM+ISga6yiQD5FvIzrgRiyxNE19EimP88DxoBCukeHF4Dgmv29xGol594u
scl8x+IHUAN1+zxiXhS1OWNiSTowZtKYhcJAcUVoQeRGOZE1VkOckIBoJbu/cl/v
PiBuUGY/UTc2g+r6XfRdPjCxvcgxW6kWMO1J6hZq9IfM/5NrrSrlKD0jzqYpFpub
gQyOUPMQ/NitrhAkd98bdjvuXvSS+pKQR7ZWm4MK6CbM9mZxpaPR2zPUwoj5LFmP
TFovqqgyawBeBW0izG35qvS0iuA8EGk2cCOQWs8r95rNYOK19dplJ7qaqfhugccM
wywq1glafGsdmc6ELCpHX5Tn3SfEyVee7uXitHvLw0FmabgYpdLaRfOQpeSANN6C
hLK/G6PLSAU16xz/Y2ARk7hSIMlnlouOqnS3z/ZU/qvATkIioM2KJ8R+GWHaW0yd
xGwMMxcLaOlS+pHsS4PwCrScUx2RS9232BZuRxrOJLtd2qIyTElrjK+/kdSzrkwx
v6TPlMgCOHbuQ73QbOCTBljrSQwEDCo1sooEX0+YRJP/Bqi7uJi7FSnxfb2mfBzi
RD9QAXfRxQ/2LOZkm2ZANz5E5EHhqz0ArBjbySs2rCxJ8n949B2nUXgiY9O5qX6e
i257g2d0+Ww4DizFamr6bPgWanlg0n4qgQdgeoHpI8kQN1iO2rRJvQg+5b8yYLti
kMF7SDKXS89Rc5jy3/ZpT4UdqwVShHbv0n2ltkg+rhti1hqxh2y9/GrSV2GDVwOo
pnDMOih/ROLc/RZ/QENdwLbb9DkoVPAik5bU+vkbxMyxRiS1wJgF/Scy3AHZ7Ui6
04Xn9Zad1/b9auCJyqIdwpXi10KRkI7vBt4VflOG5AO5R695+ofWGLYa3nDWqUtd
mXOnLUUCZ0O78C6Jd0WkRLKxFnWumOxnBAdVzR/Z4amPamgKWoZ2uHvPcbTlmXQO
BDviRm9eiutwO7khb+lpXEOKP0ZKu6poYDCw8VBhRCIk0GFc0UVloiUqgnXjosvM
8Kel/JoViBJsHIv5YpRMBi4+Jl9cb8CBnEgN79Bw+U3xrmddDY0pbcBWk1SfEgyt
+LgECgEsym85eERPjYEZLa0QgAIDLYVQ9hT1oVpTcTKAn0625/BYehb5GmdOuTVn
Puja7Jqn7vu002a8TZMyx1i06SJbAvyVZBzZ7dwKVdekiCP0imal0uWtiDftOT9h
4VJpPd1ajUxpBlTFgtzxf7DPMtMCs4XNzkI3uuDFc4cO8F0rUDUnPu8mQBd7woDi
GXFhYnxOcOBmPCD05YY8txSmipE8JgSdZtFGwFesh2JiMdh9DtRz+WG51z5BMT31
h5p1rS9E3PxIpBKzScCeu9Ms9pv1w4BBYb6TR4vKpGhsOFT3t2gu6elNFeYKPqs7
QvncMFV0wgVJ8d1hVEQsPhil0pbIGUVO5jyOBPZTtBMfmYvxASiOjIrrWseupjTy
zJXA+WNp+3hB/e4SJ8mtxJsjZaPiIaRQrMxIMygfgHdjbPbfc27PFnZnYZeH1njy
LH/CsvjVQe7vF9R9Ijqd+od3rcZj+8CAGs4yLtPa6MNYz9zFypQwR8T5QeMfoSM9
0URWCcU5Np+JaLsNaSn36sqtXDYUdE2kKlUFs08pbxnK+QuK8VV83zK/C4aixUr8
bEslJIDHTC4uU7FodydiBoe3bg99wblFFmcwU1BJrs7jRyGTC9xTYlT0wro0+Vf+
ooRexjU82OBD0obsavrW+dEiJBf5uS7W+FJZ1i2pBFc+sldy9ypBKJOb3rjcvGSH
4L2ZsHBexbEYgYTZg466P177lRqBRhoU3FPUdHQByN5Sb8OU9wfaV4Gn4lUYXkqV
3gfka52SguCNpQyLoPUd4UOPu/nlRJiUIur6hGdRkGmA7J9CTGiuiQl5YMhPvy5d
Bpecu3inwfu54jcXcEAs/xGmCxBCr7irETi/tWxifIemO0AkZYxjEy6z18ioDp3Z
ak7ZXhp1qz8f46t55MlYUM/rZFHq6aQntwNU019lIyVzqACxFp/SMUSOs0bSZ4d5
+4pNPHtZCx3jzAglEsBbwrTlKNKqraz92RLg8QmfDLquFsjqNTccFPcwMTq+o7Pn
7Y2hKQQA1cyzKt/oEgOXWCRN41p5nrihzgVc7ZnBfwpsYuUVAk7cqgcJGXkjxF3k
Fnhh+JdIZcVwDNQYV8lGWAYl3BPShueBvwn/AnM7B1xPpQmlAfnZ1p954LO75Lu+
4n7LsDwMTjCjpvqBApOybVY59dwRwYfUi7wTPBN9ibm4/zrX1bu/wQf1fLhg7tt/
Kype9O7e9IzNw05qAFFia6S/Zsg/GVyeY0RX+fbaYf1x6QIiFDW9wkxae3A/ipIe
T7UvSMIujMP4ppTgISyNOg3OiOqN3OAGudJ98u5KYv2VJdyrvAQhIt093UU3tOv/
tPlI5wdW59p0fPmk0a48gepl6ST2jdarZyrapX2oS0aGoVYeCGZna3TOPyz0AyBo
GFaJiIA+U51vrkKIpIjLVyOivmr6PRDM+KnSNtEAe1R3HrGrDSeRG/Lw3CFrM/fW
L/p5Vg3FW1uF7laOfT1z1xAsIlo7rKl1XsqwAyWR7M035/j99uleJUR0ttjCyjsn
rCAHKZbNGR5oWah9IhQ8zhKld+fBZWVcJk4bRIFjBPwyDEsnfJ6G1BKjfGGVQmOs
pOcNRucNc7Zi3YNhSHzKY3GRw4R1ey6C8WZ5YArZoazKLROximcYjQIN83HoKU1B
d9Hr4UkjjAL4mt8FWZnFmXTSJg3CM5el6b5xqyrg3fOUQSJ6A8I6vMnPHDhKFVpA
vW7hqJqVXGFwjFd1LhEtNu+yLvsxvUOfH2ritOA4u9k/rhREdP0Ik0sTzH1pRwIG
Gl1v7imtmnAvJzf6ZSgvOSPnepGmR7jLpXNvjPHa905aTwXggUx4gsmSOIlda5M7
0BSDH69iqC7gLvwnSOpUq1HELH6T7WW6Uyg9zCqT5eH3vXv8vcDaYkNJL4RjfTxh
Oeuo4xSfjLyn97xFisrR++wQsBG1s/j0KUYlvXr+z69YgQM07M2kQOU2j9U827Uw
Asy2fOgfqFuERQ2Dt7MBsXGgSzm2cnprDkc4eYtY4zwz1K5GxbZ60yYqKvPAndX2
EfwkxAK+ZGs34MBW/aQRMwQjuabBD3R+YNBR6sI3TGwV0Bd7OABzgPzNLICPgpWa
dFLmgbOjJfrsweX46lTbe1SoWP/nSmxk79Y0lTdNePlMOJASYgyTmZEgnWGIpgRd
wACtEH2Kr8qJrHNYPbtjxUCX3LPFjWjLcKy9AcadiJg0TYlbzVE25CmnizhnM6zu
6b9WbBZglimuQSJbmLZYjDpv3nswlF0LU5+bID+zLB0aw2+jgptbUXiapaVB1v+B
wCcXBhwmLGchM50cV7SpOjRXQDePuZMBNZDZJ9Idm47XI4XOvNcWB2Ofrjor8kdV
6InAqGyEiD7itSeqyCZJjCKUShA/WHS1o/ydq7n+0FUqo7xoCyx7QGNc7bRikC4s
Nuu/j72G40W2ggT03bhE3P0tcQIs/v0hGnZC3hOnQ4kd4k8q1GfF4NAPSFNAmoRk
ZUz1I68PrQHEvSFzI89Bl33mBMRgJFefdvgklhVGYO1UD4UZUeBYuuTOKG3LeAqQ
ldcc7UH13/NXr7+9weBH7i1b5NU2SJd3rCM2dfxx5TV0KCi3prOvtC9xoHZXNDgN
IzEfl8iqDAVcA9mQckZdRJZ3/IITrVl7ZZjqsrADhnbHPo4naISW47Wr+Ksn5k69
RhoPBfoZ/v4mC4/26ZO1qNLprENukexfCEOih0WqrcIy4Ilap8aKKrLMQhP515Pt
n++zUBJYTdB/ROZHdHemuyWoQ4rXmkGPKXo10qMztxMteKnEblRE5MbyXQk95rd+
1cY25VgINpz62yfXMO702TQKo5exevHXexVgsZ5N/Bgl9iP1mhgwxXHrhk9CkvtG
ucuyjLX50Hqmk0DY4RFMy+iRloIRH14UnkBsVQ+rRLgEXOIXTk0NL25SoqIj2ERr
flrLChJ4+eTiAGx5Da9YOmfKJAoBl5MZM6bB7Evj+EDdzfAiupS5yO05ChBc4ky1
bcRmbdw3qpFYVSk2hIc56ZhDsFGm2zMKRdIHtHvRBcu1BmPRNChVkRjE+XhMlq5b
jg5K+eRREVIaxSuLnw54xV+ggjxKVAfMyEpA2lfGO53jUHAUnpR8uqpza5NufB1Y
SKYy4zMH9RzEtj1t4ZEh188mV4pntllI8fO4y61nyWiGioWqKo7hOkFeAlowBl15
llPbiHIqvfHgJvvyQj97ZJoEC0X2rPqXjO8SsZSDcjxgdog8EUYf8oV44ClLMGF5
87dyhfguHe6NwfTnttMHU11zW0TbOXXDfkW6nJ0DM2eGmSiC2jZfnJAStgS8ZOPR
adZeoZQViQQOmvtg/vrDBTDAHjsPzBPXolxLab54WUok5PAKyjiBA6bVgVLSa25Z
GyigAxJXbUkiywAd5TiHFedadMtdKUzLQxKI1aETfW0UQWMBpgfoQ5SKEodOjH+3
Bk7avlpDluTt6XD6ua4Tq4ajKuzzgwZkcBXSxcLg03q3mkKPG2E75Z1i2eB7/u7J
Ke3zf4GGGuKgH/Edp5JDpcgyGearlAk9hy3tummR8ElZi10URON55RC/20gQJXal
M7zLXkdH/3b61fUvDlsSKh1j5yYdeJ3bZrWFdCoibaMaU86nIqBeyOnz+tpT6vCw
r4alTiAHVd3jEkaH9vp/77VPHQb8ufcm9YBSzjXnOa1+79l7Q+2mxARU85EGdiYZ
PWPevaraIx/Fgwa3wViDKTwtewp5EnWf5gPplNfve8U8oppDwnXZ1pI90C0b3+5P
lHpDDtQPjUlNoAofaqmO74VdXF7eh6SDHy64Q9xYG/Xbhp5eec37keHcMLOGEs47
GnrlTWnRZAOmu+cjhm9UcbHOeQR3j1Xs409b0aiobPP9RqzBWll6uZ6yJy7SPyuM
bKzPOgBYG7mwQ3R3HHTxi4FijBhq9H2aSgpfp+m35WEx/+gPfXXxAWSoZVOYhnkB
JYpW+W0NstEi3CP5Kqo840iLw0P1R3Ehwp25ZUm9KPOWlwycbN1O8zSZgX6wmyTV
WHhdY+RdbuMPGIsTVvWAqA0rGCxS3z1WrrDVZy8VN6rHRITUsoZeDCT2T8khY5Hq
MzKdiY0DI3/EATWD8iA5pi18YyRdn2w4r/vgzFF5fw2B9grn1fwZFIi2pLBmdWXJ
ixllu6p6Gwpui9J8aWz7Tmr/rUthXUVyZ4Rcg8jqqb9lxQHALB+1Y0rmQ5vm093Y
gn/XoryuGQNl8wusTR/yKkk6ZyfmEo6xTKbarbKukFIhR6YwCbBmm2QHdMpryERz
APJHnn81VY3KS+c+SChJ4UPsivZIhDPs64Rg8ePJl7zNKOxw9R57N8oWNZp57Tpu
QFIGL4KvHUDSG/U/oN8pPjBc6WxXEMZZc/0Q6vonol3YqcSVEqb7U4YN4VafkbZr
GIcypbbK2MAKV4dvPClxBXlOuMwHS//120rNFsGfOnBnk5wOb7Qa49LDxTlkO8Ga
khM9uxSjpw8/v5p8iHYuAOcYjRmmNWzet80VHoOYfmGLlE9Tww0QW26x+fE5ewXv
T+IgL5gg6qOs87B328Aggd1teaCx0nAt5jIqP+CDNmjnhNjnraPh5wQantEgXToQ
edp34i/xD95yxZxZ6QVJX5lhqQjVnG1YlX0ADvN/x2kt9X94W1IHi6DL3CUUqEMJ
aRZ5uXNRP6oNJKeENak/bryP1IXILfH3oAb3LoIJTQIgMJkU3blqfHRL7qRzuGOf
9VeA5XSB5aYxLDXLsctz8BRPGRuJwj+y5EtbmSEa4HIbG/tXRO+I35bePi4fClvl
+f2EYtko4pmUYIrLxyIWlXd+mK/xDwH1S1jnC/TU0PstkR8DuFR4xE5Kftvfy/7y
wc0rxhWFb7rYrMNIq3fZ2dheyF80G8LNXm+sw0nSZGX52b7dtSYXe7TOzgjNzBFX
jHWb6z0jFdKh2Zw8/uvaqcNiv3p+7pi9V3sY16QRxIh4X/LDkOlI/G55Zaya8kby
1flmdrkLSbLf5qZ0cKcpIKXQy2B9OhY2cHQxAQvcRujLL1FV6WSqKYXjRD/GBAoC
ZqanAUWPdZDKHAlgdTkyEw5f6HtJcYps3F1DeQB2GJOqg6lxp2YotlHsKBv61IDU
zVoI9rnS0pQcpN3+NFTNCH3sYRPrPH2KWIo80imOJNOz4BTsNblmEDutBXR4Yg32
7rbTBLBNWFrZiDJqMP1AGvmJYzK7eTfdbNd5stbz6jIL6rjTbu2O3WUijpou/5q6
7ov9VEpcc62y4nVwaxNs5I+lx7wiu0edXKRupGxQElQKIDlgCuTILnJFrmfXcqoo
N3GyZQ5Kzmzgi1ScQp+pRaxNuZR4hXE9EAqsO8eHNLv6VesD9cGxx2clqVcCxWVF
UkhPG9RR34bPlINSd/RD8BnDBbpUwgXhpbfOr/uqkW+LH7uHNw3l3+0d51F5/AgA
Cp0pqy8pF9Ir7/pNatT+lEGBUuYvn9BJ6rYoFve7JgRxVwD3bkByd3K4fMDqzfhl
Iv6APTQKDOShbUzMDSZ85J4KvS4nTCY4HxQsxbz07PAmaMYeAjxqyUg8T2WaFPi0
evzn0pSjXCNg7hnKI6XLn5H4DI+sCR0KoNJ11H7nkqvpeZHJY/O9gTemOCio9IO8
xnxBN4iNRaY0sea+qsSaXEdhQ1rLiAo7EjM0gqr9yMWI04LfW1gm5u1q7PtwJkqr
dXXnsMam9U8B8BAnWzqshhoIuKX4HHX8UaGDB2RYo8FV4/KIONp0Tv49ocv8RXov
7l2iXugLD+qhgKCH7zW2ltvhIMvYbefrEM5hJZ3nxGXmrOVg+CyeijKvAWIYyJNj
qFQTmT1fWUKFICvcmLlzlwYgZHL8DkCiz+g4FAUjoiJrvAp19/C6UfBsDLjFkLL9
oBz3pY+P0u/GHBz1tgvHtjiA8AteN+SGcI/E70rMAZlg46DYZy9Fzc1M+Y18oTMW
aojTUGwAzW6PrqFi8bWn6l5LgKBqAOcFOn+DIOydOVhK5/6E/C/v+M4tc0L248Ee
Y2bRzIE6MOxfGKVFDWNbvU+BSyflO/EHkVJnL3Q6FJt0Poh9KwZwHXgERTLbQJ02
SP3LZ0+VpKXl8Kl27DtFlNHw4x3kmVfEwczj0e5bMInSg8cFLzjY1j3daMRmEcjG
B+Yd0TIo+VHiekILmNrXF/IKZzEoU1mxC1WOyZUV/7PnnuOJCPuF9zxnQ5r7imI+
IX187tvPiCSgvFEnVwk9RBqTlsFSB7hr5fC5x7vpM7mCSEugIDV8d5lT8/x49wRd
709R15TpS5eeeABjCP9wViHPPxoFlS6mCwGSNNPi9fnANOPGWr4mOpIVrOShZ7yM
T07ihrImo5LaBZ0LoOjkHtJ2PqDqYFOx78U8VpWka+9OOHRTit2mOsUccAR7PU7Y
uIRhvKpWcJCmvo1iWnsrfSRHjYvOCgMN4qra+MOTa1i+0XpvY+AN0Deu3pFZbmpF
EcvOxP51apYwF1W8hHRI3q8hKTjVO1iJI6q+Q4MNocRB2/28whQr5NcxqMZ2nDAb
TxLk1fKTy922SBj+4AbJ6mJPWT14eQcTuBvTbUNWqLg6ehK0BFxc7XPmqnUYW8BB
GG+WWQoWPXJUMEH22h2A+sQepCGslckCpbhepr+EZAOudermCRG9yNYwC9E49KBx
OhZJHq7XNkX3vZ/cjrLR9hpnwSnsFYqsFt+4gviOIiAQa3f21NC4oLl7z5AZkfdI
X03w5zyxMHGclx5iKEEOidlzAbnTkEtRBz/ROplq1bQSz84s9kkl96KFDPdUE+BQ
6vgi8a7fXpRe36yQtCOKZ60riu64yRVMu4ORAuHeuCT+Bo/ymWQntSMn0C0lxwon
xWBst111Fo43jwBkNDFclrvdbSYTaBNz9Iz33mjMvNjcP9ix8pAixqq6AakkPvN4
l0T5ufyFaoho19q3L1o/7f6yrlOH1inK7DFmagMAv7gqKu7CGvp1U5G281IPOwfR
WoFB0V3JPeEaTJVXLwv0s49P1GLfJCwA1bXo/ArbsaZsDQXDSUYialPhvQphz+E5
TIk0KVaqQcHV133DXGeUdKeR+dY+eimDhPQ1tY3T0Y8uMy65X4XkFWPWfqe41hwJ
tGOGNvP70QyPrzuMFQuOVV9oVYONWX6IMIOci7LYHlgXvmPCxkG+SSARMFkL5jGM
D/BskYYlAAyXAs3lHecTO7iy2ts7Dpm9Yjn0sskRgQCGm4lvj6gVZwE9NgiNStzs
qOdpRp02c5m6VkCt+XptjaBmIZFM456F737892CjWnbUFNVodaUO3VBF+yheMvin
D/ckta/SDzQSYiufCDTpVoZVA5qE1uv7sZh/tPlMvYhuUS4oMyZSVegtyT9p3rI7
bIJauAsFojcju08VyNtLS8RU4jKXHeg+uLk9VAYN0nTgW3sAYOM4DNprA21IRHQT
2MlFN91Ez6Rc6Ebo7k6unaFoek3cHM8kuQfihSO8lg12PXUz+/JBvojmlYf1HQl+
yAvfRmKO6B2fYXYIP5wiYKo8FvnQv1Swrx9TV0Qu6qjgtAbP7mU269T796APLm0u
Yd3yWVvTKyNnyJq7XalXT7+u8gTGMhMYd2H/Qx5PXGcT1HJUj7Vf0fKI8kfKxVmg
rsyOE7+bPv2yJUR/oK9f3C07ahLzSi0hQNRTBpR6/ODkjsaa+QAq9j8SzWi+D1Nt
m5jjj01ODZeK///XKuWSXn/TSrUhAqnvzGtLdN9hkz0+Lkk2/IEPjl1AOVgs29z/
sAPueXC/UoRUMKM019GJn0QtkHiTchMUzKv3RkFztKiApAY9fhbuUiqLh3xpaevR
z6J6DBFsJ7nCaBAB8q5SX1NiofSmdz+hdUgKmyrWYp1FVVtdw4fWxZGY1nNQ553l
TFKcD6pHPGF+RWT4MvJRPAS4ZlpenaglzewF0RbhJAKwHBVbHKMNPMXkGpOkJIlS
1FHRlHxGoJA6GS+i1xesy6dk2ASIIJBmpM/QwIIfeALVkpRnaswWRl4wVXEdKQsK
ha8f//aPRSbmxE4l8+wyEp0VHPOL8xSUTNjAnyQgrDEhCxf2r5qswmVFpThe935f
7TsMjIb/OIJIy3f+gL0/UlGzmpT/y/wPhWmSzUFdEPPhOPWuW9jJqawILBYhWLJq
uu654rMM38S58CrNbV2qmdKA/TfGNoiLTsPDdi7yxIxv0ilelL7sUSTN4h+srRne
XJtpV4C/AHb9bDQXL8SVpZFcsIVkNlPujLZvKNBrD4QWj7vTBG+Qc/AelWnilfto
H2ubfmjMdyhaze5r6um8OtcFglJmz3WrJ3Q06AA607wpN3m6x4XdXlVLvJIR3bxj
SYc7uT6P3AsQi2fGysykOJkHeJ7kxvc2M4/A1qS0THRNn0VtKKOYBE4elmE89sV3
PI2tB5LJ6ElqNYj90UUuy/HbflMuKUMLNOLzjw03mrEicLbjmtuX63NsILdtXh4e
9eysGlOxpUTBzqtgFA90p3qUe4R5WE54hDndq1Zkp7cfaKy671ZSR158ZWWtLkAs
YLb7fxnc0TOhyqUJ/idT5uaSf6zYJS/4FOv6mZyBCLDq5V2nv8rsHKn7vL4zcrcb
AEVIN9y+5I/VXo3tLbfk4Fr7DQ7moYb7HkJFWJda7nd0lXQJdNkZBDJIhEMrw8TD
OSvwoR1/PuzEz5YX8LRWxZ5P86SaFI1u4XYRY3s6UTlra1GiLlcwuwS6+9hTiKbJ
fvRS3zQdnIvC71KIgFfY0+Tx7Q5V9um0aEncpGrzQhUb30Hc1psvexRtLXYoxace
hf1oeglEpgLL//iCq7S3bihMEAwi1so+pYAUOaCXpAfKUp6hTeev4T6FxTDPCbvC
BIoUFkDmah4fj/kt9Uk7J3MgEj/qup5ULPRqtFD+VQdhGvVUD2ZIacTJnk0oPcKj
RmjSAs04CAN+uj/Q9tfBGWGoxXjXsJSA3klGw/0ViUD8/z9so1A8alEyq3LfEBQa
1CHnPGCqDq8i+/4hZZk2SkN2VoKmmxZtqHVFowPuDzudoPB4TiKtaID6XeLbGnBz
r/4KBp/ZUW0zHhSfu0Qb7bLj6aVDZYH2CQ6kQMvXqz43yionigG5K3f3GqFxF7MX
ryIazUQB+VtVYyM9Km6E2Q5/Rm/TCqyIPOl4IVz4bNOFmRVQKyHVUQb9L3GwUW+g
oyxf2X7cXVdlgvyoNL9glS7ZMJ8dyGabcuuehcZuDxa+S4Z0m6UqSVs4RJI8O19B
DKtU9eRsrrf/lf5rkg/OxUhj4GzsXYnZS3pgBIv+rd85jI6D4rEeTVmm+30YiTnD
AZv2H2QX6AZ59TXH3DTSUO3RldikLrcF9d9ZRhn3tyqnPPq75LMhtjPd8C8Ga1WN
2AC4PUggSDKKhpvLFMOWU7rmduc2DpoAJWhf3qfNT5KmEHzaZbGhVHVo9UyggLCS
kxZeAAdr4KxbqznUofDrfN2/dzMOgZ+7EZ1Yg4AOI9bfLhvNuN40MSRePu1ij0/m
mickfC0NIEWZ7P7yIHeYfqzDNvGVRTakQovxdkT9YStdxNGPoQtJ+wCOgkyCCHrI
9npJL7rqcWrp5lw2Gi08wsEkPkokeG4PFNL1BDRqAVL/8WMy8fGVKy7tFg5g6Xv6
eCP9AM99EGhdKHI+AAAKdtSACm3/Fsi//hFSwTaXA3GVlGF6eTa0r22w5/Uei7vm
S2m7gPDbccpGI1ku1SKoWwBIcEOleZwQPISWFNPN1IeHhCO1ZVxrgZ+LsuAkOmWJ
YrKHcJRCcr/9NFH2XoP2GKEjAR10Oo27cZdSrRii4ChP2j/YFSHOnQxKCHp5ya6P
X5qWSRaE0Lb/3zP+VWPxTx8JIvF1XwHJpQODy2mI6ZCF1VJ5LAjuOIJ25g8nzEse
ve19twIPEXcgnad/cohNWESZR0MffDDnmAqKHONc3Pc7btkFpDIlTZ2dlZxeLI0t
/Jh3NG9uCxci5sjWb0zjg+9UaeQGKe8f+14dnZFSfm0cTUOUq06BMs7uE4qw/iSu
I+w4ws9BTI48Ym5T0WLUvVuco2vzhpbfiGwpEKulYA8AyZ4krk9QVmvCVWyHvOmq
Ocev/xTRCTTBqzlQkXqpuuDAREewy2VR6oNJrnpc7u8qGtBN+TW+3rheuY/Ibalu
RZ6qgC+iwkLAlG2m93ROwcK8hzqJpeiEKAXVvH89IIty5FdMEqsxgnaU/bVYodd7
o/cB+LngvqRwk69ReNpf0lyFI51ykYTBVnwq8TsNJSawruC+NHfKxcZe1bj9YCre
L4gsnoCsPIKoW9RLJjV/vMsrKhokWl1Jf0IcFzX2suZ6RWWG7FUkoyHp7F9h1qaG
mR5W92MLlOw+qJroNgGKV6BYsf46pNbXqzaBgWOjXPwHyvvxrdNDcLbfj7NXMeYG
AHHrxhoYt4Z1OVR3cgQOWH84VJfAvJXnVhggU4QMVs6loldJxM5pB8I181L6qUA0
DmidvUZAiS1dJRysR9ZzpHv3pSMviNvcrto5XmcCpfJjmPpBW99xG9tl2tl6DY2R
MWDUJLSMrjeWzWiudGimSVGBoXuia82GXIrztIW/MSShq9Myq4BUOtKJQM7GJ7G3
3PVW8olEkEQITpHjFS492Fs2HwdQUfK6pVAALjz8qdmlLSMrRzVVhmnMfMTTCWMi
PggjDdVt7guuYsL/+AkDat2y5hnjYxHFf7PZDxLOcvAxJHaee7+HC7qNOwEsEIc6
CXMcLTsbywUl/c55fsdDpx7xb/4kdW/UjAhKqTk/i+VCtC9o5tP/5csQZ/KjO1uB
/paILoUBqNv3k57raNTCpkiQ8M/Nx3atxlbk1QRf+Sn/gViCkgDcxaeeM/4vha7Y
f+sqqQuWMQZOaATjzIoVL3IZvVzxPWc7U5CxBAhMCT2C+WV73BX0JGLuAi9IA/Jf
G0jVv1Clu5tMZ6ChSqmz7c1WLGSw50RrNbDcS3E4xvzfuhdezoEJMJohFZtiqjMh
sG8GNVHtu83AnYCcVQ/WwxYhJDo5vAe6xyf7Az/+uKuppatszSIROdqUBxTKx2v5
/gqcuspLyqCDMImzf3B8+X9eZYiggg87hdYB4Srw8t4ftX3qPEycVChzYiHJyrvI
H5E8UGbSelV6Cl1XZqm/9RTntQgeFH9uNFcFTPMcq3nIOKScVgvE8N5sK6YDpCfL
Wtkq0VZJgS//fdIKV3dOqLW5DcT+OA+ywuBIvrLqDhH28ZGjkDM4usexjclSqB13
e0MuuvMITdq1YTfwe8AJ5oQu/785GMC0P5b6t7X0Z36/RJyHG/6VLlaHH+33a3bm
1P2REwIjUYxlLO0RBBxVzjKI7Q1VN6xvs6OGW0BV2ujwIVgNkC0966Hs2pTPkmOM
RU+HiUHFK2fxhgXkUXQz77dGSl72Y/VE2sB9+GVy6abtlebIsq060XzDKn60KdfE
7/a/v9l9W82T2qKDojYcBDCwTYEdU8YXEHm/MClO7Rc7gGY+2WCcrz+I2XeaqwQr
J3fU+zpWU24vCqVHbaSuEVyNWM6M5OoKyvNrTtVSdsJMthTdhstCTfwVsoM8j6eH
RIW/VF9/PczBFMY+ECsacqs9b9dSjKw24oGJCgrIDvzZVD05bz3TNKRQGekAygOT
k846RFiHwkipnz+cQayqcvF9FDEj16lWBxBaVX9kaz03VcMjHGrEokTgaYCU9c4A
pC+Reip3NUMAKsmPPSv7Zrjwt33pctN6qXr+47v0nKXhU6zvSctPW6BXlXGRcOoF
vHyn2IYV4/jWtrPBJ17i2oFgtXJ+liXz36v45Te2KWlH69Ifxr/Y37pAwZSF5G8o
lDMPUgDV0e5NVQWEhWj0ikI960uqXU2ACUixgkxO0EdrVuMK3KmYeNO92VVXPLoO
8nw7BEtRoe1m1vU+e95n7AjZPiXjwhAWqwi5iQ+sQGlqJab9x9UfGOXM0VQPaQM3
MO1F70NKEk9w0Stg7oB0lrsWmLkALDdpzbASxBIDzGk7VaH8iUi/743emNZM5XZR
cpvqiMb+oU/rHJDEoE5nJ7nk3XGlXXYjmS5p1dKfOhr/ue5avEBBkFVs1DPz/3hk
SxIsDx5zO1dKUHKLxjLyofYGAvrXcCbii+/Jb8gFxLbfnBFII0NcwWTAqh6Yn/LG
WKcjN/MzyJ4/DdpgjPWKFvszd8nIadZOGGs5FrkgMAixfQu5u9xqPLBwSG++b7/U
a0mXSLVCknnK4q4RuMNmaBmeThLcKU7SpfLvP+fnEQho0fz+7MqqMo4+flcZqN9f
DImVRTPzQ9cyrbqLE6LIyE3njypNXDADVTUk2Z20QiAI6hsUJ284+zz2vCKjrxnw
7TPfe74ziMz8MNDqDMu4aN1J4EAj/d8jRNZ/LCThHHa+NJAL6/AzM+Vkbtkuaj/Q
bI6DQ0DaqwkpBdlTb6h9/iVAWpKwDnub3nBtVMl3pMTaho+D7sFEK4/XyjDUP999
7H8rzvfc9EnvtNwRkC140ygSEeP7SzIrw6IqKPevmGyzeRKV9Bwo3OhC8f/qj6GR
pDmzp9aDQ8wzLvOGGiwPGir667wHSSOvBhkGUuGG60b9PR1UZpse/OLhDK5/m4bG
oLzLY2Y0O8RLGZdn08uAVcSELwAm8NC7sYDaw5JsdvjIsj98D7IjBDVsJo/k6tTh
HMBrBRpaM7D4gY5OcjxmB+JQMQQhE44Hg7w8egKah5cUcsAjbqnvMkYS3fcoYIm9
DUhc2so5KU/QFMUEoSsaOlimMIDM7dufTkRYvca2xo90+5gxjrPkwwIW8G2xjejw
lGybHy5h2rxZizaDk2jFg0soNGSVo3pFyB+q9C2/QrmbE32llzCS4ST6w+zwmWo9
CdVI1E215xkuIgJajJ7ejcLPWYCND775UwzkTJwJSjc0xoqfqLgRvMeKfL2/sRAM
0SH+WYX5s7V/VaPYbK0XIq5ubRZzihbh5CLYcOOrZiAD70EAZYR73/euxaaRVzN1
1fd0CCNietFrfxgQS6US527G9TElNjKlJ2JVjnW2YSKdh8BTr+BnDbkUdYxyMPL/
q2mUfeKhkJIepNpV5cZMZsNdmHXDdGuFUnTS3IZzAPEPeeKl5anLokz3Aym9c0LD
2knMQIyO1MI0FBLVQkqYDXkn1IFUhWDGsRWGC0OHld5h+aOrp003SQhoBVqrtaq5
4Lhz3iyOa4r0wvXaOipHiKqeuh7TEroxDkMbcYEx9oXt7ecz+eGSQJqBHRX49t7u
M+rj6FIio63CWbtYmQPcamF7VBggK7brYoBbNx9QW8zuow78T2w8UaDEmzBs0Om7
w7LG055YkUg8NoC8im5zGjZ5kcnfXIvoUV3iPmIf9I+FPdovjiStMyEOQpS6w/GH
fnsA0KFRyZx2wyoBYMgNEWRmaqWdnk9eCprnwUQ8Ne+Xbw/5MNVV2su8cmNFOObV
m/5Xquyie50vsxsUbJhgQNdVbL18mnWQiGgwQU2T7qmo4GVJ9lPMqbwk7ydYOodW
TZCimGTO+10n0Y4CVxJdcZxa6nAtF/El4YlMcGQ5dDYWBaBU+AVkahqCoqRXMblq
pJsfPrPUPcFenU6h3/GwyjuHGCwEdaqSpslyUczpoxCWFufSf80O0bG0uzld3dBw
Mj2c31ntGP3wIFhTe/036ja/ytbRwL+zR5e9qqBSAls59bvvn3DOsqIe4yvSlQkq
gjFY9df+WYqeF8bhLlAKydobBwA0mPWkt7T6YJbE/fcBBhlmrgQ8uc5XfFG5yJw8
og4T0XxJFCgzdX/tN0IhHScZWo+lelQt/PoeIVtDiqcbHSzCBwU00sblivtx078l
kf6supXSrWv2HUisXyuN1oSYpTHvdLm+6xnIuF656+be4DXO7FxIwXZPX+jVorDA
DjAh6AqBwXKULl8v0jhtYNqg82J7ee63sW22LHHWO+5WlAL+s22CgQM1EAYG3pqd
4YRkaVHHSrsNmVcyxvWBVv74KEmuTb1RevGZZ8LZOX3UdZ2JBmcJ1tbphkx5wG7O
ebtral6KcKgQGhg3eez9N2CjeinBbGv5YzGBtcg/mdVoIeCToI9QuTb4Cla46oiP
RN9DTMgVgE8IT+zIC8UEgNb4WXdHCR1k/JJFe/L6NKmqT+OUge2CAFTInxeLbh9H
FXf1OP2d8pIG4d+HELFx7018Qgl6RSzY9q1QfNtibWgIdcwk7Keuz6f3TX+yAAMA
FJjspHF7da8YCLZXp83ptKgjqxXQN2FH7BFtMkXude6RFcNHWl4Yqre6SUnJBgMt
Uz4dpr+Oru70jdXStnO0GFXoV6Lu4i6slWR8E9zcwus4Z9KTvq6OM1wd/dSEKLtT
URdersKMG5IgDxpYgffDu79F3Y/GQpeP9vbofjFW8wLMWL50pCNaTq/cVPz4eski
FXcti/5HAvPSGgLqNLYvnQOZVBWt9VhasfGA9EtlrvrFJjJpsdHq5gNgGCoBGwfM
4NuTvXxjOeAe4KzRwnuIJSTjjN3xhLErfYHvVMShjM/Lq1SNoJR/CMjaYsN/CEaC
TK0eFynL0GUsb0az806UVfPPvLU79LhQZRQNU3CF4i8B52JRgazOpMOFD2bQeEHG
DY3+M0CaOkulALccLf8KzjjHHd8q1YWshlMG8ktYQrOi7rbnOZRIdnCCX36RBBpC
oyImsJ/VMGj7VPgTHYIETkade/fEDIZarSaswtHMcsA6iyE/C6XT/YqP+FSJkEv6
l4hS7wHFp0FbWdwIYTUdIaGMRAkm2gGS8w8dCMzVPQjPrALeFV8R2AoMbnOTcTLD
VgNW25xV46nhf/KN1PMa+SYPmNVLaaOnhSsb1BOZFvYWpDHxg18YWXtrmkoJ4miX
xqGswXVW5NnKpQ4UWSZJiRX72wp91IN4nkBWGIJBabIzQL6iN0K8SGUdQhhOnWDC
2h15DEuHhL3/VXivOHFGXWcuDUWDy4YjBbJ99FFbEdTPkeO8WoBcc75G4TcoSB/w
A38LBq7MfuzLMPUHMucGVdXeNzDCv1DO/DG/CaklMKmoF8i5zFEklmlcHo1g1tOV
CMNqCgEfQUIXfm354MN8oxzJ88DdYSDTu1evrej9mJpAF30685H5KJxre+BXu7I5
69K4deUHdZc5l8yxKFfF3VN/n2YZkGpyURA0VWB8lbYKep4NjVRJGSQNWoKOjRI6
WpTUs3oJmWV2I0NIxGVcHzRjDh+o+XGet0Q++MlLoOqPwTRr2TNPOilrOJ4bVIYj
9zZFdIWP3U2VIGHjO9n5F8dOqAPISwzXY7FdKpEQhYXGzXa6yqhUhdwaBtiqk0yU
k0UkJmCDsm0iIKrnaajXX9qC/0fcp28mSNfou5QhD2GTyv1I00RL/N+xDbDNyK9r
l91HYcCIlrLWxxvu/5K9KpvjSaDCpHbDl0Vb/fZWjZwm5NVlSE4o3FveExHnKTBi
sHm1cL2ad7Z9tMbWDx1ZEkAL5fZ5j2QCRWXJavlE5lV8AjQaVmA3pg7K5LR1+B3U
D6ZGqEJEj0ra9J4s3JqUk6Q4Bb3XSUp10rgDU1nIo5aY7xKYPiCS+YKmlBrF0f0O
KlslBi0hFzv0EGWy6RxFnEG9vrR+vkh7arCcJHxzx8A3TpfAqIEz/zOSx3sydaDB
uCnh8Vul4/7MP6E6F/yBkbfr0oG04aJGkBwO3uG/dMBgg8ETbiD9q5yJ8L6OzuLX
+6uilExnQqanV9pHGetsVH/o5K0EKYqnM5NA7WoR6SKKNspNNSQ98Ft3zh0+D/Xr
wpABt5Gr2TVpUFAgI2hdJVTIvF068xxqwLBcxunmaJrQA8eNcu7r8TCdeGgA9tnY
/IhjHGCEzc8Dr1Z4yqj6Zt3kakzyk/rT5URqny/i1k6znGLDEqshoHsgWKKSpgea
6Sq/totoN4+OBOPp9829LXKyF6ncM1cLjuZxI8WRNwunECzmt3gEfQJk0kQTCwn+
k4PEMHYKCxOyDLIQIILv4NFSFsyG/KSsTubYIomTZU0wNggBJimpejYPBDajQYtD
hFcWAvgnZOpBXKOEFJAqyOEPUrrqmilekGUrE9eK3IvIMRv6Becfom7M4NVv+/BV
hiUbckk05UVgh3pWDaeau/YkSUsQlT2kphvn4a97TKP8e2Qvtw48x5mOyB8u5mhd
XI8tXBecjKFGZPe2fPNpq8UNmV6ncUaqRlJsaQBLQTxa3m4iBtM++szTwuvu6/pc
LRm37uAbK0BdY45mxL0fOEVbAeTo0MP7EfzqR2nZc4r0a3rTLACSKBp/jq2YMgSr
K/KYnLTG39q77lU+Q59UgFpTV0IGXkJ+cJ9drWkMj3aoQHZb6n9btIxiFCjAHgLI
38M+nkqzRY1aHbLnVK8d0nfhryix+ihFa1gz6PFJ0OmwiOpxA42gp654ImkX99Gh
LIsMwoDek2Rnp84XTISZeNSwY/GWuOzACtT1s4UxkpdFtPmg+mMqeDaCGqDpYpZn
u6b1NS/h/gQwIsNWpMHufLsP1fepbtwCsw44ecrUR9PtFWl3NReHoekJqsjkxUa+
Y2ZdlsGaJRzXQtTNSfAOYVJfwppv8zPLwMoWAJ6eMZzmRCcaHENHYfa7KY2z6pQp
k5eIRSezYaWYNXgkI3I9MI5WEYf5UR3e8NFSu8LtoDYNpczQVaql9xNl844zjlM6
c+/Sh3wd6Eu6reub+o+VhfchGH6fVkG0jvvhGL/jtY/562lGzpkE7ovZwYAYLAHa
iuVnKtRuK0ExhlyhzqqdYWHLE2QFSm3d4fLmBUoyYEpxiMs3UotE0KbHMJsis7ZV
zQx6bbYtW4ZZVu8IFx8CrTaNa9M8U4xStS7Ln498InSklg8f8MM0DvVNJly/jHa6
OTYLyuL3rg/NmRAnk+a952zVslFoZkNKUpZZg7LgYoGuZIqf6zYDw563YYKJsB3k
8ha33ngNy91Fo6bOEyOd53+s65pF3vLZ2yVENNBcL2dcY4yvlaGD0nHT1A4S5R4L
BSwg2WWDpAYrTqlefi33HMML/kiIOvaig3tY5CgnV21eVAaS+tUIydkb/9XesA9O
MbxPjTJD07L4t/tlAdQ5+KECcELD0UpyWg8OAeDWbjpKdozoOUXpfJ0xwNZiuZPp
0J/R8Fzi0VXiUnVUxTcna+pQQHvbJV0UMZoqs0mPor+m1zNY7F677i275tqOVBSE
pLMo3y/0RFC15x/RQl6dhuuc583SxUai3e20UNlTR1LdwOn0rlLpZ6u4IzLY5ARY
lPNZnVFxZWSC6PxGa/9gUQ8+OtpGOQQQJh/wZDvmCIrCfJq/nnb+FQSeHP+PCG8s
3gpmk3jntK8v8bWMh3dRcwp6MHBgB64Y/UNhEMQSN8oAeYb6lvxgSVV+mFZZb3w7
Fsrp6kObfZ14WU4HlYPSPU8YrO95DciYQk9CaCCOu6XZbEAeX80NHVb3yQR+hE3r
I5iTffvHIO1dKMvKfRcg7GRBFkl1Jw8VSZEEThECS4xVCVkpaz44Hao7PfDbw0Ll
jHrIC2cIPpHY8wVbuK2adgsQs951/p+1oPwJ4Ba1cTatLW4JcDhKaxODUZBkm6Jk
KJWNwaegNM2N1yCm1WJrr7KxHH5cQw1Tf8zWZNo2NoijcLE8HR03ktH5pBpkXy/C
zWlgfQtgSJHhNj9y8Sf3NKQjfjTU4ga4V5Y9p6Rqk4m+/xBwIqm/lS1rfc9Tk/CH
pniuPSsM+eeUr6tNW9mCv3/poqVVuCajVUtgMR+ENPQcjD7Ek6svP4OpkFqFMMqO
Z8+1Zum/fAdWY6OVbnRT607mhlEB5vO6vdiKDhR2+Y5HSz9GrsZySMnZ+j4q+V4v
uuR/z7GxMhjCNtt7OWTaHss8krvv2jXwhMgre2tunr+YtQ30bV+do0JCJn0o9/hy
DAjJnpYVqEMlRcdmUeOjVt9VykSKL8329uGAgMf+RQBzPV2gmLnj7koWXCAbchZk
nPZ6urfbAwZz1LIkX/vHYZpAbIp/UiecikuY8sgLcBQUh+MVvZ63SPuvEsvygH6p
Je4J4oyV3mn1icdy8HIRqaq/VCrTEJMALHFkQtceV6pKm2pNuCanRdMYVJMo3bOO
Lzyfh0edwIWgzWBzAhMexygZCRwQs1eksxQIsggIea9IeEpJdu0c95BfMbDNchGp
dROdudHvptQZR4q59BpV+0CoeJi05cR7+svNEBtfpwjS143Tk4WkivVXIL/3LZWN
utNyUnljXAM8O0WEi+rG2lrd0mNFDytgwXoZF5kz7Lw8rN72tTl1LeKWJLnLSSLV
l1c1KJEWBqFgeMCFhjqaWHkDPBQPXPOAj9/K+vwtAwQCv7bgyR2qnftue/iMvY+v
qnDxrdcA5UshzLETt945TDHqBo5uBu1BuwsMnYNwiNgXWCVA+P0E0fzqZX203GlH
GqQy9nTG/OMz2ci0J31/gbYcV06uQ8FmWbWEDsQLd81HEOlXArkjjtld0TX57FLx
Cqp5QdZGtosQgLQqNCkPMFAp3OIrATjgBfmeplbjcKHndrmgr4DsDLQwkGPgtZBm
sr6lnrkzMXXI0rUvnb1qtHdHRKLVe2ayZpXCusskzWCyL+zzsKRxvP+d+YZ4++p7
/HtTMWOfZH58S1qOhs6o6sNzWUiZKk++SU+/yYMUuG/KouzTOTa25+6mzTp+QQdE
xs+tg53RW2Uchk7Mjyd6xnEeUuflm3LPYLgvpQ4BY3bNmwfFHwGToAm+9V4M9D9f
dA5aHk2gXbHW3cd8Ym4blBcG3dnsUwXlkO0q3UkdLKzibQbyWjBWt2UO89R9Vpvi
kTpRJcsXBOvdpYsw0PSS/q3IWNe6pMoTzsUEnTTN/HzW0bkKUgfYSBmMti/hQJw2
OhW5Lid0fqD4nTnTbsmGNpVHx5wJ/kx88+bB1DZL9/zcKp0gf7xYizo3aOzb2RqS
S5xdqHFpP9etFb95vT8WciaHb2Cp9x8GVujw9B86b6AT8pnR9w+ATfEMp5Q06F+i
IAG9LvUwq/2REqDR5XlfBY8r7Lhgbyv7OlI0lkBZQjdZR2rNm0Lj1DZdGUdwCNkF
OW+SLAqIav/P8yBGQQJubvpySyK/kYj6j1/fLD8uvNFTjbQyp/W8zkpPjqfz7iRm
CwyFg+7OtN7jpaHdWGv4GWTpxisOt9XgAYoApk/EOkRI3nfKV0pamBbob/zHZV0U
WTRj7EoS5IuwmLXM9AuhVT389J8Ht4UBt+/Eo0n0Gnzpq30ILhJf9vta89Kbx0mh
BIwnatA1sAUjEdTETHdeQqcnZ+eJG99/R15zPfg7+5XfXfnbe2OpWYU2Hd6fVQ05
LAQ/SFlfzWKw9m6LgexnMEpvZcgsayFXuDXmBm0tJlpaRUENiWTuMwE6Ul6kqVpe
8mre7rqkxDqShBiaMvH2QfvKjdCO8Z/oYQf+TIuSrzKNNCO1m1nWmkCFWxLxvICj
kIuI+KiBXGcIhUxL+b1DbEq+DRbmOCE4ycobVxvw2w3yZbOEAnofT6M2qvpftdoi
tbEO+wmce7uT+xL3vjYmN4XoGFhSIG5VCKVQKY1NPc6aTfgao1sj6X52a8cZ70eC
k+vfLVU7i2oFcPFMGNgrCEcTI8kOxyNbzm2XyIoYYdZz0fpHgVIg4xeqmyzDP78d
V3qGM6b6eg35l4iAsofbMApGdWDxj+O21vWdM4/O9pcgJFqFUJLG9jPQjyH1pBGe
wZiRKa3Lt45D4N/trdxLgvH0Qk04vqIwcvA6FgtooPcdT/RIXnYkr3FkLW51Sbn3
AamvuhcWxO84yQOdGddbGBdqFjKn95N3nrWcEV+1kHYzV/0ON+KWpve2j8z26HnV
CWuYRTRVJPVpVw8JtrZZobffUB1uaZS6t7Csc8lM4uX0WHH39ytvPztK1aUwRq5j
tSpPTUh6enbQo+2GwsOf+8K4fhAeIBQ9d2JU5B6jgQkUKM0U1BIs5cFScLc2TUdL
jHkUj481BjD2KxnZmhPAEoGYODeueN/z8/0dcu0Z/kmCc/mgCUuWo10EnVkAIZt/
xt3MK8MAL/3+8Tl7KFTVlKY+T+FHWxtJgQvHYxIjwX31YeR0LNMzmOge++8drlIt
cIFa9F4qU+XMd9oi59DLkjN7O3qvGPVjsYX3fH3MvWnCV68TE8PCWmNauPtjkKPZ
xxcDCL0TSrLJh2CMBenaqa+D5Rt8y9fvTk82pft6ufyCVz3e1js174bk5ijW0BnK
yeeCOleaVUY1fdrhUZVWpD6KsVvfwYWjDngNjBYWBwlaCLDbCsk1/NCglGpIUJRm
6jPFJ0P4/I0re5on59yeks30HM7ZDlFduADwd05JyTEOBuLSulOYqvND35Q3peud
EtzsyVh1QCv74ujFqcKYINiaSLvBoFhnhrm0XdroXFqG1K4iegV8rm9u+YMJUxo2
GJo3vNbGGHRFXrTeeiy7J7JGaKRDpksOxln2zkVM7nwnPIsSSLCh2pTAfdsu8887
2QdDgp1AkMIKtjUj7MSkTpMbwiIKqtlphCIzdfVSIqj7vRzgv1fMuJF3pTnM88yr
UnxQm5aLQE5Hw1ffKLj6Bn3hF5QOyIx9NraDv9plJ8PspmDxnvl+DACSEZJko0OF
Bf2R+WCGcwoXGsCiVDp4nmBEh3n14P5r9XHL6WFnVOMJ00ycYWWWUtOZjCoPiqDc
89G6M5PwXgbOxK0Ri7EM5kaqGMlBcSQtnIAINgCVMeF8xqW6n5iGU+bzByHymzHx
zKrWXrkofz0p86yrdfyL+dVZlcJ1RHoIhbSCoR50OCGd9PEMY/+Mu/MHiUqD129/
t1GT4IS6a9py7uShCs+WlNAsMuoSDEInksUj9KtUVBmewJiaT7BdHlbppSuSF+sP
38uDc7YtXceOjfLU5Bju2Vrt7Z3de94/eclI9nPnraAQiwjtyJgwqzcxhAb33Gfa
izAFQ2XzEOhLMfX6/7DyZkQV0Ev/XspS8hZjIzOwtukn/+0KYcmac+omnazsDMiM
3L+ueJRFshWy+HnIHZ6EyNLO+AbhcSnVNLWkTlc3FAYQMGoEaTlPnUimIrIWgkKn
dPsKULFMNxfBqZuf/0z5WcO2QjDduW7EGVQrlSB9x3YMOWwrgjQoAl1RQiFYk8kV
rfM9P76KRbofgdg448jBFcSOcDKgk5Im4cG+TEtS91TpWDal5/N9HpDvmUe/okvv
R1G1t+MmgnaX9SxsWHkX1ESSpfIMzBvD3Fw2ZhDiPgoDrayHqIMBhFNYsXgfsaDL
iiRNrdLrbpeIwilaVc72nzwCcW8qCVggyRysb5BgQky2/k4H/Cki62JkEY6UHvhL
XRHvQwjA/wFYOqazYsVr0YXQatwkYfnCTaVw/WERZM+qCz+4retVyMy0QDhF5MtN
Lns/T4l+/0EhTBQ0sEzFpodZ7ia1/L5CTx7r3vwwLuEqwntAU98a3KLbR87fpcMw
y0yAGRgPERjrIBundZ65kLcnI9btADIeKASixv1x/2x8SYU3Xd3VXLGeSR+QQiz4
2EwkRhiFoOpCCIzOZr0ETha/x9Ssd619WEG74+v5JMkg3JBUq9fDZzstrxSYvMxd
S2O7o3p5WxNIb01uXNJKbb5jyQnzPo6l3X7mVaB/KpcjY74hX7ab7NdcHrH+FCXW
yY/tKQhc7QZovFXwgDnrgwLAXQVA8y/obMMknn3Ky/RBvvkHKzdYvANJd7XfpR+j
b+mO24LXaLvz5JVg1HQu0/AqWuUNntDJb5s7JlXQ62wppRAOUpV2uP7Rq23ZQgXf
mPaACpSWG+EiZhlFU4L/KRyAiJ3PGa2ulrf7kT3sFuELSUEPVqlDJ1o8skRJRf2B
48QdswDZwkziB5WjevpQz2l5QRpgjToTMXV9+ow6QUC8t90NVBs3OnV3Gu7/3GCq
FQpnVHR6h/raQdgxT14Ne3BafSX134hu63IqnUko5EKeNvOoY+DxFjnMnk12yjGF
/hPcyrhM84cCbS9xZARGXWtjfp6EAEWgbF20Mnk4pfv66fBjXefr0KxnJJ5PzMo+
Zv4iMKhRqrByMO4ZpiIUriGZhAV90hoEp0lcyXum7VGm59fQ04D5WIrINM6/DkvQ
7LKcX4uVSYmnVsrvHIAGVXNYsQ0mnAPbo7VzWeMk5pfxppa3xnsf740zts7YqV7w
xZoFYQsrwOdSux7vMhl96fgnB9YcvvdlcPjZ0Lnyg1TqsxZtH5gTjja5xoMM1WyZ
M9vot8ONsJZZvLg0Yu4H7I7RXILKWJ1T9s8IsrnFhrZe4fQbC4pLefAq4lBwWpkM
E12sxDfdb9SrhVojxUucoIheU6BODFn8uTYALARzEvMzc6kg4PZ0zYR6UnWJT0/Z
bBIS0a3t0SVXeMqJem8hrD98+/u2zKZW66jpaa6C1umGdWh8NV0NWBir6IaePsHS
egRPtR+QxKdjjvZ5AR90pb6ae+0Ehdsngerhy3rwGS4ODNCH2R9Rre8Rh3VXV+lQ
S1e/z96x9QCtlWXL2tOASROGhw8Br4jVf4TUvwsqQtUEe/ngVJfmf5NVMEC6+z8I
tvR6O5OqQ+pUJop/BF8h5w6J9HsnQxnI5yMF6DgcVhd4w8Zj4CEXawLajZlBZOFr
VsHYj2eo/hYv67hk7OZenO5ygUvla0zuIO6puJVWCHMN2kui8dGg07AvbNTZs5r7
hpW+Bt/GRX9aL9Vv3MdJxor+P2ZupluvMJSoLHfDiKc3zQKrf6kssev08s/vnnyH
sphDpuxcTBV5HlR5lQNOOoS49PU0ki8tL8H77PE2LHnn+n5EEubB4xsmCebC2XMp
CoA6f8eL6EOdtdCKX812r1OL7kfyBIt8Dv9506/bqSwNDxVfjDtywDTMRx+MzuLZ
NYxYekqKzHMkEsZSqw0U0sB9+9/YSvj0qp77rFCX+s9xbi95C4yFd1OUpnM3a6Ep
vl67Z2gxLPryGcO9xHsLNVavfkohgu/OMarp95vCmkWMVBxzFesCSJBXtItryunG
YxtzcWS6PIItREBp4o+H+x1L2Vm9pTge4KfqaqsBpzkRGWZawSBLLv+7UBCo5wkM
3dbybuWh9hGspRNOXOch2S6zHj0zXWkhYHk7IVpxUUmlFlI5XqpxBB9R0x8Lfa8q
29Ih+gVRtBhWGf/xNVEmBet4QnalFwa5EE+heAW/mDYEFmrgQRYA/+VfkPF6vWUh
gjvB7Wj6SG09IrWzGMR66zn65BewEJXSXZ7fmZUNJ3J16ay2iuXKI9BbGJM81xCJ
v6SobYzBWIrq1HaadHGl+bzSJ/Xkqp0pEXJv2po08rvu2PTumVL5a3+HSWi1oBrB
MhHxJAPC00mwki601NZkamzqOkvv99w5GX/+Vuk6VMs2PwN28NKQkbp7lUPxhASH
5kE9jHfT9G8/d9e5iEOVpeX9rqpUG/ElzH+UNyyVgyKn0tf1T4w9/mtabKymHE1o
TnTblc37YM8Ekvo4jwiPg7DCGWJcAamTicD3J9mM+oUBCRQvSIBE2sjom/vG71xO
qoNoIGOY+vt3Nvr/vOoVY11FQYaCGIaty7aMta0W34pj3hyThh+TU/P8t0l02+6X
foEmUpBeDUXackpLGrHVuqyx1hy8pESI6aZELgI26EQ1plsep3Xycp2LlnymWswI
tlG0thJyiIkvmRmqrvilgxGlZkoiAtMZjWKiI06nj4A6j29UyCqV4aZwi/NhuOkU
ofa2ocSPj6QBCWqY6WnOqX9URHRoydLYrDVZGOBpghomJJEHbDSQ2CNuFawoBjnk
dN7BdaVYBa6214hduOwz7JtMUAaYlgxZwwhhkx8T+vLTW86vU5VoRNtnpy/c0BlU
R5sS7TdGicS+Bnib/HWpboCr9axEVGM9JYewHbjhwb/NSUyttn+L0bXGSevGgG2D
fXISr0I9Y4vcp8AajF5l2iYSYfCTMfPiCHwdNe5fDIj7wVIF5J/Dyg62EQ2I+Uat
QoX/hy6DIEuwcoe33DWuvc7qDrf6ELk7Ppaj14C6zj2zAcYJLo2erCWdfkfz3Qvq
5T/UnS7wGRZJg1mAcXgSzdljpr67vzc2uiiMVM/+O5RZpn9neLVtjVNu/fr7f5Xj
8vuHyMfUO00U3iXs28u0a3doWQIq62DqFBauRqGP7V1RG7kJT3Z1T/ZDwqLM1+Rc
u7mPx7nSk7C5+qz1B2VzVfgGH6xQPSKQ1LatELlouWnfsfQn6Jh6Ofx3oB5WnoEA
w8RuCSABM2WvUjuGYGKLIPXLZsp1LGbO8t8uzrHeeAgVuEwRXA7tFsnZSTzNnow9
gSwMgyem0g8cDCMZK/1h49v9YsPfN26lbbmFV+ilfuDfHO1gLRa+B39Y7Ces4IRx
itkp7xgkEwh5hqcv+39tnNrrAU7Kq8/W7KETwq3Cek0WD7VNUovrIgvNrKU1oe5Y
deZeKi6wJWv0ok/PVjGZGD8XL6iPrdFNxh9YoUKgJYf8yyMu7WeGhrh3FSWKsJav
MAwRO2r5ajC+Fi4wqWvqTyxJvaqwDH4PNZ4G/9zs3mmEn1OXQvdD8FhD1CMzPw0/
sMCmpxBYDxAwUa3oeqURZ+CQxCQCkAKz9cASmS0d5kSzIo5fwuDRpxprMnr8Hlsz
JQQNskDXBfXX8kbfDMYdZwx4m1ZISutU7gJ1DMl3g5jAFn+QUP+M4wV3YNLUCLvQ
ABNg+MRwjgI61/YEK7ay5fo5TfVkDd3gfzDDGpr8aSL241TQOJd6r1yW3Mpmkkue
m5Ngt+Vv2kqOaRq9kyxixkgFwREfx1Lx9u2Mq0GPbz8HfuU7Aymfc9CiHPI+PHh9
IA7kY7uEkTLGH64qLbNIksJecGpRxzZ/Y7++KVXOOjSFfVEcl08Q589DwkPJ/hjV
AwmzdfiPafTyEKAQSZWbtXMN4yOloNvXDyEZSTzYzRVe518XD470JBM5NfG1qLBW
guAAOiP+KRrr8IPjoxh+0Chs4njqUjFm7wSldESs9SlGtzJ62U8mgfBP+XQk9ZGT
bpXpDdhUntIdB5AqiPgjI6VVqyzM3KsgGz2trYKExW4tvryS9psWQJ2x2NCov8Kp
lI8oyaX+t/sM9WTIY9IBoDX3U61W9angVS9X8ciNxD0JZjpjegpf/RzRrrR/cNX4
hmLYD+1NcFgoj3FovNHn7pEhspp7dSO14orhOcg8ON97Yq9i+QzodcBsotKlnicw
dJ2XsvpOY5r3g49GfompYEdyBs94oxlVZSe2EyZByzn5IVhzkhwwsjYOqE1DyX54
rt71uWN+Rn3bwVmvtlwyisoxcqmctPcmcaYnAhDwIDab7/xvqZz+wFNkzC3hPqi7
LYbhpSB1TEE0a4PmHDnQlpSNnQYhtcFPoLyCF9ihZZQT8gUa5DoCsi7EurMIzF97
YDrFbSBAy12k8dWyxHD9e1vrhx/35MN6lj4YgNt74xnw/G84ZPKHPBBUtypuCre/
Au5GqqUAa97Xbl8Xisbi0/mtKZXKMUCeL7QauFHpLzC/q26LIuYvTRmlHMnhA/Fe
uHzuR4aRhZadb+/ne14N5Mc0HUtELUoFUG6D4RQvAHAcqM0fQmWJPYWzcu0tHQru
4XMZFmYwm9zOB2Kzxa5pIA12sGsUx5VqEnd8gV/k9aug6FZQ1KShGAgkGbXiV2Wn
yYJ+dTI3tO6Xo1bKE+zKR5arxo4DtVuSFHQYzm2G0nTPho0gqtazzgRf6geSgBkK
Vh7C4CGMFN5QPv1plHP41quAQyqnv78EhfnQXrcgMV8lfOxWC0oB5FbTSnm5+2RC
EHX8sYVsiQ0gl59IXwHy6kzGH14B75K++kRGEmsWo+FTTYbwYeuqFuocygxIKRDf
9cKL1AMKj9Qovm+K4AX74NZlLjiHQucZbQsJ6aDR8Z3Q7rTAhR3JRgr7qmlz9+Db
nWCNnahh7zoOhcYjwME2pTt0EEykexHu1v+5mk44MaIrmjEol1Al9ptJVxjz0N5R
iIU6YuF0Oeio3RmrZEhtwBy6YafTCXKgfoNUMMcWu0l3IH3EMPGI2pB9r8puR/K4
kQTgShp0/TiyBpxBEgGR9VDt0yGkYiRynpd4yoKlTSG8DGUloMvx8Fn5SxqktuD8
zBa1n2nFI+NWbMkPkTfei/6nTECS9WmVfWowSlmYaYaJzfVxQybSQLyzNbXqDZ3g
1iUpdM2MIyABOGmfiV/6pNVou24q0NkLktJUvHJQ0e+wfOpQMM/HMAcjg44nAOq3
EgsKLrDJBuGjzNhPKKMnf0vmXK6YBQWIg35Z5WgdQoQuRMR3O5jDdtrCkxTWrbpF
NGcIq3xUyl5elZV/BWp5rYBEKU21C/XkZJwcaMNXi6ien1RKt3Ftkk2PNj+drU/Y
DZ6lxV+n9XZ2/d0fQpbx5JAszGoeRFlKAegD6bECj3llmFLoGTh9llHPEiUKsWAe
GyVLl8NCNPWB8LGRfjA5SJJ1EfSm5pEyJDdM+9O8jaS4aD2xBGmRMoU3hYkZSIs1
Ystvs2Or22xYFoJqGQ0CcprDrfucAB+Bt7Dm3TRJ6FCiwKYh2KbL6BqeAP3Zr0/G
IN305Agqw+J+2cNYn/9esEoLcS3WvEP9c0aqvimMKQ+TRe1SFN5WUZ48pf2/ISjQ
3Q+oUFqHLlC62gi0OSH7pLKfeBxqt/89Y66LPxpwlw7t0YVANKCalPKQCAG39g+k
PF4N2KA5kVvLosKpdo0r8FU3TXZpWbFYRS7Tc9v/4gMIbpDAekMuLToTsF+uJzP5
wjv/RPO+iHW6DOtu8fdhbjeOiThSJNJw/bcLikEN71hK057JaYEp5iz2LVDGBnb9
+opJ10RarEez5qGJKVHSzgIcb6f4bndbwC2RM3x6mBYmG/81eXiOZrd7sF2jJIfd
CRwWC54Vzyt0feIM6sVu/JWdeeyXOPGO5p8Bdo31fiV9AO5oEwfFJLkvR1xYBHtF
zREbfxZrdlv8jEZ6Ghkk50VEXfZM5jY4ku8VqHVyuimV0LNsusNnnmzFMXcAkHHl
FU194fShzM7zlucpSABtNIq180V2YnoRf8jK3j2KFpdjyUc3FCDwd+B1HLGx5VMm
CeULIpadfvvUTKBVHcPy4a+LPUQ4n/6+xBdiEyDInxDJX4IbtapSPmDVjcXSNgVQ
6f/hF7LC6B4sJNW4lCE81K+SZsyRRcshpndV7uVt2rZUouiqzgdQCCd2M0nS0C3S
F1GZqP9nyrMHzeKBeutFYLgnogIrwfel34XIk6/+5k38T7drgQavorgI4Cx/LSMA
iFFXFlnlmTCS0LHdAAYzde+LhJeNeS/h4AVTibjJkg19Dc8d0RzUbZ26IDUQrrar
L+nF66JTxit5Zj3C6iiTkiJD89HNsgruJo/nat4LaBgWb5u6sgUrtYyHvoOWV4sq
b7eZEhKNLI//ZrOKxYZe1Ot69Q2TdQso48vSQv6KvJ2ktRlYUQ10AHFo2AaFZaee
XEwaFs5lp1sKFPBq+fCPz0Xotp4C0svh9TeerZ+YEmGrlHsWnvowVHdXi/qrvYef
D9b0CaTNvyEqLSn2k489d6DcXwx40p4idsr6BROpNJawAvwhIvzNlqZ49TSUHExP
ImUcSJD92RqPsDHGIjfx2X3k1mC26mlsX+vpGqmEg2fZ1oNM0hsbGjPBNF4bMV2c
bELewByXLluzulJwtkK5O9gWgaErx3eiY+mgI31K3JQA5+ih8Kgo36TUdbPSl58O
bhAV7Yxx339lTaBHD/1ReItRZqvMobUmHH0PycsQMDILhZz6cBQD5qwRp0BofWep
wmepOdBz40f+JKW2huWjytaWgsmBjINKze9T9HoyIWoijBwxxkK8FFRMhdlhArKT
g9xuYYraAWAsx3AgLXm+V+z+7+qSAutc08fhwE+7iBhgz49SyU1FQIy9tCvkOwDb
t12aSds7jwQDIBtCUReKC2d7T5ggTCTyx+FndMpMc+oE1o6o5AuKrHznV3ibVujh
KyL/swE2+B91dj2sX31vFTv75Hom7akZt0kl7pzGkwYR8H5pyBWdosYTL+EHoNAr
9R4czS7c/cUc1KdJNAniZiLS5vzaNQfJ5Ie/zTGandiD09aS4f54vOwsAjwls4Yq
ZtcDPa28C2Tbag9Bm1J/xzqK8uHkGsyDIO47UsAfJM39seFveyaYPWMxxvT4vsvc
/9ELeQgNwshOajZtavMWUir4r0Q+3oeYoymcVzR9rHLKb7wjCPI6FWFZu27cXiLq
KSkfK+yv9G0Hjbc8cYmzu7uoscJdGsilspKbN6CVQ03/E/QTQL0FkW8rXsZi/w+H
x627Jie/jM0E1o68uxP+B3E2KaRQmyAkj/uMPK9ZmjbOz+taQtcL17+0mRL6nUm0
zxa5nQonLnl42c298mLbnZIhGiRUJvfL0tYohkJtbsUjTpimH97GVMAvdPU8niuv
7HdoTcbGwwHKm92Fb/TaJaYur/MJRW/Uedonp8xDN8k4ErNrR+hnUoTdE5rITpvi
AZEqNXqmW+VKHV8wfVROVCQcuouoX0QB6Af7uyee1B6sAphga60FuOFpq+UcTGQE
79Nv7HrTM49jVgpwde3X6m2MtAPKCI7H8kAByX7Lppcr+3SvsnEoTkiw9FDxXr7U
cRAL9esmU1xqWtVnOUymuX5TYnMWB1syhndm7aaKRiW70RazOMAkgukvAWO+tedL
674GSwEMF+YsKEoW3y5tI/6em4LQx+RqlR03TQzjLOOObZ6LSUkvCWp06S7U5Il6
91OMJjxVX5+GO0+QZ6Q5dhMatyKmIRrnu+UizMtiTOg6+XicZ2slhBdWfPmbIhgP
M/IxsevMSbLyN9JgSAafj/ZM3yV63+BTFcaPJ816WYywhTuBBsRk3y29+d/ipSUS
rNk6A7zvZ877UImBMuFLxCF45eDPs9jt7WTxm/C8Cm1mxUA+Q1a+eQ5WiYn3nWjr
vF6Se3a5b/vf4da8u8RRy2WvXNBGSrNrg+Q9kyk9c3oPBQte2YZkQPznSeyayhnF
lSQ+0jIbospIrzOl9CxTZOSmOztH4pX9vfPDhg+Th8lAyhJ+iciV8urqqL+tBMYm
ctaqq15I7sj8qnOAPX0xlLgEEpibU3yLnAJmpd/0to4HTw/FeMRPQj9N8Sberk26
62iKjGUlztHZwe7ojYv7Wm1Lv2CJNuFhFuL6xiBKuN8s/LF/WyvMhlCsjgHM2fbn
55LARCb9WpZTW0qAZ4gOkAOB+xQz6vZicmpYWrrohVb5hTTd9EO/oMWBMGloIJPI
xOFdkYtDX7pBRW+vNhkmQtxLfnXvbBVLA/RbKKwhVbFNAQzK/Iy/Ph3orPhSOXoO
nuys5XCd/HGEWiRYmxC9he0IKjzNbhX+MWNhccJbUgyHPZXgoL/f48vyZwUK+NdF
077tX0+8hSeFD9XI2+tMIYiCItTabag2mNCww1kx+PGT1nWfuxGclu+DUYJk9j52
NGTU1UXNntzvq2I2jBEzRBFWhZopet7b3l6Fbtd7oAXfwgrJynOvo3Q2U0VWTOKp
bAe0UGlNzdcpPCkJPNEqofGbdKG01qvUjL0SxtIFBFalJllV8L4fok8p7+dWQJ4H
DCPei6Zc+MzUrXg2/0DZTes2Lj8NOPU4NCDlKqR3eEz10p2y35Xo8DbMatBpTqTo
jt606YMgZAVb+CYwSfU3nh7WZg7u/Fd5go3hcdhLtVC0lOcQrpDnVePtcPW9fRsj
145a4Et0yGgZ2dyyKR8m9tJ8Nb8XfPiM7bv/OyxMCUP3rxg6LH7HXe0mwdFdUL2X
ZnRKvrXvAl9Sqe2J9hrGyH7X6S8wjL9jiuhKEdXDtDbzm9g74ZaZc6Gfdm4XRAWR
D4YCWhGQE3rAFCDkYET7b4X5JA3lcD84jE7NVAdt6WeRRGWR9yWPxWkpTZDWDNGc
VVZSji7LB4/7+p6Glk09PNMSmofn645LNm2D0laCsFAHCyq4YeyvUv3FUS+dysfm
72Ve10y1AJ1sWMWDiLobM2oBSHaUYdideGm3uVxGY8K6LE/8MgXe9jxRSGr6K6fO
M+8Kl9aezvjrM1uGIS+HdOcJdR+MVht9Ai7mrniXbyvF1albd60cG4IWRI4qhQkg
mU1DSk1z+Y286LiHSFWzuExkRvVEHii89HqBbr9qwXKI+3UqJTtKQtJV9B39hFSg
2AoPBvTfI54ypVkR0SDr300yGou/WihNOZhWI8uzcDEWQIl917LOaTEZixP+AzuK
MwkCERukVM6IHRLwm/IAhCzwbzb9xX213wDg9i5AjMcUFaWSbSxPg2AobLZoBhxT
bJjt6Kyt36Vd0x0cvzUx5Qw3mVE6yn3IzSL5eg7uEU6XuhAq5RsE2OCTVtpQvGIk
Jb1zSQcXMDOh98yeRstbwBmOAYUhVbprjy/t4t5HawEeErraiUIvf5rKMR4bJXAm
rygQ2E6C4PUPgS9gokbO/LF4w4IoFQpl3ccFM0wLWMydHK7dtQxzYmxlQ/JEjeuC
gt1ku5bGxg3P61jbGa+7tHa2rqvZYIIGi1awBd8RSqvLQZzE7BFsOK6IQOVq6ror
qVMRORN0Ls7wej1UTJUZL7vDISYLMrvYnDf/2uaBpnXEily7WT3o5tA29meDncNB
PsCvAUrR1/kWapQnuie5DpnV3ydR3xbar2lmF6f17bdsXrEs/KQThpIiQ09bLvZa
raQLnNkkke6iiWCZVQ5qRhR+VasAgDCYstlIGl4MGk8V2rZMLc5UPZG8mveMg2lD
w+/nxtvPwKKI7I49msWnUpxifO22XZ9s4pv8HY4gVSPaSjmqaiO13JhVOC8zgYxa
pl2tkpPcRx4bLFDk4sfV1vlEKzuC5NcRiH0zbMX2b2WOlo/eaUDHcvY1ZG4LMrfk
symtjGWxnjjMXVSir0NrcuqeMSqtTIGTvZ36Mn625CFjGppwF159Z97mJlNwCzIr
3y4t8d+ZQRLk2MZSkNmRI4XA2GhcWOJdlj1U8DWyKUCJygBm6L3zXDD8UwKd+hoo
RZYXFpMGk4yMSc/wf5MkZCDGBmB79vgAVY06r8OkIliDUIXlTcd3lr5g9x4HZzEp
w+fcJyLdH/FQON4Q3z5aXkl8teJ7BjoZfZcIWdiS8vTfjk2Ala5ZZnJnUjsZajkK
MRWZGbH1XKWRVF0bAOctRknfLXj5g0/1kskKAiQJFl/7r8IUvaoZP9ydxCnh9xN6
NiCnqWv93LrAV9w3f4OUbPnj5xeAhyJfW4f1cdM7R6X3nLwrI4Fttoi1JSoPgFNx
n/0yzqzQY85yH6F3g0JAXiEfe1dgETE76AyD89jX3VMVK3aTbItUhT5xrdxw1AXI
q7BAvzHUNsDJM9lPOoCacQS3dig/6hWJIOYk6YYaIkCJx0hLzejwCFlfhenpIyQC
dmW/9fIy35jiD6hdIQ3SjvqdpFK34exKqPDs0V4gCoAGuYcOesfGiA9XPSh/P44W
/V/Ec6et5wEtWYCETq1URlFvTfryUz9GOqE8EdSZL2CQYxeHJrffq+GaJ1Wc+SWL
x3J7b6azGem64KtJ7LzDd6hmMRy9o4+iZbqDUP9VGc+ek/xevyvl0WjVNI8Odyhl
ejG41VpzTaCgHqCj2BhEKUya9RbWpg7rXu/Ae2mbV2EPxcLQyMg873mzQ3cvs0bi
bcTJrLe9Ki6kJGD7ANriEc7j+Q5QOHanwzrA160gV/KNvyTKAPemkx0HU62zh/vk
cosW3iXj4o268d1I3YrmRL3KWGeh3A+UfZYLIYBmw9uo7xkmgDi1UfdeHwdl84YL
qOeFtgRLbfWdFYMPHW+KWWeImKtXhosGIPIcwoZxC7NMa0x+aEs4ABZdBfN6LDJo
0FRsLsqAlb3HqlX/dCduQ8wVKQj+d2mYJpsHeo44zCjhs1Oc+zgQUNvyalXru2LK
tfJF0CvUvrjsW7vv58EGswgo6HeycFsJPQ5Iwc0afPOVLsO7hGgTeM8hImk2xCNh
bx2su0IPaawI3QFg5KQ4spNsBONRNks/vrV+ZaE2TBT9q3YqCejoP0Eioh9qwKuN
cIN7h63gI9mu6aV51owT6HkcmLH6ZmdRh9o4E1OYEulHtwMzWyoaXtkAGBaYQi/S
+uZ52tkZDQ97jqkm3wRCJICTIRokI/GfARUKLOD2hz5/H3CWUEV/VjTh3ta9ZEnS
EsqqMeczW9i8OihPSFpNjcbvQ5oQUgk7IAvWaVzGDINHaua5yey0llHw2Fh5Hu5C
wEyB73x+dKM+gPv8+ooEpyJSPPs+lzpxczMG/qgXG74RcpWzo45SDr9Bb+ypqwbB
Re4V7SWNxOAb8+4FSpXQDQVFtoawL5u1MRcp1wj27iopaGHkPwpIZGV88Syf/c4q
9mxeD5pVK18RNz/05JafU/qixWXvKY6BAkafm25Y9dxYJzJTpYjupCS0gFpc4gJN
hvW26TAq9TWmDhg0aH0572SAuBBzbS6YJYUjCOxmB2sK+0YFT3kgwDSc6KIo/DbJ
sT+Krub/tzM+XiTTwTOOlXE/fbkaSI042o5FzmSM/ZZ9lrLdvNbbNMW8CQsjURHg
cXkqdyjGYI6xP1MXW9UxxGY3vG3mQRkV5yMfTBw3xeWrDsP4LOdLvAlIwPu8oSNl
BK4a4ilY2DYmGQpgCuoliCS0eg8Lrc1dA+DUlWULMYjhj4R7BdvCaLpw85+5y8ni
K9TapV0eNAEK3za/bWJZzmwvctyybVHJzi2GHQ4IOHHzKxuVW2wC30VkRmlduHiy
Zd8P9ldYVDd0kAP3d0H7+Onjc5b+2Wr2QhXBn8nWSLeIQuAkebcNVDt64S5p7V9N
NWOFNPtvAuxR+AwppwYsMQAjaMq6btjiFj2E5pQZupRvumRoHIkgvLEGMRlToYTO
6II+3r7mD4Yv8ZCwD7EHNCvova1YtDezQDPb9lh3ZvovVr54nBUGhd90tbXw0/mb
sldfSoltTQAdGpnr10O0cVvQ4YJ8qWFXY2zHy23NMlaw7DwOsFil4NM+vxfXxqwp
pTRDVITdqgxVkQklI/530laKJkRKr3CWpgBqhquZPrcF9KmRfr+2OaUD7Lvv3K2p
YoDz7VTu2gvxhrYixIWh01TR8JL9+v7Jg7lOnWu0jLRF4A8t4N7KD2BgO7xnORdK
FMuQp1uTMOiGtdayAtQIhsiv8tI9aag3pLphDa2QccI1P3fWA/mmjrbRLUazzuC3
28FEOTNyKEAGvHDGGUT5tiQKt0GBkCqtjAyOqBSrk01UJK2Phug+S31sf6LND/PE
CAzLSmX5TROwGi4alP8ZKvsI5zZVa5fZPeZ+QenV4vM2x5SmrXveMJVzhMIcSuVw
vJKB6hKExrnMYnhLf2hSlZ+S7X3vOVpisc7XMIf6qz/KbDHgIm8kKnbKHlcdUMdH
Ow9+Lwj7lAvtmUQM1w7oyCOhClMKBVs8bpHuKZBIaqbZNlsBd/8hOA3hU6ayosfl
IKEEl+6bYKsCXgNdn9JhptFEX6q3q4OwekXiC5Ks5xZUaiI4gESwtJRTm3S8fWOg
Cnb2IJ7hil85Lh6TffRaO8YoJvNPo4O6SE3LtzSZYeU8veBPS37MI9iVZdNmuYBg
Zn4Nro3N2iMAXN54NEr7rCyjCMujKmHX/stiAve/P+AM4c6daCLtjdnUHBLCa2Dj
FRvthcAhsJylP96onc1W6jVssk3woBW6g8PKfYTHJ65tsSXc3yaZQo8FmVZjtcte
HsYx3hPWlvhQAnorKRqjmiSI4VMQu34dV4ohqxRY/q0l/ArtL62m0719sXQ9M0N7
z4PqzvmGFzmMwIu548Z3IiLXBZ36mD8W44fSf6qRUmHI4xrYVGQ4+aI91F5tOBzt
4gq9rAQJV47moa1R7DRBOyVig3tUDLgZtTxHKvziAVCUznrpOmhfrFKzv1uLSrwZ
PnIH25p43Hiw51c7gduJKNyhQxzT+lnh+bU95Cn69e4UfSBkMVPlPd7FN5BXmjM9
8x+579tUEokWNlj5cNDn1+JGMk2BX+1fSkjNVXL87M1t8X01P30V3cQ5LYyVNkfQ
b+RM4Y0DJn/2R4xrcpAXh/radmfLhy5mQyLCn2csQ4oM0CA1m5+2oeSLilcMOSr1
araIkAopsWTbI7V64qUD4ga1UPilcJLm9s24UmXsD4cYgULRjxbn4eWgvVKMeDCm
DUd1Ean8gIeZiXm97FMLJaZneBF9muxWmndwCVAyhayA5Pl1RKevUW8meP8Fg0Im
TS5oYicArsjeuMwZyIrrQqFLGPd9zH2B9eurvIc2XbtM4DZR6nq9O23x29aPKTm7
OypbQWZ8pFbec8PNMyEXLfQ3WsXpC23VYnl2BCv1apxUw/0e2vvOvnrNZEWQ7JYe
Ji4Wxtt2golLGBLXjBz8rq77Ozb3ayWWIyLhG4VRp/zG4Pnidp9HiLQH3EiIFUIa
IIng7nQ5XnrwKR+d5x69FLrYhYOhLMjCdcwUYcOJQbe5qBhVYJdAledKxpQdUgSm
xVhMtuIyM4uQ3glAB/BpiSJgr/kmgbZC4SBWpycpHN7PVhLUuFj9KsRcbdwrbPzw
5IbCclj9b5Tdmv7HfbH6RltiBX0GVF+2vZtDt/YXaVcBAOtB7kxBJd2jlVM/UYFS
+btAlgbMY7/W3+R+DtPfB3eS+1smlrjhV7zJn3Lp/S9/I9HGWveXTPYYzVLq47To
qk0H5VMMCuswZjjkdYcfARZ1HoUtZtksvqVBlA7AN8plq9iyXragWEfY2RcCCP6H
daQdG79r5eTuOCJZ5Eb6GW+iuEnByRSKiODvMi1NRAKFGLCw3g+WulULVNeCCLh7
XYVNcTsPh/y3cTVVZmfgv7Mmd0GnHkFYbV+Neg2vQXkjWKkWAfj7+s8rgp+xRNIx
jsVM1Ju4MpKV6nRDJudYux3N62WZQAQiNmDWNwm/N24JK+9Bg/wVoDXh6ci3G1Mb
yIsyHoKEbvrXlBW5nAr0H0l/15TzVX1aHN39GseF+4PcefwEJjq0HnXEigb/iML9
rCYJNCI1wPjrgr/5E/TNqb7YfzMKZqdoz6lDcbNTrTJLgNgMVvr0nCNZ9Yrxr8dg
3NwwtyEVXFcwAIkqWhRT1oi83fCZW0yp/7n3kBojtKx1UVfXv2qHxr5yhcfhQeFr
GuuPR5vcsIFPSftxLawttoYwXJqEHIsclGWvCmEcFHVLCNoB2nQBRztTG8fjgzsG
ugAv0AZeViLXfgt0eQDk3jp7TuBorQHDLCkcCTMpwAZ17If3RqZTcpKie/FPQAJ3
jqQ7ZdiP/YI8q8ovgBl/rlmVAC/I8/yWbtOdPIZKDenYRVSTLIP79lX6+FB+aKhe
PFnQknBhV4AF6zXGln+JUZo8aI+JqhsLkQUU6Tm9j1W7dgUWDFZ55lE1M9rENQ1W
Ek5Va0WofQFohBMJpZc6SEpEc07mtzOiLlgz04w9tdzXyVUJWl2PZ3uoiTxc1znF
jiUdg2JATx1EihUX5t+JlYlGJmI8tQIWIR4O5bZIyCT5XHS2rJJyyBuVkzLu6HGG
JMqVRi/OEBsVSPfz3P8yN+2fq9LA1wm5HjaDQg9/EFMEBMGfOosFOWwjUUwpRXKV
QpgaP2TobU9OqsSdw3JjwevPKj0ENYJQCAmyVoOQcIpfhrwYOd3gU0PVE38HS955
mXZXgJqtOL1kjEm4kMy6Q4GL0z+7nV5GiHqWTYQmw8M1nJ9aryE1pUGzrwGe2Fo1
x5Hj3KcKH03HCgrEzfsH4bEcszMfZ1m6nFz28n7z2Zxb4kayQOaBsYJf7N9/Ften
gvZf9gWMaNUC/nAMCOaXVcHZK5TbFprKhSDkSyp1nCKEBJhRHc/eiLC91to9gTVt
Btq8wrIQtLjrQTxorGrDgu8IkhqHatIn4UvJoD5dn+k2E0GZrZQkFVcBbvTTURE+
bpGzJNYLEVXi7ppGANuxFhAM/8SFSdTV0pe+8S1d9LYGUvv152HvqfM9W6Fcmcv4
falQzk3n/l4rkklt66TYSELfD6JPu6R+fwqMFxqKXXSJ1hoUxe91IhR3ANelBiAP
2amId5O24hdEpaj7977wZhX8Bepkstjy6fN7ZjpQ3Ocsmr4uyhDRTGK/8dO78Zt7
0wvEg3tE30Y3HIr6LLMv6YeVh+m01mHomQPuPjd5EnEAmnFvTriA8PwUl590y4nI
upjX3sZTmsBUU1vKGHguqswEuCx2CAWIfGtpcxG3EPdJEHBjYy5gpsNg00jlRb/E
8939O2hPeqwpQ5AHPA/qyKmFEaJfZtwXG0vfGMbiQXVqDZI19IoA35CiktrFfLmu
exNlNH5msY+oAdQFpXH1w5Z8XlJDvKXVgKAX55xq4fGQUtc0FltOWH2OWZKl8OCX
Nl32H2CpGiNTFJODSITigEZk323Ab4KQYeXs913FeaHDotbznm4vJtzh+V/0meMi
9FRqnTcTbM03S3Wp5Q1+6mJBMcrNYtrMFVJZALNhZRFpdhlXw+/pYyVUBtCrcZ7m
4W/uxp+8u88Oif5byDhf2+TAIF7cdbfFdlExysHPw0FZj0YLcvefh0XN3ZivCW5A
KeGTazF2fiPppMmnniEdL2Xbiz7qsOxhCkzOpqhUvmMMtix7d3leMcHLqz2NTGtm
pvQ++YtlLIlECRhWzfBHq2G3kCtJfzi5L/ROUBFwxV/7EiFMsdxbFWMO3i3IPSzE
cdMJDtPQV+Q3vhRhERKJIFi1sLa8mVSDCE4+RO9roq6lYVT0kHWSL4ududPgWVrm
X+7CRQz+wYoRZI/NQq937GpW2wqXqZ/DVfz5pCUbsswS7ZPO9g+khh/aUXRFRZz6
nmD84JqFyskW7DF1Uj6PvrBxeS9OndP+RtzgX+QeawaS3D4uhad/j+WIigiezY5j
n64hfwg7vOuWkeALYA/m1yuQxrXK8Z7SfHxoVFxkNZfvI4NhG0LahQV7W6cio9xW
Nyu18ET6f5RfAnNsLpsgn76K5KquBjwciYNMu/gJkkaP7AZK/PHb+j1kVu+4FaBd
Z6+JJQJFyMO0uQ7PL6vhxR+syU3qZkuHbioBNmi5Nft6McDDYOfbnUTeCWk+EFDS
wZ3n5WxMKmJX8hP+fBeKwjyDg3nr78JL+Mgxz/n26hHH0IDrcGDnXsNJT8ttn4ic
KeVUpgvUNNhlRqnlXxTmuHDc9FRdQx+F1Oq8gTDLUM3oGdGdvf08P5vKwB9sK5Tg
MjMUgCaAAElTpHTWcahd9mwQfHgoPOdV19Vs+Cgjl0JFehVmMO7XdMj/wmWx3y9r
lFIoB7bsan612BSX6peFZbtWNhBmwMLkvN4cTs2cm1cML+11eyhv05H+H/ZnQ3qW
RIa/jpiHx4g6znfOD4XUfz8F1tW09wv87Q47Mano0kFnvFK5V6RrK1+9UZ7kXbcD
vDM+x/n7yEGQLAHuv8WdWYP48jGAmrbE5ar65ZhK4f13EXavtf6GuL5Xes/xEChz
DHiMSiaSTR7bUC6mMZANmBGQBPQ/aafPSmGAw0FWkfG7DHA1BOeCTIhvhR56ENwt
ZxkLSraherbI4rVQ1xAMJrk5t5ReRF0it/EE/MSV1h4a+bDeNKDrnwXlDBGuby7B
hqZqM+ntzhESJ1IGa7+OZtywN24VnhQwanhaAJa6tqZbjVOmmkfKNhw2Wj9kq8xB
cjKoD9YfDgP8Swx/qmAx1yMBSnMvjZSrJXXBL1XEZiZs7SiPX5MGswc5TD7qYQgN
AcK5Xilw37wdqQxEYj6Qc/D6ar3uj4uPdynw/nC+Q799LKAl/XPMB+lEWFp3V4nA
EUQrtpTn9KjyXt4QE1jsG/1SEWRrXGi6pl143gIN3q7wX/Gw/3/UUhTtn3sZ994y
NM+Pcso52mA2tUwyuk5dfhfVS+5y/T/3t70IbQIAruf9tHx/wUQrfctnj0v2j3Hh
O63L3BAOg0u8Os81nC2twsSiHNvS73ozgnbfxBu5eimg74S5VH1vlo6/LabkKYHH
yLT0EhJHmj18xQYZ/nl1BzDLYhyg8L2nJ1BYtD78cAkmRO1Ul4glxiQuGJID/c/K
AtoNKfAXjaN9iO1X+KGp4bLjIiBN3X56T/23qnZoSGku2q+tIpEufVXlq/g/iccc
Wfy1KrpS5janaYQg1l8HIAJsX5XWSD9W8Ot4TBm/L2XEBssVbynjJe7+vpxA6IGK
/teZ61uh/y1uL2O+L79V+v0PGJAnbbYj8KgqGQRrwfSlWAirjDdDofT/pENFTBIg
aNf/2ziJJf67ac24TcNKAn+Hw1M/JnyM+8Q8bn0/xp6wcfaXP5bc0tHNWeoX23FI
aPBtRYOygiplSS/GlO89DcImQ7hshiWgoPdYYTDAUCVFz+EN+gmCEnzi2r74haWP
n2FLdzf0RnZD5LtpwpXmFo86N0rjxDwLIL8efYnjnkyIi/9s2WFTB+GsejMEq6PY
3gZ9ujcV0IvIi8I/mHwqHW2TqW6X1yYR+mfxXXzL7Iv4gqV/qs4SlFjfg04Pgv93
Nv9RMMQbLAwmPV4ei/TX5uCqD32/FnFWRiRLb4WDRDGr0jyyWk4iaR7HdiCpnut3
5j0qewcxR9A0z5P4CR5B7SoEmlhAYFBa7TzSrgwtWGjRlEmPlE2vOJeg28+0Jzh1
hlWzJ87ePChCaECYQ6gotktVV4enG/6SuUst7uG5ABlzb/fl/mihqFZlNOnyXKfc
DIVKGJdj6Cy3aDdHuD60FiNgT6b4sz2zA0ZBevVodxR5P6bUfQ3vPKMi4/P5kjwn
6r9oCckSGvYFnKs0CSzAhWNPPsB1Bx/Vyq/HlDcRZlHpdrMuaaKiQ+A7jDEaSd3W
joeqJPzoZAkSv+9jVCL9Q4tjWWDV4qkfbfQjCyX76FV2uUvA7GrifV53yDnqqbE/
u06lvmDSF+C5NcV8YwAahGHZYjZ8Kf6uGN/Gv9HX668a6KDyaPMgbTi3aAlGM975
XsVeDUurXzOtyHfyJgF/g25k4oJCuGNbSDJ7t9t8QosQOb48ukFRNDjuo3JM3u59
3CdPYPHjzXxHN7y+1VOM+gc7TY6NhxQR2W12Py4H/9XXos/dOI0797N0nJD7FDiW
hy6NwxJUYLZLE0lUc1ZHaedmIEQurBV6xWvNUmGm8I/IK12It3Rp2CQrIdgsxTO7
jzQT0PEKPjy44s0t+MJ5lfZ2NsX+bg2uiommRiseipPqWfL7sIRWuO4gP7ejnJM+
iWZ+lSKNjywGkxDBMbjAauRGgB6IV5kvntVayz7Di3YldWaMGC5aanRzBZWYm5gk
8DPEbpDD2bjVkc1U2NwLkNMYL0xp6pwYgKCFBc5sYflAejr0svhDNgIJliOWrpi2
GEM04XjEx9Xz5xJ+91KhOWE/1pU4/vfYHi/UrdEOTiDhKJaMpd9WPiPmZBb5zGwP
OagdF7MJgiHq9fYmWyrdS/spa8tkHd62HKqTrsl5t7mUrQuran9ohhC2X5XXyEyu
T/jRwL4DhIr7iy8wP/aKP8ZU82esqF6ljugZP6/8p4kowv47eGSetXgmTjIwH44Y
pw4iSJb3KN8KmuuhpfhO4LZUNDJi2JxPmrxFdWpINVHMKHbY3peRd3K0OYwnR/zG
mhuTF2JNgsZLS+R/2LvwQVoavvRBAfyd5LCSUgxVt7da04Ne/SruImOiTEpotPIe
C33sanQkvXbVvkgfyLxMkQJfyMcfY0/t3uyGWMxWeLIMrb/4nyK3DuOIP2WCAxaK
4Q0AyEydweMAA2W/VM6fN/WGDq5BaEMohyffdsAs3n6gi3u+/d74m2Rik1P/VM7b
2XDNhNxpbuKmVaeIXE4Ya0sudzjpunlwSAMid7joodT0ym8vlFuvlaU87P9OT4Ni
LKkxwv9LXAJ9i97IEI279FRT7diPfDjB76RDJTwKZgBXrdJjcROKp0m8cf+uyyKY
BLegc47Mf6YxlX7DUhlhvGe2ovx0KvAhrK0n+0BuvCvSvrvPgIl6nlfCTVzeXCZ0
XtN/ipa7HLOFbL3Ot3eH4ehiaAIWlITfF08XcITZWlwiH2qGyvnlZNusbr/8lm8p
UE5Rr8kLaiKjbRC+dXc9Kjd0jWzGkRmd/KKdhiyAjwhR2C+unN2PXS1bNVVSFTxQ
lrFHIP95QQnWEhUMSmocGfne4YCiaSitdkhltu0BJJGSlRFeEVP/idsSkzw1pAn6
A+p1a3/PshkUnvMH6lsJyMug/zU0y+0Y8JPQSAd6St4MIDKGOKHMrVAcp3bL/SUh
rYLUdYaEZkw8bwtDNOgwmecaRLmu/QW5+tbmXCZXbyZgasYfVy7CB+v9PTYHcjuF
0l/sJeuEK2rhJBsI1mUkqlFSBTGwhmLFUvWbId2EaqLADzUNWcLJXz9V1WEHsQeI
Zo2oURKVYdFIgssNDuP0NOB3Y/8gwp3iL+K/neaZ6N7TR33p+xdZIXV8oIgHE/WD
+QVYkf8zV1jgBRMNeULKZF+LdYb8bT6YY54X/ljR/VuewN+PyFqyH8BTFbB7jIyx
HUHQ1ml8wQXsBqKqRCw3xmQbKuSWN0fKTKeBNyS0hgBHb17oX9jBcNk1W0nndaXQ
3rlyZP4epJ8QwHsplTd4c+IuS/I2sS7giHmgRNsnPiM7YuE/jYziU9IegjZLgxan
ym0aMBGP5N94JMncz0wnOTgisVIwZnZR6tAP5C1n1hbX5bzuqExRCK6V6llLqQKW
NSRCVaIfGDfMqSDWztvkmxZX1yIQ5l6iEi/qWyhk80cQVUogUYCuEG1GR+s4Jsq4
XG4vKBWIFIOwDzfxaRssylZGtUtxLQmPgQknSOnHk0h8wlzrhoLlQhnFt0Jqdd1N
q68vAGcDJD7ih+XbunCkMFT6XXbY0Pqp+0BdtSqOdDmM/xKHVtfFR4/RDDsnhMVi
a+REDPJq2PvaqIy6sBXpHVaRUzeoW/L3ipitnCjUagxt3+zAoJY4b/TWwCNycVB7
CEJTzWPbTgAJqO8ApvFWLnpVh1MdTHWgpRH8faG7YJ9qgIPUWYzeb4hwFeMFDqar
lFkYyHLJjs+ppAMgK0990hMbsElBaCAsg70yni/pVAH9+nZ/ZWuNMYBKfI4CoiBA
82xgAx+FdX43PjwauPNxKR2GCcj1r898QuR7t1wkYuvcYVucvyGiTFuroK/Oq0yf
oTS9tv+i1ggLlgHp9jLPBgQuqs9a7/pKlFZRkC3tV9Fp+pl2FZ4BOHlLJK8U2rTu
irso8E2i6wjvV7mwqeO20sqoPge/dsbRoKeQ1ONp+CFtyLWHBeGbY2TqCqbnE3+3
gUknGBRT7KS75QL8VA6CuT6um43avNbVrx5mc9ju7t1nNWEWteOcJrb/b2m47uUs
zrqgB3Tj2ntiNP1azk0sdQXiW2GfD3BTEZsGlIjPEfChq0rNFdiyEAa70NVtLHYv
htTTh5PyAJHsbQ2ywi7HwYpx0vSH+UjklxtT42C5rreyDYcGrOVOfLdRBVbvZRnF
B70zPat25yICZw7GPeKNMPoIyxBQ4jNfEft66oMtQRSPih6h9Igfbcfy31xfVhzD
qU/ic2/rIN2LvghZ9wtDqtVDSr1wBLGzmdM2dh1+lDCoM34SGUYsE2TWrCx4a1/g
iPpgdMu3zKO6gTe5/OLjv/ewoHoQmBdrlMLQvRK+9bX970u8KqtmueAXVL2/ySOf
m7W+D2Vg/4ahMA8PDa6gY6X6mXbKoMQtE8PrLhO7x/dAEVQlLKXWeYt1CVyDw6VL
KCe/47SLuZJ3TJTSKl8cwBaPk9+ghY+LJV5hxSE8P5hgX9BAyO6bDZlWie4qDWc4
aiSjrXdXsmYdRMFOFKcXAT1afO5h4xf1VNRKSmIi2DRPVOlqTRrOoFJD4GGxRi3a
0O20rVhpXzXYV0Xslprbsadk5EA0KUDbXceQnIUZFS4eGNzwkYEUt0LHf1RZcl3G
ALjKw+rfGTZO3PrxRjXfOnQiXUXR+tw1AXWNoXIfw1p5d/huYWYSXkBMP8xWl0+Z
V/lI/ehL/1ZegreKs4L2rSO4rS9WOU8pOdq5f6x3gkJjBuzeFQlhrhzIroGtgAbA
1uWpMK60zWTi5iBJOQG9T24pKz/gv1AZZZE2gy9MPuTSID4rS7m1FHjMSvSkiVst
0cZNC/1unsZsyfoc2XGFo5PspxzJMfNMYwl+ZqR+tBR4J02GTdxt5il32LI40Xph
jK/f6a4if5VrBmzY5qzzhQtQeQFTQ9fS+QECRG1+oJr8M+ntxB2Cia78Gtz++t8m
OpVMq8xk7BCVn3Gt5Bz6eCkTj/+rVUtkDAJOXgAlqlosbIOY9RZ3WSCEvoGcHDuz
MfsAAKG0HFJvVF7Pls2/BwvIITgVosqp+C+QbAoLOIKa8T8DC/R6sH71VXdIC7wi
PxRFzFnGFZIcshtWd1YXXLMrus9HPeDaBavO6/ISgdYG1il+X+j8GplOCvwiyb2U
Kvhz0jYvAo/AfyYqttNixPkOir0vaMSTbFMfnoZb/GaKBiXAjnABtYebQ+dG9LsI
tQ5CVCqRDBvpc4Z5z0xyCgnA8uIKuApQWWPmWJ2WgyR5mNisT9OXXXQUA6QsVT3E
4UeidU4hti2yEIirsx5m2d3lpljeNMjE8O0Ns5j3jjMMlXsygmBEFZswFmlsM4q1
v3Kmty9RYxfXaLds3L68DvcVWillcil6ICv43PHfX6OwwCYRzgOwpqDXNMH7rsXW
TG07NM9cPNyxTfo/kbZffS7axRGoiA1wKyZDXD2V2wH/C66tu91W6lc96yh0I8MH
k/0Vx0HvPisjEO61tER+NMyY5PdmzLa5qpc9xOWdIsnDLw1zLc1B8WitS8Zwu+rF
GRi4QMc0Ijt5d3spnsuhSBG9lPRjUiQxKYtPcthyYm++jHzD/K2HDRcSTiH8/9VF
eYpkFVKXAB/wwTc4KMSNn5jGKOiqjyYY0kSvF+0fWcew3JSQl/8Se02SXh6lcnyw
dh2vZldRCZuTnRvWmL2YHLweNWWYtvUAKx4J9bdUwOci4IoIQqTCg/y9LEFwFUcy
UIfxZRQJnqzje+B+zvG9fQzLeoUfNl/Wn8Bhi70v7BQVqSPJVdcH2JQJVlz5mXvs
rsq8bshs+R71vQryCyh4DEwgcMT5Y/k0pNJ2RaWs+nvZ8EAQDdnAzfaaXvRv7g62
AuYrJqKmu+qBP2R7WBFPTtz6/6YMbKl9yhM7TB7rc05LThdzCcxz2OKB0pa+fCEh
CVHpv97FA5lGcRfegDiP4Tsjmwrz1GN2OCW1R0EA1+Me7stiOy1vzu2C8su1HDTq
oXmYQNhabrA8fk+TmEH4rNqmEivwlTwOAZ5vqbOJyxym+PpZTEUi9KEhXcrtTlOS
rWQ1sRioAbwqKx0LZarHniK0KVlC90fmEkI5oG/6xz4LEVv4WRZHKc9U6cqywVxR
KK5Jj9RRnDs5zljgDKzDRRCk/pkinqs5oJ1beftoJ/U1oBhnXSU1qUk1Mt9qvFHp
OManVAsWdANXAjBKmr90jzVc+tAvaBTIFqC216L/3xegCUpkjXrCeFlYB+jFut9o
ulpsVIXReh1D+Gvk94uIHZyyy1IdiTTWknvNlD74o48xh+m+AapUUaT6FVT11ODY
mAZRJ8IfIXpFVhSNLmVbOpljU/w6Ezw0EindidFebOIFfJjuyCMbOKjxcOr5UWMs
ntYCZHyHnLC5D93Ce82CCc4FuaKHLaZ26VHqx4myfnqmg4B0uW7Ev+fSj8oiJteH
EUYhCR/DGtBAkGdpQiB7nl7uCVmi54VDW/vdmf621Ue0KK+rzU3ixxhmqBvotpV3
JxNH/pNUV2/LP1Z/FV/PSnyudJvHcyinTWpLRWEHHrv620OqAijS0o2lCU72ADCW
HDNFMT0rUV0gvXwsBDUhID7umTJ3oW4vxhgEpgtmmJk6oUMpcLc555d5EnDdzkd/
8rRcYQGWxo7uRqlCYIJGLzD/odFdQiOyrS5F3qE+R2eEF87zk/lfLtwNzTMsr07m
nc+1kvMDgMigbJypYg0dNr6jvDiA8Zfr1achnvNC74P4xjFl8SqJP1wWWSExBs9/
8Ecy5zaJsbBX3aoApJSscN4NuKnxPn14hxTA7FzAQisNBEbVAHHdK9IGoF1YrhYR
pgOkbgCpdliuIS+/XrD37Kk047dRqOrxozSNzbNwYx84+ivCSP7bUHvt9ntxlYkh
o5b5pl7Bfu/KupakYI5kl6Qu4ME71DbB7TcbKqaPW5ezTPxJLEQq2YYDcBmwc6xA
NrZ/vubH2N6gZzXFRnKBPVVA51iu20QK8mIxyw1hgJ2yPCzubTuRyuf4B7M7Co8/
yjEDTJzhDs6Xq1UNB5b6nBUFjsIA28lyaD3GPuZxthHLV4Zs4vN87Apzn9PKdIWO
kg9blOytBpQCQYum3jPpK4/RG5bvYemzMBdYk+eNraOo32uTGDOhHlIJ2W5ws2e0
u1chTqREGYvHUKaMMpbWK8hS9mGXd34QcVG/zQD9NkltPuNcUi6XBC6buOogwf+j
CNCe8+awSr+IYjnJzgzyElBcf3dLsp5+AVgL+jznGJ9oMWoCYLk5uu/SwXo8EYYE
q9JnznBD/iMSwqveflBlVHlVrt8WARnWc1N4EBphSobBlLvu5xIjIM1Qw1bWt1jw
APdhAQMCp382keKM63sw2m7DMltFzIbI6zbPwYvAZMa4p3NULw1RldqL9vXZGyoi
qQZYIKZHgf1EeF6y2G2b+oO+8Q2WOTwBp+vlvMfjaxHgaJcQtJXuVdvrCi3DmHn4
xUq/n98yQmxx1W2+7zNLY+j+beWgIG2RyRz2AekQ5OOoJBX7AtTyCmEHZolRIBIW
5QDptAfvhS1JuyNqqgUlylAeChOIIsqD6ReKGFDblJrxI9ARIxzJttOWD/lLf3x1
rn7YThbwvK//oywOsVloL3mL7Ih2ywESJj6WQJhl9NBOhDgy3fxHer6QFt715U0i
8yVb3UHz7M7lFhIK1bmL5x8VMX5CsqqMGhP2vQdr2lrQ996RMjxnnNjY2iormwhg
yGjMAypI0PjHKisEpO2kVv+0+nGa8J3qH8coylUrVI2Uh8tyjIWd3By3xaDXvbOu
VTS6SRSTsePTunkII8GM5zjjTmqNkfIeK+dEu6b0xGog1Qxl8uG24Fe9bIK+a2cF
4K7zEat1K3uk2+05Aecrad/0L3Mwqrj/3MrXMnjPM2Sd+2SshEBeBpcwyARcgxEh
AE07kuYUISBfV2VIMMd6OTzbi2BlZiqcEy8oDETMyITg7RtlPlMqoJNgdCC+7W0r
J7mAAoW7F5dDeugCjL7wg9X6d00lua14fA57eOSGMCNf5bNnw9SkEOFjVipENyeg
hk66mESTCD5EhKbwBHdhzz6ilx1YOu2Kl/BB5BfK89IpeEqYYGn6Lu2DsAdXALsF
uYncCm3ob+VFNhCQqOjgAgiWNvWscBD6Nh9qorTx0JLIPzcYB++cvN2BYxcvV9mY
9yueljxFYU402/0uvs9qyhN4mnhJbhqF8//e/eVgwJySe8hSForPOpUnXzwS0HAl
sTKBes/gaBM8d8P4FN3Lsn92sNB5+a41MyROxbxtZL8PpgYwm9UYY3yvuJPdIr1+
X/CKXOZPA39JVbs9Mko859A7pWe4YuYUxv69hTFm1zI++zBf4Danyb6sme58FtWM
LKOnzLe5ah2C0MQ7VxGmSft6QfkTGjycqGpa26xh7Z0IsJlQ0ibRODz7KuR20rD/
AcnYOKRAeaNzUmVrS4Le+vTpj+4RrfJ1nvWK/tpWKVxmqjpIaRMMNLmSfcRDVHm4
AlIF9Bxwp/a5SuygR1doL8zZ9ePr7CVp5d92id1yTqYaaopXjEZs8SF+4g6LnUGO
OPEZLl34NVvcMsIoNJfgbmd7R9iY6qHyuVHckckmM6ZO+gImTSIH9lalbVPWmKnp
QRzVAi7CtYJCctUL6DV5Yjd6OONlED4MGq/XFeIMv/nF4nbqRpV6iOP1oGb74CWC
+4RR1wr2QjPQ9uoK2JP5S+0K1MkpubN2zMaJbPmChKSmVhZs8+JRcSG7BBUu04p7
Cxq+J2OKLaUNoyH1L4OyA4VL25m05dzqc4adedghPbqsfgHdp3cYf3Nl2vTt1nIA
BtKKB0YK0w7SLdXwAONM5HDt9ZonDeieUqNMO+W2yUkD22VS81nyR9pqEdnLLwX1
AD6IEgQdDcl8cpddCPG9CAsk3odnvjdMLf31SsG3xlcYGzvc78+rLVhAaN/d566Y
pkc0E4XgieRl8nV1yNwHPeICI0sM/lRdT1ATVdJANMqxEzFPcBtBSw0RmbdPI4Pe
X0Waj0YIlWYNtXsdcIk2bKqPuqv5Qn4+Xujh+Twp2ZMzFne8PcEpzDzs6fFC4Vn1
89rKJtV1pqE3bsIr0hrCIqrYX/G/n4nT1w0/ev9+DJuwqf+lEiOKjDqPkYQ4UBgv
3okXWi3Y4x7uf/XNGPH7epe5FRHry981x60+NvRpTamQguF4pocAMZ2uOKeaSZpF
bSDyPZC0rmhFdeUINE1P7wofxzdv8YeG6GcUx76aSmpDWob8gu0WcwkG1zqfU6Lc
5K1CAaBSiMLahKOIr8QoexbYQEECzf8szUzVoJwtLN7sf/zpYPab5GGZkR0hD9QP
fRJMX5j5EAmGCr3EgU5AnEB1edwmNnhdru1NXIPxw1W3ElG65deJz0aZlMQN6iHR
o0l6cM4oXRH5T/MxfDho4RkL0vlKD2YF0pmTd6inKHI40zELPLUoPZn89Z0r9rEb
iigZJys3fQzzAF6ffoawUqI8QtCKxSKb4dezknYjEB5ew4aJLrqqhhIqXERNO1fS
3GqBo7g1qN4sIh2uPtTstSev67SG/pKHVZTFdN0UTL/smBb0fHlTbPiS8dMHxkz+
BIyZde/8AwQZzVRCg3ESdyAWi8Uubwt9i7eB9vviP+woLEA4gkNotUI2/Q+mWeiJ
Ul+i5FUwvzw1kWeihJblhB6SR5iJ8omArCJXB9qWwSAjfEYvK6nW7VPHNZN4xvC8
k5vqFdEkbsSMxrJRvhdfrob+XH+oHst59VKiPGV1lfVpmTj5N+TEpKAojhxsthdw
AfjmVsaI6nXaMSue4JmHmXF4XxwQPLhbYw2TG8XAMNvZBKCmTQ5NE09nXWEiRBQ8
cS9SQt2qhyE+9+UjIVFFuOwno7fQb9VNav+8zyfqhiEckIK9WvVRoDb4mxXDqThS
OYlA4XAZmG75BSoSfGy+LTuY4Zj44F+iZr/G/ysTEkDlP06SBEJ8lSEwIceAXvkH
l7TvH7vi2YyeeQwpl+Q7i84mXoTTMyIztlBywMTUHGNX5bIAPuawj3qvZGx+fcDT
xHiZ/urCEFQUCzh6CnYKgxeIVuv4KY2spN84z3Bn+Qv7AZdS2gMa4chIJ8ovHDnb
Y3pBiW31O0EF9ZlLHJdqu5FpipTjZwkxDHk7+tG4C7pYpgarp6Qs5vlOieGQ5bhO
G8Ww5xggKvmNSxnRpWp7z2rQCXu2kMRYCHpUG1spiihlEb6h1ilsuXL3gJEyXnPn
0McFCuK00TvV8EQi7iGezFnqUgGvRSCv1l4XaUUfT354F7PiiIn8h4vr6JnxJNgw
DhZVr1h7qEK/h4FuD0eMgUpGFCTCuKxE3TgPaXnnr3+c1MfsoRw42I7uafMiVDtS
42OWCDPm0HoudTWh7tqI3zv1HGv+8V/9F3PvdZ5Fo8HRB1YaVya98fCMcG2/akJR
zz/jw1RKx3/99gKIN1123PQv8PAAAMhIs+RRjB9cnlqgXbaSF4eVXTAWOm/OA+uK
r6XRO/O8W1BnxO2bgXJh53NLipRwU+OzYwLKn3MJ8ZwJwKA5M8izyp/7IDPAWf+d
wEbLXjrQYJAPNt5GcyzggvzJRLdM7txt+bDg94ngjMKyVoObI/h4Uj7g/z88D9uM
XyVUYodkXn5vv5s1Vmmq+dBRDxkl7UnipDT26lBvOJSAQAUzknmyviiLGntIcARI
lkNVAAE1t5R+mRtIqPZkQ7TrVDv2p0EVklU9HBguT+1GxCdx4fW9DzaQJFxSx/Ky
Q6DyWHGJ6fC0dHgf5ny4kWPPubgEKcuvIyNWrh1t1PF7MjfThVQJU4tQGep319qR
oIWk7Av88DulXhQEOahNDYp6ovzbrBjaIehYjKhPuFY03OaeACaWK0TCxSnM4ucX
fpy5Hn1ZyXT3Q3w8nOIblqvJWtFYd161Q5d4FRi0DPyLqeDFrAKkiVYNE8bqkZgJ
Tqwhf5kp49Ya8V9fNc0PfOxTu1xOcljD2sVrXVJ34DxKpmj2pRmmMWIAL+kbYJC6
A8Q+51gCcnYTrRNRb8onqcZ52i/hKyLZdFgpt84JmMFfovshqgD2dQRBIRlzCmHQ
VaCC8q8VOmIVOTdnHR6M847AD5ec3mlhBorXFypYqq/nJWxvF6ilTM1ISkJYyKdB
C1fc3fx9PDmYY1TtGsaQokY45Kqb7NqGnddrN4di4fugZi9SD/XjWaOxLJccGfYL
68mOOHScBsvFHGudue/TQiSAMa8/7mFCbWnf4WLKozy8EyL3d7JJHL/UE/SLvQpA
ma0z7IBs9Elup0zdratMD4iPrOwbxQe/tE7imUMxargaNK/mIMCAq5eYcgl7WogM
HL24R+jxZQk6aglaaNk0YnniUR1bYU53P55/ihek1whFxn2EuzwdYlZsup7Q4rbD
VLP4bngudKiOuZFPafrVYQgq2WdSPXwHE4EVNhfetJnxvQuPE8SD77DrIQVnLvRk
TBbfu0ZcYe4yxACcOIuD7SBBkHhc9RIMmbr9Xxr0J/Ofqq8YonbOea+fCaqBKVl6
s0PWYa+n/uYG7H7URsdyI0sDfmLPGs/OoVT0ImghGBTMBXCunrVQpsqZI6nXihBY
mNZwW74LLT0OCkIHlz6a4uSS6cf+DdjVZq5lOlzp1her6oKUbFO5SLNRvo18P+9L
diFKzVpvuToi0Rf4Yg8/pJMVM6YwmWGnCql2Yi32Orersp+wAjfkgOfDUGWiQVCD
bNIpbIrHWif5gexg7HiO08B8g5BioD3XK54wfgtbnYpYV2zhBGLPJuuPPNpj8cwR
QTiWUx9aIeXc0KyzP9ZCLxxUyLPKEW36piLQ6QiZZOhxxikv1lKaRq6xEOl2rLSL
H/wompZoqn6zXCUjfydpepo9foJYP0XEimO4L1+qHeDSRg42dnyfqbFq/fgnU+1G
zPGVl6JObZrxVPM6n9i5CFI7Xhbk8yt10Ic9rygWJXQ45J+cvdU7kGQHU7Ct9N9L
42FiU7ZehVm8eCDGcizaZlKeM0VSNkbn2PS6OIfXAGAqwtbdHGsiE0veSPZBkavd
J1/Ef35f8FdyhKljmTF0RS+6K0ubfufD8DKQgQXpyH4jEhUdvFZjb9QJ7ZQ0EZVL
lh3zV2RZWcjfDsVrI7P5mUUvkwLIK49rZByNmW9nXUmrZm3ilTJsk0gaHX/MomVW
pz1PcjBzS4XQ/hf5XkY3mIhk0QBYFy2q9nrAEDrhHa1i7jztmCBEvHYNkCX4h1Mw
va4hewrttklpTQypNvp+V3vqPO/Ngsyurlq3hum33QC8unwbsBMzG0EmSvOwo76b
ze8iXYYOwXtJkjwZmE36ksVSouw4zrO2dyoYoRC/Y6spGijMZktnr5iDF28ACPTU
Uht58jdi8WItBod1mKO2X3W6Wkqm+lWPIkwBUbfFvgDAa/IQSVNZboYAQmASgMNZ
n8mk3ctjiEeiqHRxTSXdfcOMcSrNdDfmVbuQ3q4sHlr1duGIzeSsj4wQiEeHpb/n
uQYwBtXJP4f4gh8DFdhJP/oaKvhu+ShcQvlIzggBqdWZvmo7M7iGWWuA9Efz+MDl
y2Y70Nb7mRN1YEkPg4h5qb5wDBPX2MlnDIr8gbBV/M1hvIYUHhqt0qGr/h1BZ9iF
YqtKKfVrlOtuSK4wl937yfNis41K4+B90cwYTVcLnxwF0tg2uiV41v1aKlUhSfD5
bEFQwOzZNK+k/fhX45LUn+9CAmfUgbteJWAKYq9aNwPKC+yfwOyqtZHWut7mbkS7
Rxg9vxuD9t2gnQgIGmCrnMFX06dVqXA61vdI+71SjhRy1J59w5ScGF5tljQ2lVLY
UuAoRfDpBVeubL6/9be9DryQgQrIdRkLJ6tKFFroHpYDjMROCEWA/i5eBJd6EyPU
uO0aXJio05GWlrLfJg/ydb3sWWA3TnY540cIFxfe9FxI4v2v2aIIcn9IBQzc/y1Y
D0hnllYJHXJbbmxXQzxiHeHfb60C2rdeAGA3FzHOqHlAgvR5kR4KkaK+TMs2kmtm
Sxzn3vUBjPrwrTg/0vCTFJC8HZQi9vHrAS7m8czJRByb4DdlxJwc990mG3ZMCbLR
T/l2FJs3MvIOY0UlouMsm2AKZi+r5ljge3y2XWXEl7F0EsTmqqldHFG9nAtKPNyL
4TdztDhLiKmEqdoqIa8hal+my1sCklY26paMXSNa/uXNvL4lL8o1HfQu6dvfm2wz
MbmzVo+u+nC7Nx3J6s2aBa37hVPLpNzsXwA3smYkY1SfEnbCoGI2rF5l48H/K470
nymCBmJnK+uQYWC8ziJJ5uX5qbChaBX4wIQ/fpapHsog2USXFhVFshgs0V+6UGaz
Po71H7zbhjktoQsnITnjwFqySTni3hE8tMlc5LJtLaHXlFQJIdP65g7ttKknze6t
kxdch5N8IbmD1oL6EuDYPWQ3jTAyRfqzPDvntA8txmmhuHy4tZ+34nagv2wc5hlb
9strfghnHiEwAEKn4NCPW7o+Zk+oTkx+vdC7VBkfo9fm7tbuGt+TCUEl1tba4WEH
yCX+WK85G0pVea4s282enwg8W59cTf3GStVZDBD7LjPNLSne2GF0mZjvoonWHtG+
gfTO7GbQbDcxJ0G0Dhq1m5wymQMjTDTy/XIFnSDjOqGWBj+kofmejVDFpVYAbpcz
CXCnHTT7Bs6cKpcczE2elonObZD710hWgw5WLY/Oy8ow57w2EcKaCtmUEcl0bCIE
t5rHuY2WKABThbVVwbMZwKAVbxdmEalfwgA0H5JUwbpXziC5VSyE3FUgfoemdGzD
9kkCxzjqVdr1+UqhsrWe1+dgc1wL9fn2jpsSYr7GEbYLzMBHT7v1qZtGJ4+vQ8W2
9/Y+7uWm2lRMce0pyHze/TfIwiui6LboDSeEyibSb8P7pBUoLJvPVUhvyn+3b4+b
gRePxUR+dUx8AHugNW+lAjIa1fyYe1KRh7z6HG/dHM7VblmnbftPmf527MgnqRcB
Mi3HC+7Wri50wyEP4keVbFxMspGnBD0KQCZqv1kBGZ9eux+QDxU6/PlJPGTQP3Nz
WRovReBlaDEsMMydGN7garJ1HUA2KI0kFN8k0eXhOViCnc4IVwNHfvrxWu/7Zkmb
n0scoUTXJkpAwotLtbNWUBWR6iCxCuTtJrD44LtiqvXlm9KRGMsJqdJI90bp7kbn
HknoWSum3KfPTaMqVsJx7WnNQIISDj3u+/CiFXyW9OFnfCj3MFGxlbgumiMYUsz8
5mJgw3VHN3GpdW5mnPGeC7o31dYX1bTL65e4E6UJl+VCcvPl2F6Q7CeIu4SR6Ypc
mrrirmsQYLUYmqsdPUClWVTif38lFDCMFd12343w1rZlNdBJdtzappQhqpM8OCvO
LAH0FvoTC1Z8faAiujRlrRZHxcYMjXeaZhbPticp+ddc/E3WHbQOnYbj9WL0L7Dy
P1UiyjJwtfcENDOB77mjkBlykcXBbmjQK2+DpYJNsSLLAsAZicCldBpFYi6IRnoM
1RTxh/PLyPckTKTKDQnidEyU1UXvGOnv1VsJO/hF7TSO3VEsKJ+Hx5/3yyEnNK+7
xUAaZuTNShBxUz5N7ybT0u7mhEVReeU0AHn2wqir9+M2L7k9zTHpTLATC0KCVgdM
fhTgl08BTw0pg8vClI6D7Z6PRfqU5hE5BRAIhL7fWuVw8ygCYiz3BWgPJpFPwKpS
LjPLwkzF+zNEKpirNrG0PIHcFzoVDmM0EdKz037bBG2ZPDZb7UywPYAsJ/HZhyHN
wfCzpodHXpXndthrMkkqTH+BxHtjl7A92VJ5IYKtd+N4R7OhQbI03tSSV2b7FA7O
sez2jdH7/3Oy+/kXqz0yuIn1xyzdz8svgfxl/GRrsvatKYU9j7Wb43bxyws7cL02
uYSrYxHFhgBkqwI2IDS3/1xnUIdIofA/2KAJmTBtU6kOxISzPKeMf51AXyqd/LJ4
0YY8vszWDVrY/kRV8dqnZPGrqGSKM0UY2al/vt8fVQC0CvZGzsavtRn3wTi54aBH
eROLv50IzZ4+gwrwsH12G2qY9eGKyvuWMjoz7sjn8i0pb8+idrJJIgH9Mh+0zsjE
3Hq1LvgoQD8zUA5Ew3294IXO0Rgn9pgjjygx1DjmvRk1e20of9nhhePJ4Wvj7Lch
bDJ44Qg3zi6CizGR2dqDqD0obscQTObrTjPCOVMePrZ3uu7bbZMV5uxiTerKZJkC
J9R6jXoeZ4sgOhXPG8GVeCmFXZxEGTIPp4lzs63q8JcBxJluYHKpCtMFd4Bj2prK
KVx4a4r2TzaRmb2lS14UuikT0GY4P01B0oUCd1fHY7umUTg2rxy25dCCdHAmkCcL
LirPVGfQosr8E/l3ddVU148tbZHvEHTFH9gET7jidxZ7+GNCaJT6xg9PowhYrVf+
31ekf6ZbaWCHcN7l98eb8owQBF9HUjGTbH/LQz8I7Ec1wlDTG5hcz8+oVJ75p5gH
VHK6rq+yRN5W8m3+Zz3iYC2gTH9EcQkrmM9XFSuxuOp1HZ1ToTFinsdgLutAwKzo
Qfubgy17E98MivYmMcuj8m8VljGQDb17qFo3s0c/zsY/bU6MmV6G/pid7hWLVVj1
L/I9KppmbzPnX6Nf72mmqhIGTTTpq6PvkfYEM+J/bRj7rClCGUsXncIrbf7YdoIC
n/t9O+cXiqDIV3Fd5WREJGBYNqBiT2bR3lrYHzEtfU9ps9O/O+8Ycf9E5YtATWnq
jZg7wKbBferNhMLar0rc49SWxx70/j2dwCbnM26O98fTnDU3h2fVVsZF0Dr9OpBY
RtAkgU17KKbIsjmZE6AKaAbOqV0d9Opf8NfAe+Q/fO/lsEggfFahRuJB4sCd4Rs5
XKNgNEkA+VGP6sXMJF22dDwNQAg4Zr2cIuax7w8V0OCvWYT3ylE5IknV3gWYUYWt
SGqQ0Mwv2ug2pbnW6Ar8jIKruVhiTPJtG4wmdEk5y6wbrXHrFLXK8xjWq/mN9iKz
7w0Lyg8jyI/3NkEtM0vK7bvTq71v1vX6CxmVlQANmC+top4KMC9DLVEuAF4a2Z9i
7SqLAhJIEUsBBGLPLGeUgtvlZ7KOMrj24tI9bBEmvbX3oAmtW9HaAFoQSTNZT4x3
y9O8ZQg5KA4L46k4auoyb/p1kfl04/2Uoms7V2XIe94rWdaAoWZEBgKM4b4SAm6C
ffgJxpMtRZixUiBY6hs995KeACUyFiKmMSmwEk6vm6NbxrSCiJa1Y+deq+a1SToL
3Avv2awuzOptnp22itMTd57aM3VwdbNotUE/s2uZ4kIyoUhcIN1oL0czBE2/DYUh
M+Z+RGZjOlFUVTQOxdgaYC1ESBXIO30obOOte14m9BSkxlxIuWcHMkhrB8lY1LT6
cr7uKe09Qgzb7DKtb9iaIH6iJQR1mKlQRj7LYXm/dUEZhDePCbYp+czu6O7+XR/K
3OaiIB3FW3P+KG95P1Dyi9EU/p/zh2yz928GmxLwtwh6BhPIJ6j60vCh7TUqAl1e
OQLJf1ql9mucCcbFBg960XeO2iD1cqPph/FgydWDjQyCJ3vQ1xSX3orZekmBPL1H
eeMUjbcqWlGW+bCFuPQ6H/2992lt0Ci4frY6Z8cZBI/rVhA3VtSft5FT5gtFlxAJ
ZppLiQnXcwtuspjMdLymiBlA/6rYHeXELQmYQoYlpIy+HgpObqoQuy8U4pyam1zj
bVIR2HuXZOzIh63egrBMhhWPw1qy8M18O8+AE8Y4q20srJkM6JLLZJiNQeoMzw31
ctWzNrZLzTyY0jLs/MAs7C6eBOsPUWAnVVjjvFapd9FAEVAs3vSlrB7TiwmiB273
eTcBp3XUS5QtGHhtV8ow9lYRiDU4K5bB74fL2VBHpWahszfmxUe40Hb4N11aq0DM
FPyl7g7XNWdlRWtNBp5LHbL4tnmmJ896WEws3O2FsVHdOtIk15vxYqCWj1XZZu5w
FDwlNNGnSDuAFeQeyTF2sq2hT4iYD6B/Jla9JfJxkyucBpuynL3A1Xx1eL9bSzNT
W9bGGHaqq7mBLUxAMfBCylJqCA2bzb72QwJbyqVUlD7bOcOmIO0G9n/GyN00TQUr
e36zpPpKnN5U/DlmC9TlHuWkCeZI1bAtDpXcHtlLs87gPYs9ksQwK6G3i6Yf3bi3
b6tcpxrWKbxHQl67xMQyiB7dEqe4LFh/ywcPkoPRyo+WsZLt7aZsqzlDs93Kj180
NqeIhUKhH8A9rGioZLKU5Uihwp6MGJqIATouGkdEGqmJgqf0eKsYERUCyWtJ1eyL
0GT8QWN1U6YBKV6UawBrgYYrCs5ys7GhK0GAomBoNxJdqwK2f8B3NpvtjUIe9zIL
TCfm/cmVDMUE+S1+BSi/kwHLlMufStx1DFTL5WYBu/QmlfLX1woG8Eg1c8CREPus
/rsTeUh9ay7n0GzF74e8cWOnFNRKtKFbmZCGmHQQX54/T4rUfOQmAuLyQIRHu8wP
X5SraHQDAUoVPKxCsHZjcu2YGpw47u6DlQ6PB7qrR4D/igtcKLggKE9nhu1i5se1
ArMpS9vHPNAJXekD5+WLkg5tdZboWUehUFOAVPRNkOj/haT7rO6Uh1EO9gk0UiQ9
jQPQV4ri8KWpAhgZCXnz3QwB0O0Kn5Qv+OBtm+2IhjUS6GdAauzfCBy6h35DZOUA
CP+/+ueKA78STTwWZ0mWunK38YgrTQVHZv5qy6OhHfhNspM4qpbk4Irbv9R6aQ/D
RxAO7nZLBvXlBKh/b9p2/zm+RFZOIbXlxuh8f0T5CuzkGldKpqnsqXF+KD4s6KYi
MUJuF2TxY9Ckhlm+4pqy/S6ZVRK0EX1GLvATJYNkp+LXHsh7NvHkqEm3BYrUAGXP
VDBC/xKqNn5eIZmkHh0jUbjD+oTBdiDeavvrwN42tDHSAjv/KYYmOhaTTy6IFylP
+k+WHnLl6oztjSPGM9LmcRFDwNgtaw5CUN1FgWhTnlHRz8XSPLG8t6CNy455KSp3
r66lPTz6B4F701RWuqoHzd94hvSJeZKeJ8mTVMD4KdtM1u24eh9+4xj2OPwVHbwA
JFrSOR49XW7+YXjRbPp5gy+24nD1us3W86ORD0gx5QZ9Ndoe+c6poi7QsWRNfZ1V
HTK7gx9y+m9CrRpXSshGQdQKfCq1yawg9DF6V9w0ikx6j7CfqEt0D1/ac0vA5Yz8
nCU7PNDvEXSmHPMsvGnRYLBfLEuLuc4Q1hQSJi9jnhahoETTm0MkVorIEOUC7T3F
O+3qM/WMAMfAvudE3lkEz+sl3UxB0ymsAf2xoeGJ8gq3o4f4yL11qI3lLS7b+J+q
8kmQasWAVkuK4qmV7wgg2N+TftLEzHZhT5MpJVmVyu9JL7LZsicbooWWeFK8qxkb
PcEsEhMs9dHAioI6ZEJfjJKQS7HItnKTVrxbJUhTvSyEqVZHVL6k8/SppmdAG5Hx
z5GRayBY53man9ui2mHmQSiruG3TkoXWVuZmTZzAaA5t/Dbaq/ij0+k+B+ZT9Evk
kUV+NYorN63gSJeyM+qFEQtAQMmSH2IWzDPKvNPJ8ubm6ZlU2TX6Ry2uQVq3ydvW
gNEO6zewF9/F4rsdvvT9OS0Q6IILicH7HkSU6xa27jA2rgXGoV7D8G9JNGTWNC2L
g7ZGYLhGMhaR9zkKttYuZeczq1qAF1O64rzWbEEsSp4zFFvMvucXKThL7pTzh/z6
kfZFQJfsswIk/wDuY5ASXT6VhoTHkvYEYtyUMikUczLSJ/8qEnh4Zosd8Ti7UB5R
I/ZedEZr7oc69rjyG7D1x+49OK0NrAMcQQc+u2TM40rZewYfHKGAdkxGCYAXT7pg
bkQUDwlIVkLLpJGcpZCp7Jqv8EaEMlXITIaud0ATC3GJ6QyMpxYZt4zkd9mkysg8
fLkRa9E1vRvSasd9iuDRUmb6L8D6oMntzweNxug8kff7Ei5e5LsxPEuGumeoCAk5
kG6fFzUgCKJEvSilRJ16RejbCfpq7nDSTg2woXN9sWtfZMP67HfbReQnIbkXiCX4
ZO+oeg50mPm5PYlablyJyLd2PwhaqUiT70WtddRIV3JOG3E+HZNwnL/6JsAh+A8Y
c7Y2eI16+b98op8n3oq2pO9NY4K9FxcroX/rDsA9/Vx9L9VrR45qPCwPS7/YQhv1
L7xNdjwR54vUx/xp8XGPRe7i1Hm2RIpt0TxiGx4fu3phubArp5UT3fbRQ9E96y7H
8zlA2cS39LpCaCm+jQWkgveEHALk5AoYhHQ8mJFZEfhXEURoV4j4HQyf+UOmvoqM
PyNisLy9ikBxg7ctOMlozX9bu1zWQ05FEgaTu2KBu6fanlbGGdZkYJXHed63CTIo
k92UHibIowtAG5kbmuoXjDNiU+ASFzdX3C1PEYc3eH/nFO1Quivafqjdi1AjlgVz
I7laUaecuq3HxSYIVk0Ghjw+TVZlp4+tSkHylrciInObwZbQQLfqjEV2gweYFrX2
iAlPzz4mG1ou0Gzj2pmSDogQ+su6z+X66cyIM6DBwAobsuHaxXgDD0yGIWAQeaiv
gAVCfVIHmOhVIDZctxbTitQGazlT4ajLTVUbfIi1J+/H2SQzZyhx1jwgLGlu6283
qIMvo/hCtKuy507S5R3x8KAukYsHqAOnDQozrDsa5v3HM2qDpaXrOJ2KJsSKlF5e
82z5QIzZWc3JSSOjYEDHfHw7n8IH3GY47kTvUVSpwLaqBpmK3vCZcbex77SZwKdO
fHFGA09/DKYSuFOYic334b/qVxb0IDOLhjvCm4Hw9eP4btTneRPqe5kBQdTl6mTt
WQV8LWLo/+y2KdAWbN+vq61vzkROUNk0yHdHvaWx34dlmxJB6rYvSwMyUripstY3
kKcs37h06gF6aoFlou0SONL7k/YQrir9xRjD6iiU1xWxa7YJarIJgOxHQU/Vskiv
Rv3LO7BnrYSKMJfYjyplog2a8pClCQk+v7ci6hj+De4CNb9jv8Sy+xtx5XcmBQmz
Iw0KmYyW1xFi6II0e+GVjIV2Ap9BXjstmu0O/9vrJmUfLo3KJHA38e4zndyWyQ4d
GHPrBZiLY9HZoswPZm7ASWN/cm+5meuuw1fpYa4OxWIBqPuu3BelC556ry5ZZ/ou
6vZ9A+Ub08BgT9/TU4m9TLybEdf5MC6+CkZ4wDzn+VwTGNJKsulYoBQ2E9UTDOLY
HzsKmtIZijkSgJ3FH8Oc6fP03Bytk8y9NVVPJrOt7iIRw8KKQhHOE4NLD4sfoHWU
TVMQ3Dk+0mdVfZXev+90UfLKuRBYaMEnyCfCXimkx6cNTgcG+++DWHhxjtrykQrT
qmTZNpfGzvs9mWSUS9dMsv/9MeW7QQM6sm0JxVFux0gLIx7rPIpC5fOUVITEACeI
F6jxFakMHufBaPQo2/JJO97vV+Vmm0yOvHpzXNpyeu20MoGHZbpwO5GhA4rbs030
geVxyfz7TsF6I59+5Hh6nWd4ZQtAPOYm/DdI0Z2ClE7bD7LepeQyL+9I1tZ5u1ro
qv5T9508L08rwxfBiqWlueMErVPhfzRhQbXsrPtjyjVj02qbqgiMNAR2CYOLbWoV
miT6Tui1Z2hOH7R7O5W66yjsNETT20TwXxto68vW6LvH6UbfXeOod+zNMeWN3tHE
7FaU7enIXpHESF2TXf7LH5sduqcrryQZW+/GiX5xEEpjQWtWK5VXbNN4Oz8QtCQK
cM6zGX9PAV+qntO8GF5L3AbrMHj6mfRiI8X4KKiNwizS1LAb7mdpDuMtdb77OshQ
SatRw+jwAmcCYTZwzChxCfGuVbg1XzL7zbT5/kHA0pJ55hTp0ph3gMTO3Jy8KGtn
llNx/UVCmcFaep2PMecY0TTyJnNBxtqjmQoALhEWhIEtxrycRK0tBIYaUq7cnhOq
XHS+NaJuBrvPpk9roNsOprjM0wlxOIT5RkMrWOCXH8qo9BmxICWDOpntNv5Y7hGl
/u3oaQgKh9+sVd8uF6EhoWpQSk0xlJbO1Fqt69Ke8mZN9thQj56Bj8mpvzCwJqz5
zombY3GruUWLAu8JkS6sqe7wm1a8Fc3DhZ3Qj3icuUHDj9YTnF17hN+dOMt/I1v5
na6RycWgcqcI5FQiO729Hxrga4Ym5L2jFDTTINZLf+qX4I4kuXsapGrwaGSVwkz8
8Q/+wUrOw9sRr9eBk3x9M7Pfr+JBOpn4VVwIjjATI7f18j9ww/RV4nShRJd21GiB
7B3tllBaXALidD08HK+WRSj81TDCn/VlCPkxda59r0+0jGOIiEiBwpAE4MFk0tij
AsrJ+JNUqxQD30+S2TNndvh7vxMpVpzZ4PhldQ8SYQNVIxXr0jpwuWsNywWr4s4f
pZ4nRK6XTsQrPHbvUr4xnGa7tdllSdvnDxedpzno/iTLZM/84mPXPYDS9eKk92FU
eCHljiBDLNEo1sQR1QzqrJeX6/VPnJNzKI3MdGbT5HQnSQ360JiqnWONAftJ3/dH
vibunYZa824wOTqNjdSRi9v6Nt5ZCj3WL1jpKbi+BP1sw3g0Kr5VagkB1D8RjN8s
wPzbncGgBaawkCBnH3h73ITyqOVbWdOTzk6lVBWiE/DDyuySgyP+Jr2FtCJouDgu
2bk6umzPtnY4axuszhmjqBzDttnbieotZtvVfCkOm9ZcZJc8MZaM2b16VnvVmTmb
zssKTHB2QDUHXp0r6nSB5ayxMKmAFi7zIIuj6IDs0YGfLhCVBeYO5h41n3kwzwNy
+0fKrR6q0s5aLGySg3/azJQI84LGUyOIvbssoDwPnzR7EfGlMphrnmZGU0W+HwBl
7LZp9iMTV5ThxFEQeSeklrMw4AawBFSCgCmLrfTYEesxwCL6ewx8M6kIDEhsJOYS
mOgs9STnq2tYxMaeUXACxE9TpQmkyUodgpjnYDndA+FFXOrYhzSyvTv922U+e6dA
VpOScJmvOwmHHEBx3INhrspvJkqg53FwTAQK8c1QMOaS7u2Olw9BgRF0DFh9JMGV
ACzClCSdO0ICuXMEUEclPcQkF1MLUCmf+A6VndTClbjrbPAEaXwe2ItaObl24llH
QgukTFUYPefT4zlke9lQKgaHiic0GR5FIQ5qz0o1rUi6e+wDeiWE05+l30outy+5
/W3yLOLh2SjAZycJ9EXUxXNvpTt4FFoMAu0+qlgl/kC4dEmYjRbUd3EiYYFBVJpS
th3CVOeVjbQcrG+94eDTLDyZ5yviYEPPLoSLj66h6K3AmJRCnYPM7SyGXwI7vq7v
Nm/KZWZ2xJCPNhmH052FVQlFphu1aLuKk2Rd7FU+lTsaFtA9XRWPr9LXFB+E/RCT
FqdMFh1oIGNUoc/rpq74En2cOHWptlJNjtSgJgQ3R2nHk1+uNYT8CgjtMPYt0RgP
wEU3WSMO3hfkyPBQnDxcNWsnbBm5EvwmZtuFgh7VCW9gxbWhR2YQ5fl0zxLsi9TT
EF/HhqfhWXNtTM5BtdRITF9pPU1ciLEHWdqmiH2WPuYkeJAUlHVGdi2QGHt5JGVt
wnXbADJGk5qAPyb8CE6B/vj/HR2XRRDvOuYSrzICBiqQAGCi9gmPay+QufeUWCbB
/k0vKeILck6COGaGSns+l3limcqoIV+bxz3oo+P3KyY+Fv59CYnuB0+zw1+W2bRp
QhAx86FvZ7c1CvoLkJ3y/0XmCzIDH+V4YmJnyu+GitjDzuw4786UC2V5ok0R0Flz
v4zvlzkRc37BejLm3BOW15TXEEA6hHcGheA5kh43NHLaVzXZ6AcGaxwDtZTPpnTa
yO9rcN2Iq5864tsNxFuJ1nzYXE1j3pkPADIeSCVAel74wsLkp0+4j228LDZcy9/u
YtUxyDK/FC5VF+jsDDdIPpKdMVTvDdvzQspvErConoxpNP6AJk1h5OnLRSqqHVTY
dQgoBdOBrEiTbesNvTdwlXzAYJQTdpgq48U+fOMUGEynB2W9v8Ud89E4i7Db/Tpb
7XDHGNT2bd66xM7PLIjTAPmAOmrznJfs15rn3/upUw5/83QUuHno/a/ULdrekTQ5
vQy6y68GSJOu2BJc+6NdPkg+RKEMOFGuXGybYLMgeEzJIyiRpxXGsXl9yvlNxpda
QWMy00ki3DhneyVG1XAj0uDpMAyAGIwixFVNztc9AdrhlGNChk71TOPGkEbTov7q
hPRdDAJB+XCSYfUMcpC1PoI5yljxnt0DIavc9QukxGmij+yh0+cWICUSRH8ESzUV
8xsrwZTchTgZ42FpUpVkXUZ0+NNujVjHNGK59QTJLA6l80rSaVKTOjNgg1ckjTFc
JkHngP6S2NyPtBNwiO6Lzx0udBusHnSGfdq+nKaqJxRPoxF6zhWee6Gor+65OHM9
2sjPcfPEXbtDWpsiiX/F2BVYNKvRy8LE8AaHwuiTJCfizIJV/oeGUeTTNXFrHPTj
OwHAhC8DzZIIz1zO8GOAPxDqEwrC3XXmnndgLzeQ20/k6lacr7eYb/NWUMLfbfbn
Wl7ihp62h1W/rTIr3nDuWd1ZIOjTgZtNkeyKTLeI5ux0Sb0mG6XpB+OHkZqMYrwK
I2GxjxnuwDX3217AbCH3bh3IfCGo1Mx1kO9zh6zSfj1E7jRzJ+XlAxos+J+EeTF3
qr54OdSMHo/L/gqCRevoZJcUHBRqOIeidKkOHLy1msYTRXmzYv9DgDGMDC9rsR9W
MQhIVTxPRH1fyH/o55BN8d+u/ziTn/Gp/v2QcArQMiH4kbZDcfJj2PQlD6j5KxJA
1wxqo15J2I7WtqkpykPROwFpuM1Q9EbVLFTxuMQ7Dzju+pkXNSGL4elCDZimqmh9
45rl/14kTIDTD/BH5iGRj4Ka/07ntaRVh2P+qeMfdYQEUhMTYaonRXDrSyaZ0rWS
dBgK9gVyBwREqUP/Ytnu++FQNzQgnXM530cVR9Atu0wLXccVLiIUMSaLjgkyk4Fz
Cfij8mrWdva7Fw7kTcfSUSMHYRi7/XRL5CWVoWH90fK1QjPR9kyraIJpiGbTkH+1
ES9ut9UeDEMGs70fkpYDiI8Z0DK+XWKg0I0HnLXA8OU09UYmU0oBt2EorN3ugQ9o
gydyhz99ItNYsFkhW9lb5wl4nVl85zpXH3qI06A4kzBLk+BkGVeIjmJkQvSY8jrw
rAKCGlB2XK9O1DF9Nm8AydUJq4lyi+5n5KgmEztJ817LElNYLDJmUkHPPAyEJ5XH
S/6bodJ0M5ejWqGDt4jiCrxOmEZTtv+xFyAsxpR0HsxZYTQjwq5rffQy21ehBuf7
NqAV1s+I2pO51IT+soSK+gGCHtXuqEnK0T0uTMkHoZd8toa8PIY0/CddeE1o2WWw
b2K5WitOPkH7xMbzOCqAVGKA8Wm8brKpawrLS921sRNj0I1upq23oyjBnz6ymNuY
1De2P4dhItCPdxOzfSHqO1xEOj3SnUWK5TIEeKh9/3bGSZlJDeQpqREQzajwBq4g
R8RAgTMf8DCT4DYCOp9WRZvL8LPmDgC9dzjLttu3JYv5n7EnGxMeAkw51GVspSxb
q5OzmROknuAx5hv1UBmjyBRHj2470QgzIvFV0kSBoJOxL/RImlNE8Lu7DCuBgJSY
uDlt5qHGfaALXgrW6wNzOLAjrtF4Pfq7pwRTnfwySkCMB/pj9La/SfRkTpzvt6nB
S0zqm0WfR3G3r/J6pAK6Xi7EPAfEmdWmWJ2O5oj6M9t21FV/GBTa2KqmKnM2r5hI
xkUFU7X5arsWyDpyhMzbb1y9Ag5jIvBYmwILJF0LMgxHCa7hgiL4Qm5G8f8YrX5M
5aABBcxT3Z7Z0Jg1hpJpP4DObilgaJnK26VNyUksGsTS2TJ9b1MYhYMhOJf3IFA/
GWOjfKFLICeYpM4lBcmhsMeErCRavBMs9SMqWucLmubHBSpKwyWE1IIK7ilHv9fW
pGywliUjIeIUStuph6buwT5wVfMpaoZnqGRiCX+T8PJCBDU7SFc5fQF8EUpu9ZOO
Te1+BhikPPqJsS8+oIgOI4f5jARbTGbzErzvINMhJ+wa4NrnYUcyFYouFppN0pOF
7bD9UpJlXNTWQ/s5vtdboRkZyfMFZMz3qOrJ89Ne+DJYlcgCQSrisHq8sXDp19DW
eY4Rp6cyF8047U1EMG97YaMStEXEhzvnZwlIEUNMoTdGrlQ2PGOWRx7EXrdkd+pK
2g5890w7LcpwXn4EV94zTA5LIMo+TaNI5S2H9AYt4oeWgKU+Yup37/JkeLsUnzUF
/MpNtpe2xanDBIkb5C8aoQpgBO1CWLshhHHqX99duKtTllZ9uLaDpWNrLX2N/lyk
Tf61PNk776mqj2/CQQAG3pSWsLmaZovdafjFsYq7U5KpKT4RSYLtX9kdp54BZ9qG
fZrTTCqUXQve6zXaJ15IkLFE7XAoQ5nm+qhaFxW2Qq44+vwy6pvCRbaUjjR+naQ4
mMhH6TWB4Ug5QyemhEqd7eJy5gdCle0lWPeFWtBg92a0WtSRSJrUbzyc/naseLoV
GR1Nvj1LBrw/zlgJ7UAUXHG9GjbDxyzwkU/3X8NOhgpVE/s4C6xqocAV0d8DHBIO
DBN5FnDcsPFXbNOq5Ou0GxNsj7zB9t2iyZBCZwvQVaZPyamn3IVIMXWjnIwWvFTt
DMS0dsa9wmTKoBQPTIWXX7mECjEPQB4bNVVIuX3JckbDQKEdfYZrGAQHnPDXln5S
xhVGNJpNfgoueVbSOKRQzGOU/zQtstRrzEx8ASERh8fbqQ11xRHUqEoTsELGqRqm
8o1gWJHWyEuzjpeaXMBpYUJoRjmIOE4VZHnp0qfY7iwn/LoSOY1RlcIx0RDW9cyx
ufd1wnDqCJUGhY5Ioi9WzZxXV3RIOL1DkudlgzcEJu9b3qVoySVspPEJeu7Y6nlX
pHpNl5nVxrWroZQ4Cby43E3fDjenkX8vRIP7L8gZz02uHnO5lucvgMvKJNuvPrY9
Y/kImvPCznlB/NF9afnK/GQk20RWxlSIrttXZV8A1kUvHboToNXfTMvSiH7Dq0UR
KJfzvqq+PXcqGs4BE+7t/tnxLd1fmg6ftmkoPke7TxV2/ttfOwG1XMxvheqImsDo
SOujTeUzMKtFYqMbaeA1oswsQQqLVbjgNg6i6bJuHvg91Yfu7qx2NV9AgD8ftjpB
VpKFA/4gL7h15i246v1/189z92We+h3xInD9PoeUHNNFKyKaFtnLrLhHCDmZFDPH
JmXbDfpQxaVlN1UToHi47pM/zafQJCKv52+YEGOzDI5uyK0by1quy2gCcpNW+4r3
muCljZ8ChYFyP5TulxMK9hRYHkYceGXdoUt1WYF1pFroeNsYkDCvHNAN3jgBQqeJ
W+bznWNriNvvr9I4JY7RLr2x4O1Uz1FA/bO+NjLCtUd2jyCJWgVaO7kH5iiyTtcr
QgSqhPN/7ntAu7uhG66BTanVGNahrvcLcb3mpgPKbmCPidI4C94Zaep3zEaegiad
iS0NCIMjSFvzmpAE/9Y2PDEkl3Co7L+nAYxPhttP90AX1kihW2BDjezfsHUgAZ9w
J0nDNpB+MF7rVnR+Abq0n0XV4oHgGpEcF0GrCie44fNTavKw8/cG7k9kp3nn2+/y
cO8h9H1ZPwXmkcFF9nG0B/vErSbgembugtuifm2rQP7roOfNuRTPaHZ8uHxIoYlq
66B3w12d+diMACvNDV5MKmHbhDKx2tt0SCWZxQyOzfnGmybEtBjv/sWbbwbydl3f
Wj71+Fj/uSueUEdsOskWY6ZRhVwhXSO/5F7oO6wq273DzPdcPYY4JxhYE/UOHyQR
930nrJbmTOUdkcUrhKf8Drkgk5N2EUp28v4ATyx5iEgzkT/sq0A7MLbYH3c1CEVt
hbjtWFx04VfTsDDG1KPa3+1tMzJ5cRHEGLfxotsLwcJBK43h56S26h5Aago27jKA
NkBSLUN9PvE5ic47AruHwEpUam3LKDrOBHYxrPFLpcVwrbiOsjqtggdKOhaCCg98
AO2oPC7lIT6xgAJT092eZrFOsOaUsUJlH22PxkrBH6dEPnT3OOFXjZoO5EiwT52A
12v3JWW3QWR/mTdeTQq95AitUJTGgSEfEbXiuGVLsS3z5NTZ6sBI9dWJYYHTlOeu
BNOQoBcRVnuc0vVUj8ZE+ZQG28jkv9rg0WQxbYtaUvF5hJwhtyBPWb3KX3rl0Zqp
Ea0RpGI52BZzTuIvqgkVB3TTrII8lqpf+elKZHW4ciipfe+0JvevbdTt8fj2U6st
4i8vzkmZ1LPwnY5nRvw5FjbiAY9768YrLdildgWuJlQOWOeTqL9Ejp2zZmnqjZMn
pnabZd6cYvSwuovp6eFQBLnDJ1y0DAYIWzFd5etd8vCraf2v0JTxgWzooeFlSisW
mFIrDv6ZZVnM74Mx+hAQUPWH+ih+mWcqaI2JuZOh6PtLaOqEHEI3nCW5P2wSYUnE
4Uu6n38XBjxXVwKRXC5PUGop5rhBZVVhL/SmgdmLtSvHHCZhYSSKo+rBkTguGLqR
aQHtqzOYlAIT088yxAeyEE0AgtGQVlX/Hg7c+ajZMGW0TVAR7KGlnQJ0xZu2y44I
TnqTuUEKOjNSA5KrefkeKKbcUXzVBjjPfQh5y/aqDom8463w4KkMyVjr58904HEP
nP9ONJ0ld6mZCPBFTt2AH0nG7lQ2PL0eIKutsZNOmYuT2yoq8z2kOvseiXecsjLQ
ufPSoV6ZeIELZlcEcGnvZsiFPgtut24V3YzMkXj1HexCcDBQpfEGuU363ZqepTJ4
jZoksrDzm90NfdfNWtKcT6mP/t6nCRvvvI7FAw6zURbiVebHdguA9Sa4xwJcWaE6
qmMI/ebksMAZ30xH67puMhMZRDt8rQE0vq/27K9OIjRDh6NjGB4zTSpa9k/9O3rD
JkpkbSO76vwPASR6zT6lLXEcoUDA3iml7hCVwkmOhLypOeixsRkMVhTkRUWWsR0E
CP+uTOzTA9abD8MgTF2sARvD7fmKky5BcACAQdUkn8FNiFowEov+UfvhsdTZsUio
eDtF3ZnEjsvCUc0wpj8qe/CTU+xTa2oy40x+AeaMblBCwpObxGeG5+kanZAQNwgi
Ur05eUFnD45GVUfqF5rmv5XGeV9/QR/RYbd4A0DoYxsoP40Owm6o6UHdwxTb1LWL
72QLnldX9TPrIEl/N1L/fsUGZGxIxp7U2clf8/VqaJ5nyGAkuIiIGuY7au3W+Ssd
DGstDMJbbFa2zwAmqzBXRV+b8ZEwlC9eUTEg5Qm/rDw38KI3pKn9Imv28XMiLFp/
qPKXch9+4Hxyh03cZ4PWeh3kZZ0Vn5DHszCBOS6RIMxA+1FyiBvn/5rPXd07+GSE
f5Zz7L32oGNvEpje69maB7Ca3U4Eu6cDNwapaS5s4nNHKzAN33+seg934EDXSuz9
NmCMiLPdL/D+w37jPTL9OTGZTteR2VTGv2/b33ZGviyGmEpNc9ETGKQMrIJh8mwh
DGogeftTEY/Itx7sO5SzKYy5Gi/9fa+0LP3sSkCqXxDzJ6CA71Vm/v3Qxgpaq/fR
mCPXf8ccHylijpU75BXjxc1WERQL8rWuK3hyFbdk8Ty64h5slfDYApBMcdY45Gzg
0hJCTqWh/IPOzGD7VisVEftnULPgXRph+jPgSmLWF7P+zlM3flHA8s5yLaPfc9YC
kL2vZjqJ/4q/YVH6IlkNWIwVDB8V4wNzSIPu8d9QcZHr1rPcKP7SwL0oYkSf2lYG
8QnRwfs1PVL/zMm8VadPlgFamwna80m3iNUibEUR92tTWODE6BlEQebEUowjEYTP
CWmt3VJkmIfEeZeP2FP3CXto/orvHVCOAutWKtFJU5iz7zeLwemfv95QMPT7QvIp
SQjKtK9LW9cyPt6b9sipHh5UOKIR3zeOgtfKc+k5j2L1KdrqDHBh4ypRfIm8zeGW
LvbAXgi+IKXBXoSD7+a44nwxxoO65rCJkHFemMWyYxeR1pWiU3MNhWcG0oPg19DO
JRaQrxlCxN3v+Hh61RA/9aENxkpBO1HL4/xbIH0W4KZ8p2bEcXDT5ee3WYvALqhP
Yd5tuLqtowcdn9lSvtNaxCKqWbCL1LUYHRwB5VN2CqhBsR9lJevtFDBeujDv4pUe
17nRLbEIv7dSyCVxm89nZAcPVkM8taX/ezZ9KEcvIOastRFQTqFxz6VC4Be6B1h3
GDaXaNoY2QOAqNzf+V69Z4MobmsHWrGQ+TVUqsa8HdeQHuN3CiZg/h7tD/JL0IzK
Lc3BCnSxaxR8ovoHrqUJuFkDYbmDxn671ef6JWyxT2W96GSJmKm+vPxS1rP5CQs+
F9KBKrtqYIxVTz7kfybFK2e7MBL6G6x62MceMuV2Hu0IReVmZQORdE5g4EcPnEnC
ZEuaEjTV8dShToDlSpsiuTuS0oa00ZGIq5IJ62lpkSce2IXD0jHdAPVW3WVICfaf
HFXSRKGXjvsGCwR05URLexCBF4ecdAYhrdTQVUYGBwgmAN3c1tt+/j4CE3SP8Jm2
7jdj89jcCDgYbTdMm/0F5XI+fn2XCa5kb8zQxj923OzCZL+PdPHkRnH/8fczQlTR
0pvMWCN0TQhOt+7UL26t3pdf7r1ZIqyPo72rAivtF/MPyrn19yFQlc3daoPNzYdg
o6NmOw2TLQIe+dqyh62eslAzBeB3JX7ms10OoHh2YPvJOwL7mSCR+VCQGsTW4DuY
/dGm2Kob2fOo8XE0bX50RNOOKvKDjzv2bARycUw6Iyfn8+OMcpa5TYjvLFjbMkBw
dGIhnM83LYxMzjEhdmyQMBn1CfheOwPe8Wmo49qJXeZHRX6dVSnd6JR+5ozaI59r
8ag71qd6B4JnoXps6hKW2U0rfYDIBspeqG5QR9/CCL+773YzZ576A2dyjUvOP+Gz
3oXUrlG+80/fUQUiP/PrMewY/0EZM8eHLK6dOuB5+RyeGeO5ndflbRiKBsLGBDMA
g8Og1rJpdhauPtz9DItjPXFZ8KC/rQ5CdlOveCaMTlPNUEvbijDOBkiO57XOhFHJ
GNrzEQ+/jntSVijbbxGCZkEbaBNTKpgSxK+XCXZR38F9UoF3vfvES7vKIV9Ssb9W
oPiJ7/Fi5q9TEM/HUE1AbXGNl7oX11azvfv9PFPbR8ew2MYK0iAoOz7ecc+CIBoN
llRE03sKISNBkmfgMSUD9l1jKp3ZDLQdrPnURT1CUX1YTaY5ay6RpTWIICn57rc6
QuG+mKCL/duZ3i+4kVnWdg4tODzzrS18nLRMBlH233r8Chu4h94gxDWhChQ2i7lS
KFrn979dCIbH0JkRMngkmoMauaRexCZuazBTJ0RWuwpZkdkaObkC2waSNjiVtJdP
/fdUasDEPpPwUymfxgyB4RMiNzhnkf8kkJdDKnUrgIP9u51Gi9gH8tC1pC3+Zh8a
WumF4WqcwrIw2TZmgGW3iJNIFYFx8tpzPZ0JF/PWYov+EzsQXJlR/ZFasR6wYGUW
1+bNlrbSmPu9ZPGSB0qE9iCZgiKqfp/rxFFU/a3CrNPUVFx0XPwMbI1XrXp1/twG
DoyjdfLUAWeTt/YcEoZP8SyOuT4QS6CTtmaCmW9zKCnZQ8tGwKAMclqNxjt/Yrwa
az95Aa+ASbR3EZqBZB8cPcA7F9qFqLGYpbw473NxE+dDSztswRJDeWfPv7JpActX
wKZHtY3USNFXh6bQxpmdACKsGKSyYuHSVRmwiOBHlG0nr3UTyEDHyucwh50tzl4r
bJaYtmofmyABpTBtuuX08pdNoDSaxwTsQ6h/v9CkraEGyVn5d2zx6440h8s5t1Ni
7qcspsULa5cP3RcojqBljnhRAFPR0CoYa59n+0YemOvgg8PsosWoH2dAbImYGqnv
p4Sb7x55G4Fd/Sh0lcr2OMLqdLeKvLgAr79dXggp34Qw4oQch6Eq6viHm0BfNnl1
azo+Fwhmwdvw3FRjofhVxiLJnosrPONGksJJop2JFvEMMN2HI20ZslZ6sAMXjT9j
O5RVNa3PGHqGcASCXRLSUeLnZNtv4Q1e0t2z4rVUp1Px1Z0LJmE2C9RrQmynLUHx
NOD8Zl7j1i+u9uIVMe7hr93H7JXAi3mIaRyJZCjsJPYW33kq4J5nZrLcwQySGCFO
blcL88bgXBCwKNzHo27SKhJRrj3buQ36vkge5abEo42zGo82nIMx+CzVAF3GDhpI
AWBjpAl2284OlPBUJeMWbGXUvfSDfqUrIwTm0Ho/Fpn560r+PxSzPXdRToxDrbZO
heNBAY7dSNmEmFuiTTO/EBvWHD/ZCjskn8BZklxJqejQnZjLqBC6bh/u4HLG5y9O
rP9geU41e/DfGKzNqHc+q5NnRZt/avL+tze0RncEkF1LRjRAtOqUrHx290HI2aR2
6/pKuFCNMzJ2WIvrHIcyiHKDIr7xH9ZgSwyshazhmlbhTT4rX5i0wTEc21UcQgia
46iDtxbzjycNMYXXXRGnSkjfFtDMMg3HYI9bieenAXlFTaRc3mx/epkLggI+w6M5
ykXQnNIRlocuB2660WlNEb5TsG7T0PEOseGjs3+swJUKb6u6skqp90NX0MY3a7Wm
vxszinyyaC49nCOaAa531T6uKGcGk/yA58MUzsMar+7ZbHEYQqrAZC172ocI0KwB
JkI66/0CdWCtrvyI+tSo7Q4faRXZHWWxiZAaLfpPd2Y1hCJ4rNZCPQaNbQelHeCh
8INg05CQWOZs/Th2hxCKasUBtSRVsGJfMD+AhppvJOa3M+RZpKwllUC0wf1+hdN4
7kOGYkcid1OItHLptjr9nY+8dmu1zLfu97I/JLabpbOszMunRdONpp6iL+rAKhG7
ox++QTdr7hzbQqOu18HUUDyd+7kXyMbvLH7oi8TlxM2L201aoLjkMEBT0PZL+f7p
69lMLWbVbPb+cDZnQEUrfpw8kjGXSREbpSXRBD3jZ2eeQT4yXlWkMxXKAEHT3HOL
aler+2OT9IaIGWa696avnwFaqj0hzKkFUHQRbA93LJBDTBINoNiG0yMSi6Q9FWiF
lhIgtQF5RgdorSJvpl0N+nDEYwMbZlV1Mnj7xto9nrWrKWl4kNzTW92i6dLZW9pW
6k9l5hhRlvSS1n6LyaqIMNOvaQj5IYJ8RmbXH+t2oT+UWouXB33KHS3ogomFx1RF
FcryVnbzAE70CGh6LrEKc93fRXGdknAxUI3yOh3f68tFCE1pd1C2yVuhKEb4E2hO
UxTs7KU8rpwYGih7g+kx7F+EogTHq04m5azhMuTqe4n1D5wAdZd840R1v3F8Ym7b
OFWj3yWlU90Wl8+ZzrWRvrh+v7gEc1SwWLc1el2EyztQKk1wX7luyOIXFcLQIvnM
zT/hV28UdFKOKwaeb+iwTozIy7aRDJ8od3WpJgWPFPjcEfCyk1lkjTa1zScWKGBv
i3XmzsBy09OPWD8WjkeBSkp2FAdIS4GbgTgpRtUXrR6os2sCvZDYwWmhx4ShEY/8
0JBttANAE6Z4laXmUDgJXUwr2tsXCX6l73+phDlQnLCWxBkSJQ9srhvdDomV/TE4
PVhdEJhutkXNdXu91WyQmzC2i5eGUW9GIovQDRQCslyu66Bv6EohIc86n2qKIOzn
wFk+KiCFdPDgTC9FuADCMf2y6nkCRs514MkvvuC/kgJ3TDKiee8hbpf8Pf/z2TWJ
/4dtRjIcpD1g5s7bTe/5vpp/gH/CKbu9RMcTYAtGp3cxi6XAIZKexMygekyK9oqk
KcEsd61alH+kMTOoGV3GbPnys5G5oFXOQGSU1pm/I4yq83m3setT0nRfb48a2yDT
thPVRoapbSZ2yzW7ffYYAzLKKNJPNmD6r8EYrkO4bKkO82Gn4VDvA2qoPKqvnfap
Tw1n+uyNJwuxDmIg/QrRKwSMAg0J/DIWMXSUA/78NM1hnI8OvsgRwW44pZNP51UN
O4LLFjwl4MBbzwk46NOpplRnH6PQ9QacC9jnSUaOZjpidx39+ior5Johkd0PCVtv
dOmTocUQPHDl4Vtacej7wJA+QuUFn18FcpMcQePa2R7hWYJnuPTm67t+xY8DRXKE
+z1a5GIDLXIBlH8KjDhumpu6Z6fJkVecw8NCytoCNt1TRUel7u4ncJOmgaEB/46q
yCw5BpSC2TGLobjTWYc+4SN2geIxmwVmn7BGK4dBPY3ddcyfHCxGPw7oQfT9pnMl
JRjA5B7naFfWS2nZOevXK3gmp9tI9+jdgACK+F1Sy0l6KVnmBVukMTdZEpNSx7nu
6CVG1GfWBlVKotY4SXyCCq3RaAFNqvI9yNBDVMnv+sDicRWlgypjkonecMsefdOn
f6vX/hALUXMJL0FmH8qjy0CA7wfgUOneUsJsj1ZS4fq9BqqPwK8wu9Ok8Lb3I+fq
xtPbaT4+ctkplDLPd6pv030MvmdL1XFA8pqYRSsAW3vlfzHE0xAskjbp8cHCHSWR
kPrBKuV+e13Bd1Eqf2atn7kg+/e7Nl/XC+3q9Miw2IPBx4PXKuZEKqAPtMe/N2nm
uW4CpdNTgC9j76xfv/WGuzeZ1LpAi6RIUCEY6FYkErUV70Ttb6epQ4J31zCWvfiq
rzCH6PC9OLcoL6IBMxi5IEDYNPnXmJ1IP1Mp+D4kxwu682VDE3gSxqWxtw2n6H0I
ByMNHjKaEEE9lzhxJpQazwjzGktofgk2/LIVhrWEh/c/nkGMg3F/UsjOiusBE6l8
4TncHoVDV+fRNGaV/Jv2fsDV0DQ4rku0D/T1r6i/2EGnm6ZF7eykxlBbgdM6qfiq
PL+xdSoHstSCH2BLNIpOV558lBUxA+ZiWccSVHSCjTE9LqPnwOyDFjkYGcdGaPW3
f78E4wrP25X0mAAow/4VrN9mwMSmhQjcZS/A0ZlRRmNDdXC+y6ROVZ/ArnT5grY6
MQWBlEiv+98LIyDq0P95B9VNfMv7OktE+tNLHRv4/L+snA6LG6jfMZy8kcY0v0lP
d2sKlUSN8P6amX9Jdy0fTANzJe8dMbYjcRNJZ8//oj3uG+2MV/xz0KtKlwEyQqxr
AcxkvTUhUjxyEczMLcRILfUvEqgXuOwD6r+joPhsVwIAuFh/QZT8aWAuPpYHHmVe
ZjxpznrFrm54XNM43quz6earZUW+XF1IjXGPGDzhIYkA/PKqSy0LTDyp7V2xJQsW
KsMlMDvePK4nqgKcatENKcX5ea4dZtUGAQqoJtGWdAtXq6cUQ/j7s496U7AI1H34
B2MMNyEj8JYnx+xoGGLOc/Hz9vfxH1FgNnkeEeHbJhe76q+TCBzQEHrm6JKTNvU7
R5EGT3MOya/tkE5xw7l0GkjixrUboc7RViqjV5GyeBuBpn+PmzjH+GCHwis+ZhWV
7bkroXeltw6rzmIWEebB6rPK8irmC8Ptn0lA9WjqOMSPp06rw/Y4u2jVSNuZ6eGL
zdGfytOtE6VQsPdIcXVVtU5wRqwXd4MszwC7eLfFY4kP5GfylLxtbYHW7VJ5phCR
uNbdqr06brv3bj6ZCpZJGdU/KItE/jIGnjB2PzYZlbG7ClU4C10ej//S74pAf+g5
J1sNQpAIpK1twoCzJED9GJnlndIGUEMJkenA7ahz2IhfQNdod85elYbCl57ozx5y
jRIoEbrEDWI2g1j3cWD2CYagAiApMHqHwF21HBgWm3TOcb6tQoDWlVagnuDxDSlS
Tvf9U2y28FH67JXWREEoMCALqR63wWl1LuYQHRld9RWQVRSzg4gLS7gvg0u6JUI/
FxHNTin20YFyOKy9SXKGYnirZ1SE7IBajj17JSoRcQx2Qf18n5930PpdDeDt45J8
3guY8uK6aDsSSpQrJrtV/PUvyF+fZb+j70kwTHBC2IzF23JWOxh0dvgc7lwzV8IK
stJAzZiH9oLQr5MzKgcEVEI3b0z3+RmcY59iua86XR5QHkaKb+c0kUruM9F4Rkyz
IxnAhNE86/xN/rbt/2SxUWiELDrB6tHZ6GgUWp7juaLplwaaFszbmqdbbPYl8RMZ
JntdHtoaVtic9avCqgwxuVxch8gtPDgSlnoBM5TZ4BeonxeUaGEv+bXO9mdrZp15
vLjVXY1Cy6ucQpOt1iPruVdElhZibzwkiejEluH31bXMzeAzXNv8e0N6LOjl/VCM
3Iktl64ieCuoGOjRWy71hTUcRmV5x2A3odGE0PWMXcHnh+eoPjRxyI66si6jNYlr
G4259ReXIEL94CkEvJvSmIPUKoytP+91LOcpOE3vPhHROQ7khSZ3TVDEjDUAA2hc
bdsZgymAQnx4P8Nv2r2f3BDZIf6nPGDZ57EknfeXuBFq12XHEzzMCOwlycSOTfrO
2mpznh+vua9qlDHbUZmSQBbPHlIcI/Ag081S5fYCFNyY5vNKA39nIiC8Dm35wkre
ppgUm67uhJnzneqXd8d9GbrRxsxbaQQZsWlZr4xaCnz1kEGjwZLbdD7PD669iQfd
mqWp8VFkAF09UD+3EaOeSoa4RlNVDKGvnGIp8BQx/FaL3dyLY8tsOUrlO60BV7xw
2IOc/+3f5iNwgWJOObK7/cJOOpc/S1R6ZKlYlUpLfUifxT4jZ2Jg+spseAfG5zow
kKCw1x28Kvwdd10RK2S7FOyqIKScDo7Fln8SF4vwYe67i37c8KK1MdWn7F5I7Vh/
8xnLXenW/6JvSMDDYbrjcoiARsYzfb+IZXG8KlK/+KD/zh3i7hwdZz6DR2DKWihC
i1wAbSrgJm7the1ppI5QRkmeoMeQwbfXotYKpbwln9cBj4EfMuTT7B2QCeMtk7Us
IIX7RT0Ssk3pTFeckGwLtbK4Avj3y0KT1sbprutNQBpZjpV3WMXiRn2bB73+56K8
0hssWGGwHQTK1t66SQJigvRF/MeS/p6h0L6vnsQHkHbwzS+I4QGJY3oeJFU6pfrY
R+t3FbRSgsCp/ps2vX4iYbuMQarqG5jhyxhThXdVd7GKWY6OCcb+biLfeHd4zpY+
qlmbZ8gtN2dF1GFGhn56SeQUuobb3zo17z4pg8tSWtJKj7U3YJl7EbM19R+Xvi8i
x/YGyPw6UJaxLjkbJaKIFtnNu9foBzjSY/B2wiRpzTopiQQnbYY07lAyxZZ41v6O
WUzDOYY2akGlnV3d8P2ExuywhZntZcw21ltRAvTuDtVjejC8mF48iVqjH3VjAELH
WWSL19SfHHJuYOnjmzlvIq0PNcqUxnvzsiDszi3QUQp4APFTwv2uf6wSgzCVIAfH
g3llUGOpAGShmKpnsUr3CegEpCLoQpEgMJeHMJjV6lwJ/kJjnPp4DPADb3NICsf3
OrSdkNJ160ELYlot6KJw3sxGo5CbNzSXLBbBgmihqq/Sxh+RjYDnyTIv93wCy0QY
OMqV0IPCiX2s/zEKq1PEyeaQ/WZm0M6V1SKNycvKSItdb0Ue0jEhpVjOkaaeZrKL
5RHCiO7X10Vu84afRKVUt34ys4+V07OecohhHlmW3TAsMh4Coj1sipk/wUqN0tc6
XuhJn4OtX3nizoKrxb4/5nYggdQds9QYK/NZBWh7jkU9eH39BXzUA0rrz7qYyuD1
ZdLfrK4U7CbH+aFrexxJF9R6NBxL4FvWJ2L8HsfJrCjZb7yY21Z3XgHioFGvtL5f
N0AFI8uZw89Xil4pE74BGrg0JwrZJl9UNGQ0bhVad7iftqlOv/usSC/rvMecgsYl
9Id7/ifzCbRorZb36lFcd3+MmTtJIUkHWjABsiiO4TSTxVZUUVTimHf7Vvrfyn6/
mjI5MaT97kshLWf/8R/kOUTaPW8/6bhgjONjNFAZ92LTwJnB1cDIYjXYqyGfWSXu
kzQosWo0tGir9CuH17S55HqEcV0wTVxg+JEJU8RAB8qNG3lKjMAOBOGhzKzHL68n
bFsiQmzUCm+Jak3YuN21oKaL6SBJgjunASJW8NXGpAHTQrrAjxbjIsaGmcVN2XAu
GrPxZx0OXpi3BEW7NtwZMMODWpyZ06LqsKbu5aYx1BFPe3FjNhHIRrfRrNPiu8Aa
FoGgJo8XGc8Yy+YLBWmZZTyaBlbX+Icrt2ZZ2sZn9E0X89ny5gGxLTTDOrBrMdN0
/HcLZ9WF/XW6yC6epVIUdVIr9E9bEZLlKeoiNZDMc2avzqur8ZmksMwVNVmBcmMY
Wue1kPnA5NNJJj+uQg7rB+F1my40BLjr+D9Nbqusr0bicZE6OqNvTvuQDz5DrwiC
0+v9pO6wSkQRydIRO4GkEE3qX5HrGKhpo00uDSbKfLBTL4HnULl8gnqi6N+pmljo
9owrE3TCvkyjhOu6MZyQ7LJd/945q67MxKAmyiCf9yo8ivqDlWcVEH9u2THv94Ag
aJU9ZOBBWHLm0WP7d7SWq0bl6/Q4xS5BWvw+gr9My71GCzpiD8X1+bKsqXXuZWyQ
5sLZyal9tuJeLTvsU5bUdXBJDYs9vOAkFsejvS75JGAdM/0Z8H8/lDxJ1Wx2TakV
8UShRpUxObvImMrEXhn46O6SZR6/WbdDMrJJkIAnKRUCS6X81rDPkGZl1Z2arvCh
kEa+zQ4KgaVVbh6nHfM9zbmjCpRhoaSnnV3k7KrabUgtCrsyobRuM7FCDw4uzw6N
a/hK+BlIjQfCtjxr6qZhi/qgX1bR0KqLXANlVJaK1r0R5ifvMyVGGPGlVT8F7Dx0
g77YrpW3TKxwrLldiqsQWRCTq6hSOUjCFW6BfBUlxXBcpH39Jag5HZDUDsHpx0He
HqIHnNbGduT4MMDSMUsN+P/kV+bst7UaJLPDtBr794QnP9OKEfkyyfQWGVBx0zFe
iCMt3RK7rUjUKW5IMiLL84heLL1FWua71uhjfUi3vIStmoQ1wbzjXS0kesUnQDfj
JMywFYNDuEuV/JBvp143pg==
`protect end_protected