`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 4416 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/9huKRhRMtvnNqb3Z+UU7TahEoHV+T8U3P3ufru7l1O
3DlgtZzb9QxCbOjthp9+wDkjygH0eUfDrEl1ovhZG61EK79YEzKeX4THB8tjhW8V
9yRc1WJVV4U5lQc6CykgYAhIo3xE5Njtidmsfz+wH1psOVC4erjZO7TGm7oV2br6
fjN8dJHTtyMKO+k+PmDuTD7cO+kJPw4aXANo2iaQmakdawQnDedaQX4Krhqibcxi
mCXBsqM+3ZuIDqT/xwcuwQnyQeVIwZx/xRrh8dx0bAWB79Vyspv32y7jLCAepAjq
BodFlt4IP//IMDtp4N9yZZ45ZNuUfD860jKgCatko4eMJ7BT6EIj8CcxfL9QzBhJ
qF0YPaxROm+Hw9oL0vtqpd7Yz66ouWy829PXYkpFIfImjyWECcJjjxDc3+YQEHWw
E0zlTb7xvtHbRlIMRD9AkynHsMMPWkenZJPuDdELEY/emq8sdFLF2jInMuTeE2kt
u4lWq+xRw10ybs38+ttZhADx2y6XUZmr126RWdVHZX0MZz2cVSSPkUo+UMLR+sQa
yHVryQsWck2RlZ/M9or/EA4jrMFxw/KJsc9BoqNR82DrlNDHPA8mAcYSu7oSVi7S
t9ZwLJvBNzCY2tfrOm/m8H98yphYVasgiafqoiJztpaZx2ufysirclD/joOn7+Ci
2BIYV4G/nLeaXrKLNXzO2ggAOAuTjmd8PTpZIWB8Uu0XY0ZA+KoVSoXOZUHnom1v
LGfv7I8xo2P001g/LDzYOiIcGVOPt7o8qDhrz3Q6RecrAfVZJ7oLSdEyI3mEASha
OushynJt7ffz+1tELsYTx0Y4f4hbQq5kF2TMePtN/+SgOACgJbNvxjliBflnAzUv
qGmzAXoiOEvPeQSRvzMPZcsx3oezXFQCh2XCjVYgrqQ8uu3o0nM5k/70t438l9n+
Wy8VNmrI8sArwvHvHwiFI8LmNssqvbxQMVpE9wX5Izh94mJcyoxgdTPLeOoGEFfO
kcifUvHPd8uag7uVmcNCY2O29YJopdwat0usih+s4fhNZwVBUz8+/z1tPDc4E0Tq
fAcOBfuKfSA8fFO+UwUzh5J/2Y9cj5ufmaAvOXneevIgNB4w45OJb5uxqd7i57TZ
t/cVzjqkDOkQLZlMyoEyEd8Ez9rGvXlKPbzTHjgLvhCSIRW0d2Nf2H60/tWgv8FE
2995DM0vZFo4wTyid+96jGyLhvqL9FeUzs2dBU0lU+3eboh3vFIf/U27OHy7jfVQ
NjZsOy74a2eUlsMjjZ/JQ9AAODLQqHt/uzNoK3Ymi/FakMsNioSzfzInGox3HymE
i9ouijDPeCg6ajpa7fzBx4kPq2kF4S5tUop13tdPQpnW4j/fFfaZOJcbMMsIQVT3
rcL+d5ltU95Sr+l5pcWU14BOR+3XSrJrt5gQj+XfXraHaER7ullaoMnTQQ17Gzeq
ycFwNa4TWky4tRK7MehqZ2p4ReJF/JQ+C0aI39U1RZiNNFXH86QbeK2fxzBd1SO1
YD9WmwRmyg7wP4/Jj0mYfu1ZyYkcDVAWLP9utAHVsG4zC5FNwVrTzgF/oPS8MD+l
dGuoTdy48PsPJkU6UdlKkdKUz8DI6Xz6oIyq/3kzfo8+NxwWk6QZZIqaYYYnEdsQ
34nKed5h9FP3jgYEoroVH7bV2KoVT9bEgIfJr/ifW4GlFInTbElus3kYXd/vUJtw
jX4Z2kak091LuB0059bjjgcQR4NbRlGm1L1Q93nfmM3tdOmEoeUFkRUgbjjquDSv
IhMwMzFjhH+gcZKQRC76zCLpwXFVGGvkEHzIH6bdUXy+s3wU+TqM2wKjOI9x967S
kHuv211vwkPQJ61W4cgLIeTCBJ3d6XzoctzKx0nx8CVhL65KNK9tvT6lTdDt5HxZ
j0zRs/TsxOZY2HzAYEY2Iu7Cpv7BoMnTOFwUQu2LwxeY2j8B26dJy8je8JKWA1ge
2g1ow13M1yD2r9c9ZXjB2MR2f9FclmeadJzkyefaDZyLh00y0pr6Eg/3/QFh+ozl
dLuiFNvVWyscLuLVZ9ZRLhYo5TSFhMtrOh2xnInMjm3YQkYHIUeMLEIC4g+DgWB/
q43X14RAvfNqaesEYO//f0aIY79lRAUXjS1zcZ2r+RsiWveRW2fxM5jdlZCJ5iiF
esSkwQYeInvvScGW5LV/O/56jUzmy/oXkC7SpzWkxVC/i+jvvPRYe9tgaVCpij28
op7ZqaVrLPAhzOClRbbcHaQRaDkRgv9yuAR6IsfV3vbu9TZDLeQ986Sd7oyhn6Tw
ls+eisTYX4IDukVx9ISydug58MbKIkbTB2pW5RT3JpmE6irQplKIZwUe5yFOr54r
919ayckHjDUndc+9QJrYpgfBA1JVao/SApOlOiik1ZxANkmBpiNYhdEWib5dx1zh
6UAYd6kiIq8hKcWVcDw0X4lMtCj1S0UgiOooRjong6hwJ1mIaELIv/mekzOCMu5L
eQORNGdFT2dg3MrgdA01dgOZYyU3jhmH2fs4b9iupQ2hwSwHvvk+xTC8LKaQwFPB
eqYY0DRWL/HGMf2JD69TZsnHWOBlEnmP9eB6lV3/AF41bgoLnKzovV/Jc/4mcwM5
MY30S3XjReAjBirjK8dWA5LV7B2u6Qa/UHWTeLhzKt7bkQf5O3mNDlV7SW1H2l34
WlTkhabEEwMFYLExwhzS9bcV5G17x/7Zv40XZvpPdsFWRMQMcbin64nFBLAHYPH4
vSgVZMOLYz/9JYdap/QAaVW6fwgmAsW1Srp73ibCeoYEDd1kCPXP/7qLPY2ManId
OOzpIOX4/szfrlM+eldyfVVCWch+/DD2PgvVy/Fcwu/AodUben1pEr6kgC+R+L2z
ZoBPTZhHI7iHXl5qiWOTVd91myWqvtJicEjo93HJ3ftkYy6GoDA3oL+ByZh34fIg
zQiNIIt6I4DsgV9A0jB07fbTz2rdr/kPcUjZSjvdHjp+bEAU08bon+hMhCsutuVX
gdfheT8s9mlfqmsdhlgFs6ylAmeF4C7Tslna7jTwgwzit9QWylyr8irARC28nH4m
FV0f4v0UNe5mPxJXzjym/aYQXUqHMLOB+sIfjRlqVdr1D/pWmoYaD0xVYitRQfVm
b4XBcnDtrwrgeEd03Ftk6djqE6B6MY1T4yjT1Mvb8oT885iMHcsp0O7LkPehHJRp
sF68VaDBrZpyRw59g6ZsMvJ6ySZkn5zBdbutmdUeXAPN7XrlbBsavr9KZNtRsKiG
w7/MWRsKD+Qi2GOmj+WKgVKSFyWLZ2EjYlxtu1HqeiRPSCUpFnMEBGW6lZ/jBBdk
FK1Sz7H+wDeXNiu3IGilhjW3dgMCn0J2qdFruFkSOzVr+7gNKaHVBXRpzdQLjk6V
+3OWbS81hh2pXrELj9I3g8k2i7Fwae7PVBKEEjuLK/Cksf4tHbBgdUcNtjTBKMHR
lRtgudc52/DeLoO15U/qOOxZs8TK576n780t6Hs+qbMuIZFfum3MtAMgnrdt8REs
qIDo1+MHiHpyeH0D5c19H9pRrd84GI0RzG7oAVtrs6bcIxtJ5g81bH62hKuiFm6G
6waKdQCq+lJQXjbmOgrryioKHLtsuKbW2vyZ0cDZw2zAwYSexxFnVMrlvzuTKs+Z
MdHNZjfYV67EqF/VHWGU2A85cVcAnmp3qupxcr++67L/w7v+z05QIuSWyub6wjsk
8hvBLwr+pnHOl5zBZmDY73W/Q+G8J0uLvRpiUr2C2h+k1WT7xIweGUMzj1V6Jd2+
zZMAeverMGauDRBLEYZ3shYLYtLqBiAofCPig7CSEOU5lpgG/ABsTZd/v0DGeGap
m+p15BmS8q4pFrcLCnRPWkexYBYciLdHpGLF4AAhUEmBJ4vuv8jyEgUKviJn5NP5
+AZM/N67LZdTQjCELANWCUeVJ5usK28eGarnqJcKMuLr7/05gq8ee1g+YIY8uBbo
0onKtLGov0ai9XsaA3uCHo2XcJfHRUtjT9Yzh6m3Gfnn0A21h4AL5MTZjlKbkDvS
SEJ/3oSMw6adT2j4/pboN+Px7I1YhxlHBCQmo5hGokeGwsxckGQl/W1uP4Vdgt29
c15s/vFRojSbtRfVSnHr0ZEtBxQk64zj4B8Z2epUL/QpxMvVmrETUnN7Wjf2ocUE
ZEZ4a0pgcU+Unj2MBW60jij5Flc5qjHJifC0bm0kbtczQpVA2QsU2wgTrFxpY4yJ
yZYZ4kA+3VetoWj4OzNiaks+ojIkHCE+HNTjvGacqHUbUh0oq5ndivdOovhUm9dq
7UWHNBi0en03wAZR3rwiU+p133iXaH99ZhXueOEyPKsGM84lNugS6KSdHnIP/N0f
z4QoTyIZFS9A4byJ4LGP6WtOfb6volcTbEjPj/rvnYgjxTklOAnq9G2cvAkBZzTF
etzw5JHhQW1PXB8oGaCFWFwaN/TaK2N0pmoS350cLUw9IzjXSKdjDF+mXOEzHJ/j
g73L3eO0kidSZ/KGMnpAlG++KlIwyfAmHuJDNaPSKvX8LI6jZ+n9PJOjkztyo3NZ
Bmc5VPMWgHaRJK+VgjwfEY2hloa1C1eWDNmR88Vj83qOoI6V5OANKUaV9+bGljbJ
97qkCHPubY+p6vw2IpjKkyyz9HOifTGX1B5+hzyf3hsJA739Vqr0TuoUi1PRDtPj
H4Hgo8r1tL8/VBIIEK9PqCfKjj6PbVebG3CJZzFu1BSuWc+Ghb9t3ubSnKKkr7wl
7SYXRzHQYydGBeoxV8A1Lw9j38mAkVDcxIH+L2IcKygPaE5SKo6TKU6bu9b2D9XF
tJXjuekEavz6/I1AC3YYKN6KL4kGzU5pH5k6YTzDzW6AGVT2rCBplzXfCVXa/aTw
OulI62dX0fd01zEFJg04RKwm18UMZSqoSAQA9VhHGNa0XrxaF1qWwUVAazXopWGg
D2JYZ/qu/7OA3xz/+u/ccscKl20OHWgHh2VhiU42DOTjrpebZEjRoboGszjVKyiP
OVFyp81XAJuZX8E6lyeuP8oz1rfQgBRehda6qjoMq69nKk4NKWUwY9lzQggmIiVq
Rm47N9o2Mu+QVv6TrJtd2FpsIcf9KhsuB64Mpa5tgRT6JB9ZndmbZryvidMe7A8a
uSoHe6AoIu0wffj6XGpj9FbEy/zmY47FYc+9gEDhXncUhBcHVzzB+hL3jkLpTowN
VZrPiLnG4C2d/Jd8INqnyX0WT7DlXi6WQ6SVlF1PnGpwuygZuz1qYRmVZcKUt5y3
lDxByu5kmrEf+Ug1RMK3laXtVgmWNPqflAW7nfRYe+MZIdQXC4bV7YYbCvnDEcEo
P5UZN0QOZ0JByAhbklTcdYieSQsauKPdT7vZCPz6Pafg/BL71cKnMYfHi3smJJdP
izkBT2KYsmpkOLaGDMwapWk/cOgMMAdWp8Vo5IjEnxlZIpmThxXCjIoNFqtti8Ns
/egy0h762FEayanWqOcF/pzu35f8o0a/VMgNKB/8YgGTu5RTk8I0P7RmI4dvJeQP
4q2CmWthh3GqRMK6PFw5ovYL5JjL1dfVnMzpLiv7XRNmF1nNZe3/KqsuDovD0Srk
U8uOQC/pW23Mey2C22gZ+qy5ug2FAMU55JnA5naMFrgO8PixuOJYnGWL8fDjS7BS
DXDHIO5SHx9/aS30rNhf2eMlZjcQOceieTiqFF68CE5b+dpJ15MVSvWhBBvLmZO6
E5Lh/q0gZWyBSiboLi100WaUIi8gjXb0m+KfVymY98gZSGWbshpGvbstxh7Pt8mp
4CTIrVQimiNVBhUfbqxp6hspwfwIwCd0m9YcokVVPSh9fZfAEsEhqIceakX9LfU1
CfLO0FWqgrDbnP1rYxjmpvaxiciQoZ3GqAFsyAEQ+/W1TG8JjuxDA/bU394AghqV
`protect end_protected