`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 2256 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/9huKRhRMtvnNqb3Z+UU7TahEoHV+T8U3P3ufru7l1O
3DlgtZzb9QxCbOjthp9+wDkjygH0eUfDrEl1ovhZG612Qz7yxVrQovfAANKeV/Vz
fBw0xvm8LiK4oKY9F0eFVMWhFZ+fGG3t1yC/fJsV8DBfGaMC05t6U190nVbJeT7M
I//+jb3iTU2XsoSwp61h/Bp6LMqrAi3lJgf5D/T6m6iLTYsTEWqaEyENsBuB9Df7
4sTXjExuiSEkUN0cycNrMh13VyKF0CJ1sWwGxzyb6ASR7A8yXuuiVTkWZUQXfot+
IQTtfr5d1/rO/q56tJ5Yj9v5ry1xmnKBvDboInd34gfWHKwit8O0wwjtuNQqT9Gl
1CqSLsfwXWpeByhEpBcewaT56j77pOWeHPH80W70uVcBPC03RFpdVVXy1gTqBLZC
++vWk6t9LwyGdambCrGhbVq7HLe5TdZk1FmgnrRdjL0zxDIkPbP9ljIRGAlJSNCq
GK7+U7eiR8F5acSdXiS/bDQe+xuvuXELtC5AxIBrARGIDQL42RYMK/E95vRYZ4L5
BPXWZtPPKeMaTk93aVaXMVCwdIe8qB1+J3YsVUDIVmDo+n44jmq3UUGSXrQyG7Ls
SUIoMxeMVo3HTh0c4Pxw+OlBF+d1aX9FmWTmMm7m2BkRis9zsLvyahKJsKQuxJrp
T2nIlnhZpAD8b/5QdCOg+AWDNqux0ua5npQT0Gva30tMDKSnmBsb9WLEAqwsZ11C
cw2isyfJGgSUIwK4zKgqjZ7uv+RO+9Ns6Ex5ZDbArs09TJGWqhT7MV3UL7KGPgu2
Nk/eIWpYWxgBXDnmisKwlBDhPv6tShgJY5qBzFWQNGaCK1sWU6NwPBUQEIFugBPb
m5B1kdslHs9FXlWuGt5LCUtZtFqH8RmbaMhW612XlYXSJtAKJ714mjqcQBPNWt5O
N8YKG3XDOz+8QAcvpg6ViITd0JYcZIsAVY9aWEnZcbBlxQLTK+C3jGG8aNiSskyh
T3xdwX7ml98PTQwSt3hycr0OLU+j9l1Wdklg3I238bqsSm3UlJXB01it94PzkZzG
FJ0bdf9muBHvyvnzhnI6apCwI3FHoarlgQXuO86pH0ff6+jjPLKDuGMsSZaR/1DE
VoTzbcnE+dyIwLUtbymL6aZVvEi4nvhbP7lfSodsVwr/FEbUdfb+R7xw0DJJVWur
rWeiuZppEiRJYc6Em0aECKQLJksMJN0JVbrQHYmX2l+dhcyEHiJAE76/pUtIQ76H
S5eboqwOIBYGMefccIbPn+jSk/pZMsafQWXwzoMsXoZXXY5e7xqKaijMAQK7DXqF
uoOCxHQp+aqxNf5SThtB/QEcTEAoW3JQ9yJ3TbVV9g2rtibUdnmFpdPyRTmBQKNZ
j2vwB85SiwnuNSymaXSw5llLYVSffT0Xbp6XaRHf1yO6uRmswI2aGjxU7Py3xZ9z
/YHD4rOgA9QM1w3b3F4fbl06wZ/O8Lu2coILvEpIaQ+djRj5yEe/Wi7rWHCl8hrf
gMe7iN+XzkOIe9r0c1mkJ2WaQe/H8p2d/WWZnviDhmRkd0Rq16ygvEBvMO7VeHEs
JfysWNW4GYdRM/f5hCIwuic0ujEEodisQUnki9XXrVkBQfjV1gkPaNCxNXLeQA/t
+9KFxoicdat006ZKX2iCcYCl1iGwhe4vAi8BCJ4F4Uxq18wWrQXl1vohATH3YxLj
qBocslCdsc2GQy/0aMFJ8BL0V9JLF1OrziluL1CLJZo/26gpRk3KPaiSUkfa/xkF
C0OWZmGbK6zvtfBqaA09+Zvcj3j5xKlr2e/MJZEY1XH/xG1kxycXaP5Qa0sqcq6U
44uLJzjy+Q+ysdDSO+0OFzXAezC03EOSX20YwjjhM+1xxkWbm3l9A7WE7uTO0YIe
VfzjfRT6ev1T8LvyRl1zR2TN6L7UjW5ky1HKGH8+elER/iFg3V9sziVFPI/MmNyw
GJzyTM+nPQUtMHb/PXs12oHWsbxMBr1/naXtRXseDb35x6AVpZih0gJspVhvh42s
vcYijUOMp8kvychr948P5tQIenyhIoppjCKL4bQPcIVxE/5yxM9XIPzjvX8P6kkO
TTs1dOv1TpQym8bbA3O3QKW1SPpXXUtibXSh6SgmQjm4KUgq97l6iaofdBLu83H6
jxCMIG25BSLh75vcTJ91P0vjM59j+Hppdk858EOPqj4oMnEtDu3eJzzGPfY8ZhQS
GgcPUGO0tcxlQVf/gvcY58GL93mZveTRl/Rqh8LHmtiFoLqF5lzMrKYxxmHhyZcI
T/xu1JIyDPEnC3M70uJcErqPADVZAFPs/qsp9yLuH57kO9ZDI5QMEf4EKjH8Q55J
M9N4U+KnbhzhMzBzA6KUMFb/vC38SzEbzDOif/ZwSAYAj3sPw1gQLQ8iCr0ybk+L
iD4wyjbtOqA9Aue6TFvlHMU+htcyXN1bCSxIz+o0MRE17VDiIWgLHyRC9qmJu1ED
FWwDgEslmahTOSbXDqidbd+0s5P/w/nyH45lEIk1CXT7I9jB1eT0ZcmPNY3yU40U
TpDOu7xp/VZviaMt7dx9wvQYYFdc/oSNDp4TDg8GCkxruSvc2bgXgHSM1U+vDl9m
ZYKeShr3ruv1vaE00O13JAaltx+WCW3Rt0XMDiZIwoPJRSH0qK+WGSXL58rvW7VB
hB1rcsOBM0PiSmhTgfFgxVUp4wYopWdpjy2z0u+Tjkv+HOaD8vMQSOlrHF9yPdZl
rlxyBVs0r3xlTV2cgR76615HKwa7PTSAyxbJ4uXRFkoAKVsiLF9FdPxUy3VKkHuZ
0FTLbtIIszMne2RwnAKimpf/N6XaB0PH19qJW/ldv4DD6VZqnbcvwKKEzvOI8eK4
a9DMll+3S2JC+oTQoMdkh1fEgtaG+ApPNAKyU3nuF68+XOovN7uZa5p6jEcpIlnN
2/Gt+6UuaXFt9eVC8jFo7Cadilkq6L0NYaA72WsW+POniXiUZZJdzc5o+wah2rah
`protect end_protected