`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 1872 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/9huKRhRMtvnNqb3Z+UU7TahEoHV+T8U3P3ufru7l1O
3DlgtZzb9QxCbOjthp9+wDkjygH0eUfDrEl1ovhZG63XYnqrmE/DcdVaf0FWH4xl
Bg9j0m2wtlJZH1tyKOnpBR5kIYVbZIXVEMsSkod2obvCX12P4d0fCSQHM4wqsSjO
iKYxX5XCKXM2raFcRiVOwvH7AFnFquDCTRWK05LV7vqbPONUOo8PBZcmei9l0fgG
3cLBMsVG7KdVAuJhPABnXUKqdSRdLm1G22haYXRgTA3u0qhCO5f2R3RDxPYWd6xt
KBLTiy69Uw/L5ezf+sl8xF39NhBlSkJYxZRTtEyvZvZOBml+qZ8UZOe/oUEJoURe
YLeftOcuyW/kWi9F6DrrK7WTFovx0/Hz7XPJtdMv84iSmwl5IIDAvcababvaCcTV
DpcGUYhHCzP88GDqjPYOYpXR0UgTuUcEvA20NxlJx7lPcGBB3NA5TqVkVbIAB6TX
4lJdWMsa45hnGCFozyLJJgHoyRKzLaZyF6zUIayS3n+tVzNkvkBR0aOdXjF9Ht+z
vc6Xha3y0YbsM+x6TCV/c9Wbz6xiliCr/2oxfVUhPC+oiYuBzNS5+sZKGWWwOElo
hajGUk3GUPwukMahRcvRMi/6Hw4/HC0Eq9Piye282VPw1yCZB1ynjn32aUp/0Fnj
+27DCFWe9P9gIbg8sKlZZiJ3bB6gr1gMcS/Jte5MSh+8nd8PPntx1yGPcTNG7xIg
BjSRfWF6t0IAZO3dHRKatCfuAIRLA+gMGHCb8PnkzexVr6W268Sm3zqaYhMGzN5S
PLrbfObNXMqJGX9SZzYQy/KmDHaqJf6SHGCQB24/UakBvc27xAJaflLzFKD3vN3/
pPhWIiwO30otxMtiOdzX5BXYIAaU0Fnz3KDK/4HU4zlV/+l0hf1/4kWeBMEGST84
u3YtKtDM333ITyVPBQZcWLe45RzD9ehChoLjIt8AdwfbMAA2GUs4zVNmiOB7Yet1
2Qe6Oh6BqCkMuUyElDpS+4pHLtUCCEDX6z+hUssaN6RCKJULVcetWEA1daixFDBp
rYmZg3C6lVRy3TIoi3Rb6yljXQDKOq+jVwpLnRagz4rKzpsVgTSRi8TV0K8gHm0P
LccXX1ZbR9YR86cbrnGf56o2/Kb6e0mdPOHU/Q7DRxgCpPGhqKUWEZzQh5XPUHuu
cvQ57enHrXB8U6zLp3VN8/K3cKDuXtmOFLi3A+4mUMoL/suuXTsDG0hSNcv8toXr
h6Uvo1qZgoU/yDneTUCu09ysu5ycKiU4tLEw/SqsEOs8pF+Y2MEm7E5Ju+M9Q9Yb
9g/Gw+U/mjXDD7zG1cpfBGlpUcond0+bSI+yIbnKZKrk4SoyfQ4ddWvEmiMG8FDM
yx/X4zqrRBfeP05+byBOJDaj5rDufK+CaiMp7/vtl+5jLu8zwCbSe3PxUIFh75Tm
oqLw2nuftOz4eVQFYXZsOnMYpGYziqcLRvH26z6wxkcIVnH9Tmda4w9fWswea/Vu
YWR33iKm6DXEscbffPZ5oE37h6e88j+oZSwEpkWY2i/XPhLApbxxWJEUwXyMANSy
0Gm8T6V+u8d491460y7WDE854orMBRgJt9iqiIWcTupa/5Tt3qLyi96QOoZ/s40U
e2Dx0yKhFUa0TQUzgO84VjcbioZeZWJz6g2UBEMPebfBnhaXnu6ZZJcvuQ6cR1zW
Pf6O+jSVIh7SpG+B8iOsvJz+I4cZlxjP6CCWSQs6q82LDXftGFBdeCTGGsXXb5B3
jRGc++qTHL5eUbzZ6kCTBQpVRRbBa4CnHioGhGOVWg9J6/6pdnn5wB5Y1LhhQ/nF
51y817U18iP62l4Epncmpwx4pZP2Cr3cdUz/z4IMPi7Uxv/VfLcFClw8epAK6H45
kwmhRRUfQMwcjLvfrOpfWmZrktAni+nele25y0yAXoQw53+OoEdnpbZ+FzkAHdRz
cIMVCsESt2rakbd42tcN7Tg7aTtse/yooK9vcmF3nS064tzgRic34D5Dm1nYuIFI
s0f6zAJpwppMgdSDMe/JP4ZVxUR/l3Wzqbnk0N53KtwePg+28HWHD+JAZibmkOaY
7M5OvJ2y8INJdVIzqYsUdxpjqAV3fuTNcCk7QcbujdZkZOvocMSNxONccVe9busC
NvUG2tA2NOnYok1ZUT+2rEnRDDg9pk5Lb01oMd/DbsX+mQzg1n36AsvToE2Z8G65
HvUzyYDA4fwj36bpFDzwRVBIGdMI+wr7VqEtqPG92vJTKX/r79PqxthfqwONP7oZ
2upKqO2e3I47AkgJTSZhUUuSnHTb/lArxkzvojgkzJ+3Gw7dRdQ+48IjZzx+hAf3
zWC77ZwYZ8IHB4RVS3SXAIjjrxFLe0coZ3cvM+OxA7MlcHcYqqSoeZTB2AzuPH5i
NxxiLlRdpU+zJGIlBAXgIiSWTL05ZBomszJf07bNfPskgSutSWeU71jPGjMOtTCh
`protect end_protected