`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 16688 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/9huKRhRMtvnNqb3Z+UU7TahEoHV+T8U3P3ufru7l1O
3DlgtZzb9QxCbOjthp9+wDkjygH0eUfDrEl1ovhZG60mIcE/QXYR5q+Zy7/GbzVc
cIvqTXouboLomrtSj4O23fz/P8lkBQqo1zFZLtZOhzdx31aFS/Hko1WN2Xc3PWC5
nQuSNIe543jiaE5W1NPQyXI5DvRYClEZmeNC0ZZp/CQzADUFS6uI8l+jt96Yquow
ue/mszBTD/2zKosYfNAeKp4FOkK3ocir1kxkuKjp24dhcoTL93XZ0yK7pHv1A2jX
xsNKXYzTOKq45e5SDXkMdYy77xILQj5MMh+T6q/DErhfblv6tvfnvvIn8dxsMMJV
nIsKfKQ5DjHl73D/RYgEMHrnNYJ6ai/70nZyLR2eg8dA2GWLWBcT4KbY/CSGL6Ww
oZVsdbTw0vWgwUqanzYS1HGU7x4XDoRhqH3ITwDgHZFqitS1F7DiNKD9XqLVQG2E
CMeR942c90/IRveYaEXUioo4YXs/iVKcgx+uKjc8mWVNYnR9bQ104kVlH17izi9w
w71YgCHC8bnYCeg2+2JjVzMPRM0sgBpPd+xV2GowgeNzMXqq6zlye9v8YXA+DWZr
CFNQ4H/gu014MQeOcHMTM5SvobNIZZlzEXkF31PjUu+2Dimogw4OVpi6S8cPcTnK
r0am1GeOGFyDf2CyZQUKFaIXBpM+SPlNyrx3Fy5h5bi69T5EF6p2Y7sLe91I+wCq
JgEkJucGD/Neq8tGzzqLYLt/O5U8myu9eodfcs0O9NlIq++fDj7qs+oaimUcZHYQ
nSn3L/vQDgtCLU+6zhRdoppbGfrbKAE8q2AFdnM6YSYoOaOyvOer/0bMoGRley3p
qVkdNX+YoJYMhcKLHApe4KPqR6g6l+cThOQ+FrQifJepVDodp57jrCTXbJWoD7cK
6ttgM4jL3B1u2WfjA6Fi/KEAz1RE580Gl6CdKerKK9h3+xKfkvynUqdeQPL+zpEb
ckQH0N5qw1bAOwMTGbbsmUbiZRPkWXScSvb+IwWR10dZa3Rrz4GjMkP8XQcVtJ9O
EgEpb5Rdo9jHh4euMQRWVgqrsEqesWC3lxxxnZZcy1WixtH3IPqbaopYkyloeFF+
Y2cUct2Kkv4UAz2XheUixXgK5HtjcVNnnTHV9s2i25vl2qFZrlk0Sbs6c+d7oFx7
jKSk5ykdC3C6cBknv0dud84KkvbZYglEDes26iVXMgfHsBvlh+p86kKQ+vBMlzpF
0kMlfE024TfTXHPNy40JWCmMFP8OFBgNQJ+KL99m3JNgIjco2uZqctx0m2Qa8Tee
dL8QFLwhykQ45veyQov2naD9jIikRg/3RHINpb4HJkP3JIxED7yt3qcwPMofyhmm
o2goK4dE5Wm5/StWtGGJKoGGdZfOJLoFwwE2OnBnefSla/6KLHJ7/Glfq/dV+F/X
wkqSqG0aJZ7qIwJl9QuQBHezlU1T84o3S4kp0OVVT6DN20LyKpEW0fyMASpct5x9
6y3fvz7En355cHejocbppRpsQ7dEvap59kHdFvM/fpbwbwAHUWdBawtrFSmDWTlN
VqAxCJ9wSyvVR6rNY2llKLAYzow4hR5NysfUiZ2yRRx715qlhK+ZNSqF6bUHsg95
GZBmUgQqGzZIrxK79WBC3yL6tMFFYqZMFdrrqjk+99A0/epQEj1kP3pxCornnsVr
bklTgMdYUyuXynQQ6r3uDhvxDa1WjXmXVjQ2foYAAom2ZnXg9vcWkNq2N4uE7ZXl
epWLaaOGyhaohdU8o1PuX8E6NQ9HV9OUdFZ30sv6oGI25VR1L6rQp/J/xHRHmdyK
sAk1Qz4bPi885zYu5OSSCBl90wE91JDaxDZsnGh5itfslAHMjatYiZYpqoog4cQZ
mJK8ooTty1s9usvUeqccu3rqr0xtUg9ETQ7n1V4R5KqlPrsu/mYWcPHkzZUiBOcE
O79pjMKjl9whjFvASBZd083A5+eRj+05a44cYeB20v20d/HAAUo9KD6klVYBjsc6
9sXMu4mI5Li2kK79ZQFuqPrMZC/Odn9Khp3iCbPw4mDYjyGQM1260/1fgbLWS+bf
GajmGXgLpKlKL7Dekxa/JxQz3wsOEr8WKGJvdb2ebx/NTEkS4dbUG1ZzJZdQZca6
Zz2Jdc0Fo56Cy/v6GTpE8DGIo+dY/MYMXlOvPaRu1wox3o7LvhpiwRzS53F0mjtP
ph/nYxQyT2AJZLybni0hs8yzb5jaQZvgdMLvE8FnQnBPnpPQY5CJTYD+zfKOvvHB
Vgm3SBN4r5BG/66n9bFKR7o0QYtqbjbh/bMVobdAVrtja/P7+DJthTZAMMpeSbdP
DtqGoNus4zgfgtdF0Hk6mfvGFxLZLifeP5dxIO2XNqmcBCDDJ5mEWVPBy3nm+QgE
Ao63d7a7WoyEMtp9yHWpB+gfjOrZjiQH6hXqLyqRfEcRLPZMOyMo5rGy0xemANPV
hBlqmmfkwGzd2cTSpQg5Lqwhtv8jn/h3+Da7xGecYT8j1S7/EVzA1GF+JNotT7Qk
5RSmaX6ojeFtR+fYppUA8IfWI5H91ybZoQD+EY0D++zdYnZ87qvkOe07F4wH2ynY
si/cgINiohuOjtx5hPV8y9ViqdhggwyYOUzjesXGJHZ66VACH+K7zJult1XrSf/a
RlwhXwFxY1LhLuzWidKJHYDpueYJcDLlclDpA7g3XhN2weqauJmz5Rjr6z4h1sxj
71A12DsH+Qf3MtglYObcbrUZ4Bd2PmL1CNz4LcWXuMzOrWHV+Z1F3KG44RI8nec1
AB+ok8kXjIJMzrl24GwI9Inw8S6l1r/R5TLqKgCjFE9HbAW9AkzmCoZVPpedHTGe
rLC8YQRWt2B/i/xTNYqFFlzkRURlKGB5Lo87LQ0fqYc0KRJ/6EpZOWsLac8slld/
wDQLx5SeV2vRwQlDAUUi9t36pVxX9Z5MrMkzXUDfCONbLeKDAfwccrSA95OdFn4C
mtb5gE7GCaTLWYz3nwOjQPqzXiK9aT6PYgLzZu71zjgTzSmspx5wucujkoLVSpVE
KqSoRsoqYBkfJZUllJ8dmqHhOAviToGkVjKdB5o4uDfRzYk1OYKIoxVw6ty/++NF
Lw2y678MqD3zoD6wgbmH7SQ3mu9g9cgN+IGuAjruAiZDVthPiQddL3J8bE6ARMVO
HFlS9faxF/p1IkdXkk0AbSXbI8i4usHD9op5q4wdhVyR00is4/lNnjVKkOeJjLP9
Xqx9fj8VS8mLO9jz3bKIM8bY7MGX8GDtA8/S87zt9eU85wNbgPFakvJe6Ce3hwiW
Fb2aykzZqI6nC67NZpS9qkrQTVfMhlNBzIXtglQUCkRDUsSRz9jimVuv9hrPm+3h
KiTPZhND7ObIpbwJfvKpbO2LntizhEP58QaLMANbIS4pah5NiqOf2nU9pntjksab
FxC7/5W6MAMI1S/6mfnAKszpELsecwT6UZvbnNhghKXzT3iOiHDSFG9GqzF0C+C+
5QjM3Rht7JNP7CyqUmLU178u79FJUb8sxyOAt8Y+tBuc6MNAeMjqwe0AcXp/GhmF
ocuemHk6pleGKzE+Li+d2ZRZ2q5M2LppyX7LgaK9Sax6lydg946ToKHdP6CnwTOf
ANWkfoKZj1rR54buRIp7RnyKoLg6IgYorcJTNc0Vwy075a9JEgzsTJpARixnWtb5
JV+hh2tQkpz8cHScoao0P7P4+8PAp9mNMLFoMEd3cNlBe5/7wwkZPEK2cAS0WnJy
smRup+HiA5JmrfqrRhEnbLPisizkk36Sc9196SAV3zG8D8AduzE+sa599qGEcuil
p7dR6Cn7+oPPTX3US4kwXIa3GbEtmbGsOswwytTdoO0hTbvmXTl2RbEdeLHbJK45
Io4teyYpwHzb1v0o/pDyJYNf6na7P06Hry5iUjJx8MrADFiYiWwJiCld0ejaTtix
WzH3Q3OS99l13KSth+gqPFmwjy662PRuEB6NSxJWAVtwlMqD8mgXhAyTaZP8DgLs
eZbttLLRPAu2ombTWbt1sY8GxD0fonxdXzQUe7rvaIk4qzIkhsjv3EdIHjvyUnVT
AFwQ4105pNgjAJnMz+UiLkBt9QBAYpqmYbBGydlqkDU/u5rDD4VRONsBq4tJqWCU
5N4y5Mzqdq05C1HHwZi6Rz+7ovvCdxwDEzuk63nDo1VEMqxOQCRuVjNEd9qX5hmV
f9LyaBTdPFkh+Xrkp3XwuhrBwMQIyWnyPpTNNXhorZK207QCHd9rqO9FRFEGibz4
2wlBWJ2DKJa7OHlZK3Gm7mUNn8asBPWVMyd60siIWAgS8f5klFul8CCS6FuBTAcu
ccBIUSBOKpiMjTHTGXImny5i5sFZZCx1xday5Z4ncBWKn2WHyXF1a/q4dfaC9m22
xsnrZLTsO61Z0SS7aaaB2iVm/I+ptf5YXzkt+S3kgKxalFZg+BepfR80fkaBPZFF
rUlHPcKuIpLxPtY3vhRcNkpYKojT/WkCJNVplMK9gZnDVNHi8Uw847i0SQZwUDXX
SU1brImH12SBdkGhPMBFFEyRPczK3mN4dMwvLwMU4zZHLD4DVir+iqfe0k9XMnNh
lagFpdYDazd5QJv8MB2CIlrKTBIfHBpy7Lk5cmr+bTN1lwk0aBcsmukLG9OK4MOH
nkErL4nutvkQgods5pb16Vusygzci7OJhMegadiLUd6xZvejwBsHbqiw8PZrtF9+
IfMi/dTIBOmdCH9Th2e4nl4VbK9f020QUffhwhdkMrNro2kXiwPaHpKK7Dzdiega
2Xjk31DeCcman3En+SgCMMxOPkHM9lvS2dCT864P3H7Qn8U1nvKPX94ojfij+Fmr
NkJO2rS5sVxOao08ULXRsa09W8+HJ445ww21NL8Q0PLnCYK4vxegk9KIPq5NjLYz
EPlNA46po7HZTUQn+jLO0ZUI8innwDUoOF7HpTx9GQv6oQUsU3kq3uppw3NvL+Q5
i6bDalDSRBN3jnb536c/pr9QTnuAUHHet9QWPTQDDtn2hMsFjYUiR7DdXgFPZsgk
2J+BneSvom9C+t3UV0/J8U2ya6llDoNzE6S3k1lFZjpLJB+A16iwq8PFHjojU71D
DssFbMNCy3ebjpu5qCzjNKAICF79vO8yzinceEaD7yaOpQqubBnSxJVOFy/U/RPn
tvcvz6ZcTVc9nkCp4vZQG1w1NqQgzykGwjYJH5MmnLWHw+dvisOFlY16y7Bzynay
f8ziIIAdXm1O04ecsKSQ9XloYUAbuIG4iK7QWdaCoVfMQEE6thOeZkBi9NSndAWj
i5QYicNBtTmqWT3H4iBjijoaRKwwk9ep9zThZp5EkAWhJn2uFkirRZYXQxkRqRC3
fF/PMm4hOZft+8gTjJtDtz9VbBt1EDL3FvmycWtrFBHw9vU1jOwkxsZoGtu+cZ/w
0pJn3y+ttksFgVQ3+VFuadnQJBsYSCShmgfGsx5erz2eqzpjKKN1ds9lvjthTrEv
PrejT04EB/SQ+DuKxyxz72HkD0qiXcJCnN28163EX9dkDt/PPBPvOTef90Em3I5F
+7skcq0ztfG5qwpKJcuJ0gCXegzS766l45lDk4yeJ5kUBMC6tahS97PPWvjNd1ux
PmyeXaFC8L7kMATTDCBfkK0AhDvhMsfHFWwG7htUiFQBqaOlyDrDZbP52syFkjtY
r3GQ04RVI9OdNhEKjN2kDuJR79mPlo9ITyt4vEKtvIWVw4gPy2JixBqqdFgO0WVn
+Dm/PpWEVy1G94yreiRIImdtk5/K9JlJyJwb1r+I5NgeK5FfMPfWyVdaqVscGkqL
wlC3noCBcprpAZlrghjxUU+lkQuc7h8Took3uiGhHzF10GaDA5w+gQY6hK/LiiVr
iCGQVKs2OEAbLS6fQlggCDwhAjkY00kJ1h+9M/QxjRpfYqzaclvEB8TC8Mc730GU
SPwFzHdz8XF8BICHXZEhLcOtW9OX3U7oss+FIwLEMn/k3o42Me//ujWZyBveLqDb
VTRDJ8MZSqFjuFwnRH4dlNR9yQq8iThyjZgo79hdWpXZ4w9/vVu53prb/5s0BYid
kilDMD1339bssjjI4pzVc4oYy1iNQsq6ShELSnfm2QGjOlU371GMYLzHOCefr2Wq
GBElqfKWbhRcyExeW1dXJE2hJKZYi4AWFgQaTF5UiHD6awsJFZ1kYNjyqBIhBaSh
xMbse9oZJ66YSn+sCCwSaxVsqz/3utznaZB6rP3XaBNlyTaKNbpj7S/VzSLOCdqY
hn9b0P/cMDIUhqEBuvj5K3eoHPhICRzGFRGFu1Yzk7+dOTutKwBhGe7VB85PNsiS
lkFrf2vqhA3Gu0+827WOybOtGyk0YfTFQ2wUmOstoIh8BiGAiGvyZ1/nWYzJerIQ
175nz18kZqq24iygy2P0OJPbSVXlOS5/NYrIrp9atw/dKzIDMINrIx1FFhDLJePM
teAUBBlPE0yMWH3HXtzSQ7aQ4zhcy+5Yh+cjKEzZ7hqWBpQJ8Edk4M53vkl8iC/d
6NYwjBdO9QNUvE5opc6crfvqfyomc3PjuFx9uXjjKM1YEsUBSDvJDCh5GEBmuy70
MyD7/nhaS+qGp0qOJCfEC3Kc+i4ceiw4w/i7gKqWQ+Kuf0VbeLO1KMmUPJDdoh1x
REOTj0L14ee0HEVmQ/teI1/1LwZyN7Ydtq+lTULBIsa0CkUvVrTyO4m7CrgytOHC
hhutFSBf2V2OSM/pcohD/GsD6hNWrZNyCp8oBG1l0Ty7cFu+wKy1KNFn0FCqSTVG
0HM+BxfF682+R5hdBn8O0f9fXdIv0f9arz52oDpmfSMUASRY3x60KGRng6QCF4Fx
X+n31SZpnG+8NpUN0XCzGQdqzQQnNjlLD1yWitJubi5l8eUuCmg8Eia9ViI+Fk33
70F2LndEmvAzXZMY+9nZIgasl2Kt+9vjiaSI/h/sWJ1PBhbGNb5g5EzgCIopL+RY
xBMOCYbG4XFE89KR2STGgSGfm94CLNu76XE/OjO5bFU8IWz6uHSJNuJm019NfrUG
xGqKf9xRePRNwx+noJlE4xvucFBRcKFNjGoX6mrwBv3H+tGdgEawr3RkZwqh5X6J
vrKIVJrpd94JVoB0R16awLzGbSx4ewD5y3H0ngLdFT6VasgYgTpiLXIwn5phkxAh
GAI9Qmtehh1/XsCpdgVc6xQ+HFaSoe39cApbl7Xdd7xrwZbNA3XZqgC16dCmpxaO
XP0AT5yzjLxW86icKzdsQYM2I0V1CYruyjQ74tN46NoaSEjaOe0vok7oAaE/FEI0
LGCs3wTlQb/NCRdyNrPWAWLzfwT+rixCnxzHAGUQte5EqjydM8i2W+RK2KDE7KVX
XkK1UGsFnyWzYkAz0ap3nGn9pAYioiRVoqko0foAlarTPAdRA9LSFQ0XmCDDIQUX
ZLHgmhGi5cfbJtwC9RRjZP1A0uGo2193YclsaiJlEjx/ZDG1Rb+f3p+S5ESUdbtO
QZj5gBubCxUG2YGcofQFNsB8mA9fZCdT1KRAeXgUNCAeek0cijPckeV+X4fPtCW6
+EO0C/CAPrC9zFBQ+jt+qdSRVlG5ConKLoPGtYY7qAA0vH96r91235uuKDt36vsf
YCVsqMPPB0rcDJCnAXGOb1meiDRl0m+oD5EH6v7NKEkrEl1g+7FbhryWpwzO5bVd
EANuXmcxJ5A/T1Hd9K/Fpl5EQ46igwuJoa4+tRDS1cnq6aSyjoXX5vP0Q2dtys0Y
c2WX/WEMXK5GreSm2uJ6n+2G6B3c0xEzpDqz8UFIPKWeNjZ6sSMz8XaiozCdPiw+
2+sYej5QhucVYWcdG0+FbNtrIQO5bMnjXIBBYmAob9/FUJ1oBVjLnzRLsgUvmLIW
0Qaicbxrlkd/IA2zc3BzoWZnmFEYq58JsAM4wefJEfM9svzRc6ospda7Tg+rls1F
myvkPthzZCNn/w5QJ1nNMbPrOi1wGASFmGBFJ/4fnujubldZmtmwEt8NYaWIL9Gp
Hr6v/jFb38YuxbArGrANsE/BEiX2GuV3wRKEgVnK1s840RA/VqgdF68qxIrgt+Eo
LYfxlRB9ESzSSS6tmyH/USBXBayWMv4OFPTlm79KYA7ee1eeSaQG1PLaWYw8ZTFe
jHbtw+o4UTAaOuvjtX7NCvHne+5HTXbPFFkTzRlYxf8USp9YEQaznYBo1QT0ZTxu
KXHO0xUUBiYtWJxnYI6Wztc+CnnhxzvlXOVSU2jMZ3JSWQlphZlGFSuBElEbDtIx
o9J8TV569eJ6J2P08CB9ycDZGquf5aFW4Go2P24ZdVtdpY9Bv53dwEbSoIAqILgq
slg4pM/vCRnf3NlJj2fAI8F4akAy+Y3keUpsk8cFcDDFzhdGnAqINIOmq5rp2JOQ
K44S70v7B6/XEgRIk9fCHpIrzILZxFHIxJlbUokFCcsSHyYcmBVzGkOolaW2+KD8
1UrSgFdfA0qKuC/rnfCNN6kaWPT8wWmZ9AgeLlXXrgiZ3zkEzlNf0KYgjezhxpIn
kaDTvKEhItdXVTf8wPhoIkZ957op+gK2TOXqDj/2avBY3sFTHsWVkrLGlxXmHeLg
TKpua5FuvvHW8K5iDE7WfLp3mEQ4yKWzLYhwiPXqk83Nc0sy9EtvaelhGw7D3gOF
VYvhoNIezq9pxGJbS8swGf2GovI6JFvuBDH43sXBouDApG4uKF6EtTMCmiJ4ZxOA
alTf86R8JTTtyUvTZNRydx8Fpz8lWSYykOI+celo0jjOCj5wWcbzQSt8J7B5QRek
2bViOrV0+rFHYNv5irDaNLo/ALVLIcVAycGBuBVFcSpY9qKULIdylrgHQQXEAhY6
ynHUq7kdBxor610OsrOvu8bUQDKjkcRCtbXA2emKGcvNdNOB9gUuDVmHksi1mYtL
5HntxPuuMB8AYGYf8qenfdIu0pjGDeBX/eOWdgvwFxbMu2mLy4TcPBsPoZtDbIQQ
t2EIdfowU6Yf9EOPibuSMahRhXLAOxr6FFwoIDEoZL8B8DR9t3EN8YiqefLlePKD
HPkcz15E28A9+UXWVYkgOQhPuEne0Flr+UB0Brq+8TXFfTCvZis9TXUZw44vmLjj
IoVi5crq/sFh6/Y9r8H2eRQ+/omRN6gLa41CqrTDyBdlYhNEfc2gHNWIWywTvhZe
mUtoJvTSHRMea687PVigjL9fRK6utNjOyS1aDrpWeH8CndHzkh1k3wwhy5ubWM5A
onnHSNEwg0YKMfXBvOXUNG9k67CiSW3Cv7HRISk5stBERCpimbw6jEgOkqIfEUKB
vtjqk3sDTR3FH0M847M+4PmTt3X278i00ESLAaE/JPsi8TUApcKL0033gDL69nLq
Evk8Lzn5fFp0meTbge3ujfrv82A3XAM5pvg/biup7BfLmA3yOxGFeT6W00DKrifq
5DHQ6u1Se309Zk9F349UHJ/qEUG9pEo4V8aiW98ytyzBlTU9HDBaW7dJhLtNkD5O
qOIA6JFT490jTHzssRoJ5MoCPmhU1lqwEMOHAcoITgKd6dY4UjX9v19jNjB7Rxbn
BRM0T3HmM0zJ91p2aAbCl1Rrt7j2mZEdefw6I5hoa2nmD8VtWTDCj7lEZTjxCzhd
ERDhAQT9Zx7K/RdIb0jpNUpQs1ny3DNsSuFMg8kezFDBM0cV5FBlnUUC5gDzl2Gc
RTrF1sPDNoLRirCqujt3bb2VV3HTaDI+yNrAu2WxSXbEm6Vw0KWHFm8J9TQwq12e
nD13RPNpcQMEyznb3x0NQEbENRZpwk6A2xA2p8pXz4FrPBrI6cfa+OK75um7g3ct
dynynPOEhj8wXAjGZROdCSF5KMqxp4mZ4kUgmVpCshIArzJqmjQQK2+Bbg1pzQE2
o5Ieu919GeFmxg04dcnYnYAak74VLHKhcQufuXk5+bXbIvLNKr8J0T220URgT3Pb
UFnJAGvVUi6ie7r3m4E3uxhuXG7XE9QYvqMVYHhnDgK+2/ab1VN/jvF5d+9TqHlL
fVwu+CdmsMnioW0n6mmUdW6Mv7ZA98hETZ+wbi6wzKPyrHoi1jwR2zfTqgbLRXEk
nSl6Lj9RhQ52CceH8Oa31aJgeilK40V0sFDvnWm/gkxrVaPmQ4/hq+32vYE6vcpG
emzbSFBjVwYVWcsPVHDvaVJSfO4axXkbV/mM67aQT/gwUsHm/irc8jRWCpK6fuMF
YjNI98ovftmOV9k1hAJztx4ipUxaZKAgZvomnHfF5RVxK7do4t+SHj02+nEf3pNb
OO5zo7SD/RiZh5GDnzCLbV33zbLtB2b58fK61J2DMbWZ8jHPGfUyYqYdCTIA0gS8
wUDpJKcVZbfZ+1yL4K5HGf6UYbbCjhOe8GrMVBm28kAo1VShCeYJliSoTQ3XuBjl
H11Ir3PeOZdpYZwWP2y7GyrfhyWsc4iUL2NJQlnj1KwcQ0sOYdcVytS2+xZ/vIjp
QtWmRsSAw0xJgGEqeTaOWSjqV2YjHFNFnNUw7r3JgHEr8qZ5XGl6baFXXah0IAbY
2r0PzbGcIWE00AwXNnavgGPVuLj2U1GM5QpHIFD3db+JyzPiIuqeXrk8R0q+L3nC
upYWQnAOpHFJyxW7lWOKV5iRhpYrHwLqjxIwkd6mWabae3qwg8Trco4gTFWz1v4M
xdQcvnx8HVQG0P/6O3aK0wugLnyQDl4x7ImKqNhHblwwTtM1j8YCoprZnXf9d1cl
uNaLdwKP4Du+thNnpGEDF0v1pjmdRNe9Em8Rt7WM7OGz3lAf0u3dPqLkZYbH4Y03
Btd+TZA4H3COv2SPki6zi4LjN8xoHmb2cYEUMSBCW6QoEF/E+OYXRjbjDAlz42PT
Cc+BmiGYr8GU7kgYqE/y/sTZq2rF8cy8t0v8DWEFyNOyqF7jBiMckH6C5sLW4/Ok
N7RNZtLpRVVgMprD+5Un0liqHr9T1SD3/wJc6YTOC91Z/6d7pi/S75jOdcauoToy
MnGckM214LLu9v1T+YQ9ub+R5VD24SpwiOODO09b0h3xhvqg5mdmSLMAvwbBYrv0
sZ5GnVWkbkFTzcdWUShAGvDZmUPCkbhLL9kRVOs1Z4N9u4wzwtbpiTYzTVbGoq2/
JnkdazgMKJafZJ3BV+vW2wTFAYQmUH1aG7HuTIIitOiFXLpuHdwwCcLZ8ieN3IiG
eGov26gjgno4ql9BQ9UhMvgiXYybXmTAqkMxViX1IY+QtFN4gv32PYQVvJ7mjR2K
Q7Cjnzjijcu6HLfPdhfLg4+fvYereJ6eKaQk1LJEP1K3PpSyo0W5iMc5j1M6Bl/A
oytb9oEwng6d50wunwFcIJ0lndojLKwjQ8F25Z+KoR2NWfP4nAuBce5ocUvC6oeW
PMJRl4bYXtbtn/lKCsAumeqgtFVrenB8IH6X7WNcpucvQjfm/nNTJ+Xbc1U8z0uf
EotFOV4U4WtijwI3vfWaVxNwlGD+ugLmyPdMK/5QmlG3yXF42Prflj4L+S2m0rzz
5emXJ43nJg9XfMgyTixtCY5p3HbCAxNtnJGPedV6OS9pPLI5tHJ9w68J8il4OULC
rV3gCHNf2ohOZwrnr3CghSK7LoMJYXdTybC5f8rbqmjOGLKZKgkQA9YZhaoOsY6a
IrLj4Hq1xuM9mAE1UKgWE7BC7BvklS+oxuJvcYKX6fk+L3O/gRDC0QPpXn6e61I9
s2Ct3Bow+sKcHDEBZHOPDgVfW7OGGC6y04qBLQ3rV/LZG2JfpMfPUimNsLFiatGt
fvy3h1A8G3n8aADLhrp5ocJaID+JYLZGfvbXSVbDmbrFTvwKmjJJ9jr+LlNBKaaL
8D8UhL6s5+jwmJrxOffE5k1ymJcdCorXS1VPBCW3QbFKsqaVG0K3D4XVT7gXhKdZ
XgxCY9YM//QaDDGvI3SCs3fPn5Y67W02zXqcy+y0+UbbS3O2MaBWFqxS5NZyVcHm
0abjXK6ugFyOQxiWVFJPsYrNpMst3C+RYljYG0Jwa7SCjut4a0CgyNEFFxfppi8C
sJ+Lq81Cz+w3nHdBEDUdKacpIVqhMHHN8TffilHxIFuQHFcuwuv8Llr/aAkxYcT6
vtggHIlsBaZPKjlOsThumlCvB3T+DeD465JdEQ+LXEiwa9w4lPgeSS4BfLqXlYzG
btvyWU7Uy3FSkNjDJY4VXJvm1tONzrj8N6WSCtlbDcwKOL3toiHxPbe2BQeYpOuQ
2hOGlbuMrPuaQk5mI34cG8KwXX9Ka/zadl3BLZ8unY+G+rLN2ZHLsDon6XE7LIdj
apedS2R9BTsgWQ532JAdGtDNsvogl8qIJ50Eb0adkqcccFWvL5ZM/GkP1/LTgtGf
K/+pDc08iRbskmUW1H9oayuYq/BShkiv27lpk5rSQRV8btm6r7IHsVFk/J69EmL4
Wz3nTKGHYS+b5TWROsHDIGPX0Wp4kQRLRVl3vE6WwLMPDIHZBuprvVnWYyjGPEYi
XMhR0KVQ4+Ep374Dt3TVsS4AIpOQ1qUsIM+euD181EhvQG/+a+tiynL+B40EtdYK
6ATNdIEADezqGicSNYU6usQENT7/fRXyvauml2tinPszWB+5xpJZ7mg4Z6Wwpm73
ogPBdMSB6oT5fteffM3gwc6dmX65LKjkc6q7rHfKUYk6pV8muN4A3ufZVPUcvZ3w
p2xCxHqryOTruu0/aOc9lL+tKY4z/bZxXb0yTrVsDUx4T62vYewV2E6X0/dVMikk
OEGLYx9ioL+lZw7IrPs5UymGmF0lMxP8skUPPzoCM4py427d1sUqCjreyyDNouzf
5qpzWBg7LuI2TbIPiFTX33wgAll4dDkTB0djFiK6d7fdH5yLDBoNicISTnAe+MLz
2PqrZFqoTyz6ChdhylXf0KdCalfUR7eDWBQgk8/vAZ2YKuk7sAS/eD+La1KRO8ds
gCNCa4Lbm4pYiwRsjhGu1ZeODENgGJsHz/H7wZuJNpP8bZD0L/toNbjfoodWLTyi
1JUT+GpIpNgAM3FT66FfEcegLsmG4x5kwzLS+2Y8tEffIu+NynXicO6YPD8mBRON
K8RoJrpa07otW5objwzRS4NRnrmL/1xuor0xUVfpVzokPtsuZACJx5kT9J2lMcAT
JfSqnYj05Es4Uj8bWVrqaDthpAXYLrT/Ji1clZvinOvOaYY1a1bNLMhBeniXhrQA
Eyx6pB4NXN0OBFLkRoZ+d+Y8YXXqMiixNiomedJMGkAb0khABX6ApFCGLyKpC54z
6RHRC6Gd75UlMa+xce4WsWUZAEA6JKGQi29UiNDgzccN9XBMLIKnsfaF2Rzw7cJ3
QVUdXBSUlYOCmHTaShRmen4yuGBP1Kbxqm/FBOEhmVNUwAYi6IHIHgzB1ACu/DHd
pPGsy5rg5Uyc1A9YEsAFqtqyGGd34wI6+a0fXpIrCnfe4QfeQcY2XB4BwfYlGCoD
BTUOjixEcT/o/cSL3fbCSTpnUEqxvRzFRcUalquZ4inZ658yaP7OQOc+lNrUgPE4
GQub/a8lfvHecYT+9JcE1pV8N5XNq+2B7GoYRgIt7NWYHm4b1aLvJpVH5Uw33cMf
S3t8Wyg2WXIMLSuO0QakjfBeTbucNReGWWojg0CnTYaN4GDNRpA5xZ5cEsm9Lu9t
IZy8elNsu1BpbVJwXZguMuUNk1JwZomCskZ/MtwovHT5XfxKKVl9I+L4Y5/a07Ma
v1CqboP+e/XpaYJKSDdCoS9wtqnTtYYum+FdIFfaP05LofCEAxp+5v/pVkgm/Rtp
58VM8rIKv8I+fT06L06lCEeWIrI8KeHAfwC9VYsfhn7p3U2hqYwGPYIo7qk+urs2
LDgPhfpS+cjZ9GpMlEkzDqgDdhqUCmjUVsBOEpIcgzU7XhJtqdYMsKf/RuvyNfTG
VKyQtFn3rkH6aVVDQdkGBJ/0apOaUoH6ItkMdTDGfQzGHC+qTi2uQW0/JztfNoC3
c9cGlroNM/TGnw8fvAB5kP7yz7F88UwB8RQvwPmuM5pj5Jnc14ejUCvMfF3ap6Sn
9Ceh2N9nqwUx28kW3VloJxScAMPe3VeP7r80G0yDD5TMxRs/cuKkmqLiBOCat2yL
zidqY/NyvbwiqjqR/n75WMreqmgz3b47i0CaDR87gxfYK2oJFjM9RL6hqXRMwfrH
rxvG4iu+x6SnLB5AuAPKXlRPQrYsaaDOepQV40xGa5G070aptzYrwhjt4fIi4AKG
+98VTMjAnfSLzfcJhMeCCf8ArVGn25YlCLWugQn+dNoQb8/xf6Tm9MVJGYOrA/Tg
Fdb/4YBl+cOCEzzsul2SerOug3j0Wj4/xX97D4OzvgBFDBfjQ2g1pSLkEG437k1L
thRACduTPNwfD85K7vVFrEhksPnT0xvFf0U2IBPqCHT7Vf2WjqP02X3lb19z8WjL
LSzn/xB89IlRpzJP5rYgOqQqx34FSs2ZdKXKhxB8fJSNFuW3QSoxtkhrycWNeUMg
IRKPIzlOngu5ETjoNeg1NeUOp53xW1cSbKw+mArHQpeGNSPMcYmwbGE/BiYh+2Fi
5HlaNp0WYZZ9VQhsFUxXAzJEZS6jC32bzblr1Y4zVRD0Xrj3pkPtsgPfJr6zq+lY
4kOQiZZNW6Asdvq7CQjJTLkA3wYV4ohtpEagHZ7RQUtklmcQKjug6bS5QpCy5otP
NV5U6zM1jeo0DmikBf2dndd6NIztZlfdJN0NEVFS0CqNHT9IpcI9atvfi48W0BAL
5z4XLBNN7z/T7joadD/o9NHAbKqmwK8FYeWysTRV1uphsjpq+SDT7KtPYL+iHjMB
oKwNF+SomWhiOFPwt5J4VOGIj2O3HgvKhBdUvFMu6Pcd486nGVl7Q5vkBDuROK3I
0iEuQPyRuzq5pY3f4LJYUpOnau2OGGV8PsnnxQQSCmZy3d1X6SMnma7JPQNGkgwo
sqN5uqi2lAa9RyliiwlEH7CRbo6/ynx52XQatidx5q7F+rjosjVfC7N6BNmqT1/W
t1feY1uqaUDCuJKJGGYfjdasZ1on/hhD8g1D9PSaxJDjN8L44TZjrw+wWCOXDefU
JgmS+c3oYWpQe3DqS5Pw6s83j41MvJJvF13URt4Fdd+KT0Ys3YVz+pOUmgRjTZH3
0lPLnmvIKePXkDLY5CPpVusM5SSjoLwMObF34wwz9QAucRuzYlE/dgB2RITkGSLI
y+ImF4a5ojY5beGcGpUY1ZNPqQfRnZzAEc/FSayyNTj+vUL7T/mdnh19hB3Bfugo
7qkYUgq2NycF1jLFGDCj8HSVvRrv5oMSG84hieWeyE0gUfL3VOiC5PROwFLnq9Qp
vuvX4vzfbLU42YvzKHORogghLH+P2dhJaG9bnlkfNDUrSmfgr3DUdtIxOiddTXvH
PAU170sI3mSbm86VQp0Mm7edO6yFeKVytNN/2FpEqzwoa6VJBXgsYDiix0VBJKdz
IfOiuAuXMb9U7JHow4pg2sClnBw3X+0Na0niVOHAj/wn4guawY+KuW5IMzGEEfBT
nLXQoMrbRsL+Wrb8rh87el4PHS402xumWNs4wM1ZOcT9oykW8rYo91QyN6OGadJD
oz3QoSz2MNYf7VtdCwLGxVo4wCXz09jNKChhOa/6WkUxnBX3SYC0gvDoRzrG3sDu
C6oF8aPo4Ja8k/5XQc6cH8h0I31AFq1AyfT92d7PzA0O6ekgqV0yJBPAvoOMwsgO
wklzsPx1BFa4c0hB2SSULlKB8ReA/loEAgmt7cpscB3Ns7+mpCppTSEfOKrcD0FO
kgpy4sgSAPYMnj+oSBS3ke/EieFDVAI1YXe9ACAxs8ou6qWCvPzcrQ0nLnC+KBbI
Wv6ax9DZJXN1n+hZ+dYPD7KVwFbmFM8zx6enPXi+G6VRSReP7R7UrHnAT0k7llI3
8e9j+JjtFk266sGs9G+ZVqLeiAELpx2ZVOzZNc+7bLjv3+B3Ykzo0enORIbuCbkp
CZCIzkV4BADMoPwOkf/2RgF/UMqjAZXzbEYl4X25C9d8I6ZcO1Vr+YXree6T57rU
cFjmYhxDCPq+PvfIA90JktwzrFS5FO7wCEur5o7JJ/OPecArqD/QO0+A4XZN8jly
9R7a8v6Pg5X+KZ+QwLrIN/+zhughT8TML/EYBjKSnCs0zioTdYfNTAfRV0N2ki0g
pES4JB6HbCetJoNr0A6t/Uv0E37BWT0Nv/lrespOgjrSGKEcQqSpG2tK8OjGxlJ3
KAuUeg4/Y6VN0fcyLobYZPNB/4hI0YQDSHpCRXz84WnuUAERVkDa10lW0qYoYEzb
Fx9079Vj3ox02XqP13TFdfnl9LCDhNaNFNfIm/ETXI/08Jc5zVaN34TQbo3yfDE0
/z1RIIGdd25iTbKEq2h9aj7rsqev2QkOrNaDdVlvSjoVK9/h8CsqWOcDQzuLUUG8
y0WWET/UuQ+VcP+Y6lJH95TNTggyzp2kJyui/UZL669lXqIup06JN3qubqGf/YnT
A7W36/uxSFsDlAqEH8uqv6txZ4DGB4xYfY+L9fT46SRhN9lVZx/+dkxZR0jqVoPV
6W0I99z0u3DxRXSkyMIL5EP9KNZDLSxfUXe9Kymfrqm/y9/TMExlpvIl702Jx6CI
B88+Ypfjq9gmbuJCrmv7Upg/24PWxpCZJcRlDP697Og5Ikqe/09fBW+mdXSPPRL/
Jzh+BNb1ZdxgVVLubfjjmEy4QSr4Z6geuqz+JtTLEwDCfp+qZUNJDiKUTzA7wo9N
e05UdMnJLeu+La27G0lSCJev4emqNZx4a4qAT/x0pDIJFOm5E1+3B/2dzx0Q8YvN
5UWsv+hbQptDHWVrmcLDkalcArczqMCZQPkqurBidpkg/7OJMCwNabb03EGuNH4U
Xx8uhBLdBf0jG5ZWAX/nJJ5emk1onVPtoGC6ou6LAidbjtn2g753pzxfkk5eM3IW
q4NH9+kN8JBYNtiDK5bXjA1tk8R8gjkgRmFAaK/y1nTcWy6oHaRwDwchUmkfnpIM
OkfeAecP5nLKGeOC1UR0LpnASm4dfO/Gzd0sKo/90IzztfijLCxa0nnpK4VAgV5H
Jksf1e7dil2RvykB3M2ZVnASh0yOpP48VlCQEfuQ24OKe+nnNPXS/4EQppAGtrGb
8z3bT9rMNwvlv+q5pA9jYAoV0IXqHZKutE2fyU8FNErYjURpUgAcJNiopMuAPaEA
kHn6GW3ioAdtovKdRLg0OwV59H77dwFMdil2oZkDx7nMNDwq35I8Yg4Y801tQy/r
8vkTJEEAQAisTLPj88CaO9OkXgl89ef1/DOV3sovHg04vhNlzggtaQeYy8vtpHqp
tNt9qZoZVnQvBU9vCY3xdzNyqEWEZme/JClstWycvqv9hqsVS0wSr8cTrYuyAS/p
XoxhfGsSQd8vWVz9dYMfNewwx4QpH1cK5DMX/sKKdPcERAD9jNuSGH9ZzQfXPXuq
yHQwpoSA32mCVdpu3C5nFJFWroDp5scmyWsfALU42xCQ+KDWik4tecO5JN9XKakn
R6x9bIDaMn8x6xSEwtkLnq8UZbaHL519S49kyD3DfIhMi8aJ3urt2PVuyEy3YtYj
i4KUUdCjxnG0nnC2M6RXRKDzA+lNe0n1jMIcSfAT4j2o0iRCFOSvP6pWerMAUcUV
Jl/4CNM+aG7ycQIrSgJp0B3eCIdAc4R1o3lhkOhmE8hG42J0Dlt48AIAbeWRZxLk
gcRe6KWalyn8u3OVH32inWUiKUqN0vUlbZsnt9ZGy8C8Xs5FW68LTAdd3+kIfTDY
kLqeddYPC0GttukDORNHANe6094Aq2v+INV+4WmIgSAVYsuaS/EIj/mGgidzx1ra
KorAOrzckcBsD6ae1Ant5X1K6oYDopPQO6vqow/wwJ3t1Lk5bD04tBTRlW0tOOCX
h71ZWRfSpe8HY7OtetuxKetWQSzsThDL6U0/fXH1zKnfPVNWuLI0TcspwIm+zcAa
qiKNv72tBXpEc0fT1ZawlVJPjvHYK69ZoCpt89Xz4faOQp+rbTGZ8i95qAJht/Ok
07O6sHH57OxNAiXhznRt6sq0AcLPbMUfnVQkMT600+YB7fpsXao/pEx3AgF6MY+4
wBg3FPr457qWoQjCaGbseWbh+blFflfGXxd6OemK6ajWYMsYrzkTaySnxBNqU19S
Sx02ywe60qAIqbKRD9j6Qs4IQK53WVoLw+bwmLcUidhEfSwm8kWMSgFwkbdjZqDP
s0GF6Ev7ylcHNwD1tsZwd4qagM+qk8IMiMAcaOW4iun4d+rrTH+12Pp9AeckPBqo
XuI0HxEbOkgIz+kPlk72a/pJ872Kr+mTwaJwWdC0/8UqvgDWvGKHpQUJSx7zGuMQ
FoVZ7tIz6Um1k8dqC8KYGXaL9u83hD9U+GOdtbAoj4Wexe+1jP6smwdLPTDJkYGf
nLMPTAX/m7nM4GQ+YnhDyWZPZU4xCfIdYTChvn1ozcZ6/afzOCOWoQvNzGvVU15C
VE9sS7eVbeKh5+EBLenoR7s6Iiwx4wyaBD7EIEgH4ZtiRYVRtZ2ZbkWPWLr/W74f
eE09O6sedcmj02D0Xw6ieIyAihGfhD6Q8OOn6ga36HDT+0kQhIFLAGSpOQlp9Gi8
X3PKHZhJkb1dCy+vx33DU/JoK3KpQfA46EFQtr4d1A7WNPw6plX4f6dPAH9UEe+p
vm06GeUm8F45OdKTLrxeA8W+bsEq3IA0t6Hvv0AdzbIT3RCdmHNa0cGpxRZVxuk5
YOSZGTKw9rpcedCm5iNo7tBpnUeXLBVt6wNx5Ko8/MvzXQKfdbK+NEu5GNSqIZVl
Q25XJOLd0ayT+bWooNWAqjqcPM2a+RiI1vyyeIqK2oBltM3MIrfSabgJLXHJJoh5
0Be5ltIwAnOJIi0g2jS/c2bKFGZ/7xm1dO5OBnlewkGiyeBoex8RxhnooPqI6g/q
/wY41ajY1BEf5R08MsnNvfiWtARkRNuxxmKx18/K0jotMwvwE+e0DMFFscWJAtTL
zovXH9KMo8yv0iMmynoZDCz4HK9puj880HXxoYYT2yoaIuzeYgLkPPuwdna95hZe
oPnX+axa+t9KA37SxEkdWzYuRQvjJlxHVgw5n9Z53OPBUPJCtSS5DlRENTaJxr41
omIFUTLiw3IiY8dyql5Fwd6GzgnLjTqsG8W8dpao4mzAkbqDPROTT8BFHRkZ/anu
nWxdOxsuQs4RVkjhHr/o+NtdfqzPJDseSF7vpCHIgwijfKVSrktuGRyKNZFk0UD7
SrRAa+3tLzsl1TtOoSfNXviDzB2GLykqs1P6cYlopTw1pSsayF1E4UWp1VGpkFgs
FzkRW7Rg0yjkN+pwmTQ3vICzcu8hqBz5ASEo61kwuFjpZhCfGZSWAnfM4b5tbbKz
wWjtnYALkvWPcp15N64D75qPyrd7RAmZBnx0Qz7WV58xSDnNUJ/Ii4XXz5V6OyRg
UzEs9huQpSL57kMqUzUW6vt9IMiAB6fyZYq0J5y0acW+RwZtn6SvJJtUdn/6gqy6
rrum8vbLI4gBuGcKAOXnWIWPorKE9RJpaCIZatnXiNL48TXOnScvD0u1SooX1POz
Fb3RiFN0oBnaAPn3fw/9KYolNUuZA5TjqCFg8R8EQxDeM4ok+EUX0FEqwlLbI+2w
IfNIGpuJlJQwoc0w42GuWCptfBzoOzkD9vDZ/sAjI6mlJNHvYX7HhPQRgD18MvMU
iBOZ6uuN7IYKybFMNotPCAn9yZ4juQT8stD1z5mEAyqdPzL4dkBUkSnIb6D8aJte
fWf7qP+ks59bBnuyat0MJO8YXNIB0fOdoG8U3iDsDMJxQFK0jJcmt+eYvYdUTvyV
92tFcN6R9HRzMbPK3lKK63wBm8/vIof0cfe295xZkPTA1RH66+3+AJkebt3rV0Lt
MB/LkZsNmWEQMkeFG6vZss2/pBUODkxjAS+NkjN7PftTiiq3bXIeIZP3QiNG85Ad
e3a/A80pKjHeThIyzr9czR5N1g4SgcUrnDEEHP7CpiBastwrfreEae99cJe3un1V
VUmNodeuRb1AMeZs1h7TtO6+7QWUSZRhaBjB0roHJ++lCI5qKgx5StvbhKOCMGat
WOb7HUMYO9ZDYsy2oNHCQuJt7lo9NvZlzbjNGYbfGkImg6ogziHW2rTDF0oukCjf
PrGrUkEoFvimxFiNGPMG359JTY+rm4MFNDJ9A3Rg+FNCuqO5x7QhsaIT5yi3W2Ry
p77mq4SaVxiSCYv/dIZnwUgm1CEp+MyBrTvxiYYxf0JoLQHh0AT9G6K1ovdCy85h
zu4y8Hz/ZHzT5UGTxJTggfPGYm7lUFmLYA9oM2k0JSS7l0ry8TfTfP6tMSl2IoSP
IoQHNpoNVmPPQMaAZCP0MXclTYrQ+Nf639NTnVYo2cglxoxBA3z3kcs66adpnPf0
8oMky2S0wdkzk4ZL8jWf8dzUslgr2eKQLe5hZO1W+sAn7kr+XR+s3c6uiNMprKX8
YKkckAqHTi69GCUNzie2MaLJem53oBqOFmu0+m7HxtBp18djStnckaboaU7baAKc
Vbr3nNHLHGXcoyNPm0/uamIKfDaIkzxK0tTkIfKmckl4882+XFbgv8lsLY+O/Ll2
vGQt/MUKJjsljLVOmJwjZ29rc70RZAWrUEt8VU8x27VGmm91rGCT78fMc0v0acl4
XHiGagKur4yE6WpERwCtGAvh1aF4kUQslDHmmjAqUqDw/n39FE33EhHdGZLEmblu
hwC4RKdSucL15bGb0xz4bzFRkYc+I4fpdlb4FHsXY3aEC0eIxEVswg7di6pkwsyy
yXpGENGt+DQ1+5xmQ30vf7bBQEXo1InhjEwMPEVRP/mXA0oJdqIggjkx8C6XVVp6
71x1kwCP+rGW4UVIXlhkI9CTxj5ZGa5vmIHchxZJ6HxiaLQ4OR60jRXCDGsdIv3Q
oW1vFpNu4wtz1pyZzcWwVihLo0xB+l1wMjBsitOKW9vk4h9gvL7Xo2LQhTmN5/Lj
Wzqiw51J2LsDG+tmT8nuVLGUhsz/RSbV0aFVGSRDmw+jYA0JSBmGeS7oN7yj882X
en2w+DPgmk2noGqHl56vrHGlP7MwiP8iqbeWGuodYexEFLLqWv6rlIt1V0IYiNKn
Yf1shrM256GYKGQyLz5EXytVHsWIhTamG4PK79S4FLpRkG/0ciJAQL2JVax3xbzh
CQ2cbkVAz0O6FN221bIZQAETXnE/Ywfqxn44I4rrDmPwfDzFKTOF5MmmrSeFGK7l
xTtexrVPBKkZlgcUxsVs3oyqljtJZDoUne0F07gXtk3OisLkEadPrghjLBrzK03M
4p8QoD3D9HNk+/RmZ8fn4KrAiBl34Y4i9oX0mKEsPO839p649XGaPc44P/grg7Tb
8TGwIsqMl/t5KS1wblDKkdyMPRSCrGLOHnSCBV5UQV7UGtWYdZPWFHmd3zZDBJQP
rVyzGonQDRggqjkQbV48p/vRdUDCTa58afuXSQfQe676NFEs83SejfVptLuTYPiH
DRsI/aJXFsb/VAVmxqPK3Mdav2vdbqBWKi1GNGNpebRjXsrWizX4R9ZS0ednKryj
y69kowRsX190YnG4gXaRjCkDhpNFrnFXScA7TqGKwa8LhJM4+dCcduqdrBTVqT72
vDcv9mPnSRK6NQ2CoTjRh2Epch0L+lKEG+Vm7uPupoW+kqYeB/qT/e6sOslZ7tPK
+YdfvfN0jF6I2e02w+YL4yVBBzzhcewY46vtEp12SFnAhTVA3pwLFHWz4Iqu94b6
Chl9ERj6CdpYPEEwtvq2gH0hEV/ELqiiU38aQTOeSXnSHexxQ/dNmogdnZYWlU37
Ad90GO5VT7ajB+WKTKbmevRTZL9xf5XwiVUv6wlTGhc7r68IY4GzJm3EbMTBIFAf
die29MSRQox9GoC97WlPtVzlDDniASwSLw0+BPMieGEOu7EuhMAIDjnykrPeOdTq
/FkBmJq6pq8Wt3zsNfYv8pver9wdAeZPFxAKO0D3a9J9srzugycdtF3lRG1lA7RP
5eXeSHaNGwzZaExRc0nRxdqoQCOM38unFT/e0Ur78UPrSa2bMRXZkVmAearGMeET
8Ofn0NpCSRa3M79q8lRQNK+AR1/7Oc6EfVk2zj8XyV5uoikas7jAJdnO3fRR8Ulq
RRRuE+EhVsnDFL7M7hjDfNgFsWRKC54MiT8SqfmQPFy7LGOqdGJ7/EOhiXbuhySd
kwEEBxS5HanR9uhp8SE4XLhHdhm/qvNSW7LXqszh+P49+H1MTzVq/RE8+FEM/8rv
P2gw2Bnyr07hOGJvqOzX37YqhoIZD8oOpjHlALB44j9cSroM8sVBjGGNvSN1fOzM
UTAaJsz185xruqX/+yvJRZ1sCffqp3tOCNBToqKG5tk=
`protect end_protected