`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
C322AjKOEq+k94hkAB74AtR+hRiX5ltWnE558kk+r2+AeJwVSXNa1+pFYfFasfHb+KckKbhZdLwS
fW8S02TnYQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ofzbFY7L06zQH12UEp8T9MQk32MkmgyM1pxnYEaMMkxVZT7qmkPcrHlezwtxvz50P7J+krNjLBvl
9WnXn7/AVK2e1kkdihNcD/4z+pWtcGzBZGGpjSR4cYoy264j4wSVdvBpkGSKWThPWbv7c/mnbW9A
FtDAWg+dMdA9gA8q5xU=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
IXMd9uE8RWu+CeYY914H5fGrv6wBgSGy7PE72qSrhvha977IgXL47aVz8iDNHhB7cPWaysiOfWe1
z44Ah2oDxeU9N/ACt4VELUAKFR66gxVBnP821bIV6lnEuGuDJl3Jt6TLksKBst+9iGTzA1Xbu8uw
awvd+dRvRdNaa6kB2gp1KE1bAYqbNMgDqNruZkGtFniASJW3xoeV1/4MY6Ke/rzlIV7+JMoBT0tI
DVQ7gnZUfCWyhBVbusKBJ6+UH1IGvBq18CzC6sx2IxEAvVuGRv5jTaSOssqFhs+hQyG9sUprjXLd
hxcLv3YYPrGUu2v60tYT+2heSMtU2rW3e31SzQ==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
gI5rNyG5c3drysVsOVroSrr4ZtWR1lsLBTZK0baFAq41KkpdWktaXW1nX/+2PBYQd2WuwEzYgR5A
3R9IbnThHfZMUVpTqmm3QCjUOIk8nTQkx6iS7xUYHB6IvuSSVzwXQYY/LqkXQLggQMmEXSMTtRg7
Ork1pXzde9DisVtwZ4c=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
bnYreZri/8cxBtUYrMOxeBRiusm7ZutmnARaEPgJr+swerZuyUOJZp6ItrV3CgROOAJPmjtZ5xM6
8p22vOpGw0kyktH6b/I7eW+xyPhz1bhIfjHoQkmjWC3hZnK7QT175CxgyM0a8/ioZcEqkVaKhUbE
nSPalwFiTDeR+NMIeZCpkb1Dre5ForqsAJpX8FI3X50m3/VkpVarXzYDZwRV0rJ2y1K/44VnyXVj
mQsPxaPSEaNs3ANT/XC25M5+aakN0smvIpd4uv/LSz31BvQiZAUA4Sadb8OP3AXdb7KKmDrq49oL
v0kfRFYGECoXJBlDZldG95v21lyt8fj5NUetxg==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
isiZwfumseLxHBLiIld+QGY4tmJ5ngxpWNiK8ApOc/PKzcdGQqiUXP+VgYMyH5NFXIvrL8Slv/Al
srKlPMKwyAl8QV612cY7tc3fHQsbKD5ebSpDKOBmvNA9WNpA5PTQRl5hXDd3GpUhPpxPVx+dfsVv
YxjZACjWp6636QxL1ZtwQk7em+pvgGpS0osL2Cxkq/x/Nu9nXN4mo9pBi0mWfdIbZsWy6Mdjzgx3
jW9wsPoJ1Ne/n2S2xFex9EgaCrfvH3v7tuVNaKtsd87nvF9atFT6vcr8VVLPnWW0lVCmY7U49TtM
KcqhgUB2Skt1rkmdS0rn2etqleC8vdiEnTMhsw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3504)
`protect data_block
54C0tOwBZ3FVAkNcRAZEHNUk5qN0ESwZd1RYHp+9lDBzx5AWif8VQq+WCnBo90hq2g8WR8QR5Vmn
xe8V3GwOK454IM3BWqE00U38+OCFL1jweLPsniDVZK9Z3KTqd0ea7+YlVCXLbww4JnXMbP1hJkrL
WO0lIT46UjM7Q6x3SaUoWDMvSU7mMrp8HIrpkAkJ7snPaQtJ8RE0SzaWCCngdgBx4GIrEPMvlpHQ
uuL0NuroA+Qsk8BJjJMtUHafSoM4TI49bJNTX4bkaqGSugL561F6magqUtvNXKk7mZ5Cu0oWZXbS
bUCn12xzvqIVqjM7XrWAFMHHHjHeFfoUKpHVLrans2L0Cdn11LYdO3CPSFfIFgejhsuaztDOznjK
x7HgtsO1LXOMiTH847OUhY428xby/XcCAylxKd5lJEUgNcioNja7MIWTxTwHGrpNgFs7mK8/pdyK
w0lD5TzNpB1Ko5IwEhm7Rw1EcFORYFx5PAjO7k1dthg/4aN5+/kKsikDhbCzLCeYrXAnBb45ieSk
x5+dDfn/77N8OkFpNAFLWNzb8ZCvYyD9NqnwjxZ6o6U/eSUKnpTfvYpajwqIkmhh7OU7Whjcol7U
Al8ro4apNy8HhPXzBwY0Fryx6r8kWs/rz4A9ovQbvMkW5IrynMUd6fPVxJISUin5MWcXlk5vpzqU
bMZVoQrrlRmeBILdX3x5bfYynHq0g2aAxSxrav13n8AhgEG7MPJlDWJYs5KU7iGLB8/YG64hj+SA
F73F3xxcQ+SbpRawJnYBt5gsfapZ8puU660wuE2VEx1T8lhdyaqYJFFYuV0Oa/Ygb4S9z6GeMcnC
RSfLzWUG+0cOo2/me8enRYRzpUUAIjWWAbtTIVRekx0ZEn02zpBucYMM3o+kqEeo1OEBYJqzYj32
5whb9n35utUN+Uw2EYqJNkby7/8Fo/XjMo0RE/7VcJ3R7rrghHvQ9gnOtXXdGuXuidJkxrbA3si9
Jkb4Q5dE16c7STXhNwOC5FZj0/6lOVQd4wCJ7TZpf7kJ0HFqxd7HyDpeuszp2qQXNcJwgDu7dQmC
m2kWNO4VA4lh1t8lxGvjUcnGaH15a/s9lfZch0sRZK/umAuNhalfOg/1l48Zy9os5AuAeYbyEK/j
Mz6wu4aQfwHN1ZaUkdnmMHHQMSGWxHmudiMb8X8Un3maCC8YTLOzN0iC7zZp06PYvWbiILWEBil5
TXJ6UUdUx9nHvBSENDCFPfNvK8JyKwCFg+0CrS6+NpffKw5Y55oQY1nq7t+F0m1+aw3XrtmWfCSX
7EH3GuI1+k5G2HO7rjaDL35A1ky3kAFmSgWFMFzz9MTMK6HS2akibKkkjnCzNnKDEx0z6X38n9Df
z9k+sSh+ZOHyB3Y24vW0CCAtmBB1ZmNE0K9bU2sLUF+iXdIEClvqQL6wTx3+XPtehzladQhV+7AU
2IcnUskHViwAJFCeGH6HDgK4EjZL8HAw1WHCfsP4fSYH2hBXhBsP9aV9lUXXvWyoPGYOASMQSqIk
mWHGmPhM+Xy6JxYKpIe9q+5HxQR34ZxXJbX8DtoVmxNiqPk7s9+mYekIK0anIDiT/PkfS2hiqKx0
ho+/hKvsoJsubA8JI63Ev5YnkWinNVqz5iWjqE9f7WSI1DhYQTyjics4+Vse8K/Hb/ynCyndaqaf
/SkY/5SKzoAJ04VMJAVoexghs8WqBdD80QUyBwkECu1HoMwRz8jI809YwXW8nV1mDZMsX/LhjQiP
O0qRsk2eG21PsCQY9iSG2jL5f6K+XOeKfkzlhENtzoNCARf3qqaOYo21vv9LOK74oB7ZyFHbU/9j
FZP+rHT3ZRo/RzF/y+S9fsU1rR6r3WxirqIjSJVNrCIHSTE61Mg90eEJjYbXbC3uQP86XYWowFcZ
VeEqQ9wqK0Z+mCNFhLlciRup/9ZjVorYUcESe8gujVihveaeQqW+wUDhS4gDFyJ78sG6h7Sx0lWz
EaqW/waYoq979E3k0h6a2GHJdGn2ji8s1cpvzkvaBOzGalQI6UpXFgzYJ2mXZkZfaPWZ6f9GYXS/
3indeJUBtmiIwSNP5Aawa1RAsPXJpf/4miPvcyfO6JUQVrgeOpFFFABx6JDuCkj88aHBmsb+CxMd
wujtIrp3z4tzPNSZbGqXu2KGyk7zMbr+pj+LsEwwsdi5isrLifbNgLblRHnaZ0WoljHzGPnXTgzX
YHvIsJ+5Sch8B4jllFGl4x8husOx97k2uFpXaWf790bBVrVGRxDipcftSgbIRwi0zdeKGEefsq6J
dDYro5Why9bhvuNV7a4C4FPXFgrfXxMo+w+OrqhCmUd6uAK8X7sYgDLaczLoWVNsaIQ5kA1JGxgO
fVFSXyhz6p9X+8IMRuaYW9St0FDINYugyCs2Qu8v1JdAqrndVh3VikSHAhw6jWuWmhco+1sS19Ac
iKXiPlr3F1BjLQ5fEMaM5/CEDW8mg6GXHGl32wNzRsMkcZ/5MLC9df5KRva/z5EzMW2IQ1x46oIz
zlXtI+QHHzCpKUpgVw9Y64gjU128AW6t+TzGUboFP8ggArHLNRa4XA5j5xclxoWaTXO+ulHTUPYr
yvQYTtK0aBs33JcvNlyGp0TnohWQksruHTIKd+NW6BGXA9rbRFEdfKqZ78gvGaM+Qpggt7UINyFr
JWW8Ka/dlYTbiInw5iU5b4ec8gsjQ0P75Zm6UFMCj4rbzrJW/hYPWnr0QSUJSjERLzbNvlF4Zjrd
w+QFRuCN2srqZm+x/hijErJ3d97svxhYGCDBaW75ijAqYcezg/LR2ahG2qABcWIyA3DLHNKi49oG
FzfbtR5Z2rm/uo7JrsL1BNYYjoa8fnkbqTJwI1ou9uao06BpJGOOh5eywAQwzYd+1rUIx+6r+plg
vVENaSrz525RgGn07emHEQ9TTRNTUmxen9wn/qMD912XYOX0HHQN7doY9fJP+8YP/2wcHQXbuWqM
iK4QtSymapHMVlICX/fNhe+fv2rZDpzis+rEVXQlmgLNgsogTOwE5ARavdlMxNxKul4LP+Ul0WC5
LmCXHUR+hRyyjCZV7pTdbQ3QuOYtoyyoI32Y/1Fun6t1DtQoodDBRgcMNbxlDPbzGOfQO8/piok/
VjII95k4qJ2sJ620Om6v33O5osrq42vmhQBHMg+LN9H6hjfYiqgK/OKh0BicllA9J0IWqbgtvvx0
cBvUC2iAMKn6q6zm0iEGAzVwWxofmBkym9xT3WsYc6U5f8UP3DQ+3Awx70xJG4reAVjPJRddFRaJ
ciXTaZfZoIlPplTf7vAfN3TziWSFs6fxusxndIal7ptu82Vh8rNtPtfASh2hE2wISYYkERKnobq4
JQDb0o2tu8GJQq52PodYiReYWCn4dnAXc+DgjIc/LvPhT7APbPjE7JHhleFoP0/4R6XlKrbvon56
PLPl7M8m2TD97azt5JilGJZb5chs/sY2xBw/pkaJsDjtoE88A/6ybVeUhfndG2ugRM/B5lgBDBf7
93m6oUQRzBA86eyTXjume8Y4CK605A+GsAMR6QoqCnuJk26UXAMRqPtHI/qQukIQxK+MqAOvPMHX
EdteRggtgZrjxVDifjsRa9g2nWvi/cYAi7qMOhCXvUPzL01yQ5PApT5pZbh08gzaiiq+lPAw1Ghb
lxYT9Db1URy5BA3RfsZFjjXV/x9zNGuPEgGUgh/A6TLr3Ei4ep2EaifpVVgBIfYYmDao0cNUYMaw
Pq8VheNdYdOBv44RTi6PUsZlJWEyIVgHOpZt5OxbCDHfN2+An36eLIjwasiUtAsk+YdwkqNg1eLl
vK41cRRmmlH7FlY7WbHjlT+FH6d4TB6LyjkiP9w1Saxda+bd2XXt2P+Ppf1KaXZ9jl3oz9uVvjZF
xZZ6MNiIpVdmHnnZslrBLYH+7r1wbpk6h1k6asGzPfkVXzevbjznpRM7t++cuUZZJVzf0twHrB9X
TAWeLoC5jsIncYU0eTgPi4QJRS6k4xBMKf+hEvQNJHxtTCfl1NbCyOUM4O8fDwHEgREn4H1z7UGn
MvvjznNRmXwc6YAqmW70l3mfAV7jwuuQrilIWn6dQiNYM5ItABIdpntyi3CYKuWDgmr3eitmKQzI
jjz7RCH2r20uaawyOoDHhwBAgX5UVuXwk+BXn2Xv91VHnXjDr7yKRpdf8n9gtk9mw8UDPf88h9B0
x+9c0wttncKysHZQot0p38fwvPkL3U0Dar/pZxQK8tzqe2jqcGrCrpCJM8RDX6tgWN7A4gyb4ZdH
lZE5msncgcFVfIiTEHLwlfOfzAzwkSy4zJ/ut5C2oie0Rd4x86Il+VPDGrrSw4YjgfXcPW5J2pFk
p52xakMMlXSSXi5WDhnvXZ67tqOjCAYv4tYw75Dn3lyByUmWWy2ABCXXHaHXZrc93iNW6x/ERFe+
FqrVBDVmt0+CvzOR/PrtZx3Y+2jJE7/UZmO6kiA506r1itVGT+UP7n3OkFcSLzVvg6xbdM3XNKYQ
A8PQU7kYsAkLljBg4ZFtPJmHSuzHFWfm80owontPUWe3SOFSXxSms+15e0PdKX/YLtU0K6CNswfO
3GKsynbUO3zmaCa72UzNuJgqkvbyLR3Oj5A3rXsWFPt6seIQGrI+X7Nm1+8D1Cj54nnQVQbPNdiQ
mkLCWhI7f3YHu4j/ReYa+/XySTijO8oDZTpl
`protect end_protected
