`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 23952 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/9huKRhRMtvnNqb3Z+UU7TahEoHV+T8U3P3ufru7l1O
3DlgtZzb9QxCbOjthp9+wDkjygH0eUfDrEl1ovhZG60o1iDkEMnY8q7HfLjEqAP4
9MMI6FkLy8yAmodKSVmjZgs9+5Uf/xHOapKMJLL9LmIrQOKSrN89VKY/S9XA/0Jy
KK776Nl6MMYaqOmYUXUZOe4KHJcH+z9cNlwNDB3R1kwJGKI3TK3BcmPIpuVXXlNa
2yt6M0F5HGclIcJwsC+cYn5Tz4lGAIR2rCcCPpVR/m1a0MQTyvu2SvO8hcSEJ9qY
XDAMFJllOgrktGoElq+tR20gKnq/jdEXf6mGVmywXeA3qIJj+kfujOmZkyHbmGg8
cHGq2cadKImItf4bvQN6n6V0pnQxMiqrQJgA3F0UU49kUyJyIs+kBNnsKKajWpi6
UJ3meI5evtDvhjS/uimNc4x5kwFGaQsXEgzjlnx6W2nJhJpO1IqOfWaOGQ+RvFPz
YdFoyU+UF27XjkRvD722LGK+LIJSdrbh4ciFw53g5o5LwAXF47Hzd3qcNird9FV4
0//9ryOHJ0slWafgvXwKssRMbMfqi/otNK4OdSuqQd1zoUZnIMtWyQBXyaYvNKz2
PSRIchYhVDV0xa+rCntLZk/XXOSerzawVRJlDBP9rlTEMeFMsCZFvkOzPeHxnyfC
W6dvUxHU3Hjgwt21rzcd+IRCXwcWb0kt7q/czn0kgQ8tXEIWAJlgt7oY3tMVXtm3
v+Y/sA+ddt310soIBMcYgoPlbqDymwYNII1XLJMA6oDOGcBUcodPi3LHMfJUgunl
KZOOXLWQsyv9AgT17TalRaOvZNHLVnDDlfhD0U3XVz2SwhrfbPoiaRs10ixtZOoY
E0151KFqeCkiCnCmdlnHbunXlbbCHkKZ7Z5hCK/eY+NjHatDyPdUAqvzK0Q4UfXl
xjhCiszHtu1DIprYzUDaKGqp0LP6Z4AQ6rxDb/KxHPM2k1Li832Y8FQJdOlID3tQ
/Nydjp1ARI7fEm0emBA3YQoc/cuLF139VNrivLDHrMFcPiKq4vjsflgRHEWIxf8J
VxO9XkZjBJY4TchCf7+GK+S/NKy3BCLflT73y+O8rvYbSY5g0D+L+5/jg86hwg9F
HtqDeoSnaI1+qt2VARN+RXpZigLOTQJOXPJV36mLVo1CSRwffB5lfVaow6JpXY7k
/Ki+8ePjm73Z7aE6IHjjET+U03O8LKl3tYSIX+cUSxHD+XmCDEyGD8X1AWyPEeav
Nuh46IAAgRKfsgxU4/VQrePq31XlJUf7V4Qq4d1Zw88Y5FcIDRj0l/gf7JNJ49EH
3gkAar32NUg25UPEnR2BQXyHJxpg4bz+GnXiamTeRaKa6bIkfMJqEZ7a1aoNNj2+
4kb03BihSPUZBKwarRn3BzZpGKTfYPsYsDJM4I8ZyDK2Y1xCe5e8b86aWT8nVMQ3
JsmVO3v3wV+N/jKJuMBzf1eg7htg2ZpPddZuRxvG32g688wuJm6R/NFBLkpLb6hU
bCEdrpc8npObmxUJ8n4+s0oEs7mBR+oPsaH72zMG0PEfbvHq11y4BDqBSoLVEdYB
AxNL3txgnkl25q0/oniLJZZOpfyjfEPaFXd/hedCaswqxY3Fct4MFOyv+lDY+ol6
wauUA+vg/wfPWI6M3QgnAKAXUc7UcfnNZ4Md1p9pfMXqRd0ZiqJIckVZkFjts//F
f5+wQowCe2tkAJ00NrysgqcXcVUp7KVVwbAE+kPHKryLFVuNvBVbNYfBwzS9J/cu
l+mnj403cFjrMMMi+y08krUXeomWwZWzJEUJlFy+7/Z0kwWORP53tQFQmF90CCus
TEwzqYt2Gjk5SNWkt1shBKw6KhfplCOLapsdbwe5D1NO3j5oukVc1MMFVpJELFF6
Mc/Zf9ZZ0wYMi2duUKEPXu4U2R0TYnuZbZAvX3oiYZ5WA2XRtul12hJ6KU1b0NQk
QXUknOlLI3J4+/Zj5Sg2Ff3e0JOs/tfsWxQjMfkXHN80wKg/ZVbU2CksJzSZK8pE
CvgGmF1ZJUbCFNE9+T4qTcGrw58hbHEY1BNRp3outd4/MhA81B8ClkWQedR0DDBX
DEDwNiFgd6Sk0EpvvohWKOTgU0P01OQemFyNaJIg9sdrGx2jYeiLgMJIWMbLzWvO
XvEuKtEbqhg+IvfkfLWZmr6KqgIPHtutfyFSV2n9cDj/CDC3hOQHPVsqOrlO9KR5
rTluqV+HmXaguf3O19+WcG9b3W5XOEoWEm59Ro1C+w8pNwV/XX8bn2BNxzlKw0H5
bTQKpUBqG6FKH73YrTWuGDb5CPM6DHPayqHoj44koEtVvZytXWfus9Ax+IrAlmFR
xh8geS9YBEFdEVs6hVQjx5g01hukxzL3jFcYINlpAnm1ou6D7E3LhfzlScrnDDxa
tFghKIkn7B7Dad9acDoU7qu/MRK6sFDuELX5I2R915f5byTBT1CwXf4l/+CNR8Lk
1gA4f10ryg8FRIJjl71Epk7j1A/BXZZrZGPSNUMvizaM6fO9Ad70ONPygN3xxkjw
f3S6ybhcQGHdpFBfLPCwJC8VAqA7nJXBNo7fZb12oi4AYUUxFGzGmPrctjKWgNPd
zHpa8a5F154V3Y+d7Mw+TZLaTSehH9aCSeZ6hNn25r3U+sq1cqy6udXfg32PjBRI
w0N95Zcmvme04Ki4tECqk8neY5kgfMOergsW8ExctsGePtuouRtl0LBYwiHYpgl0
OsCU+E1vq8rUGlX2372KBqkdrRJPAaaEy8o7rlfou/t8fdFVQjBC5zfWgBuma6GH
smZ8L/Nlu4pvLLZnVVTuEJwMgvljrBiUJkAGACBzir0NnUMH9XJqQwAIAiWV5jiW
2TVrV5oAoaX1ohbi+kV3oaNkTbZonhGR+ilsOSkyYaIJ/C6m2koP4+J4Yqo/FpxV
9REn/M9nTKbSBjzcqya74spWlroMZfLtEJwkn/xus680zkUbZQxK+nhAZj54Xms1
hT0/sJjh29ZS+nFT054pMb1TsS6hDoNqjOl61WDGugREjKosla/5kFy8FiPPSGcA
u41hNMpfDxZvXG0SSBgHeAMp7SP4AJsRQy91OGeDteMaiysYGmCd3N7EbPtame7d
9w1iUbykldqzmZauZVqwjSsiHu21zsRFYkJBb/a4rPwMtHhFbT4Ic1AA6uqPUn8e
rp431wTBRBfvVY7lzIzR/Ni26OHvc1Na9oUr+GM7Lj7iiiNZbktaHlcqF0kdNuND
oEtW3y5ay/IfSnGuILzj6BsOX8YIorpfpnRWy7npDq13geFITTajlKgsJ8ruY7np
t9b/8mgNueFYGCruXfN0AicmQeq2g9fuT47TzGS8Ezb5CvwFiLJb5Ar5cPUleMcm
VdJDVNy1H8QePU4drzy12s4xWA9j04TGf2L9B3t/PpunYT3kvvY0tAG2TvSpXJi4
mVxjWY43QMbM6wWM7M3oHzXQi6zz9mpSdDNuX9fK8Sq9jmnWo3tCfynjMQEw1IBx
h06xlcLvFdvsza/q587bpQONhItkeeKdoLXdP5GBQ17RmYGSLreIu+tKHbWbEDm1
3dsAHHE6dAaAGF2RMuwhvhQB1ezQ2xNMmWzRO+Rz/kAYROY0VEfxhVF8IFY3z6J4
X7pUn+Kecg6Wao5eXaDo/4qGx98oEKwS8DPqBYr2lYfTElAzb7/gRJQLwDH+TJzI
T2tBsI8Oqs3vpMIz5qyE+cIZv4mFK9fa5lKlH6PgTDQpEUlsVwXeHKQg+bYGdfPB
ofGWUVq2J24WotqLpIMy1mzND6eG2EnGbdC0g026dK5CPLirlldG0uLWkkGgzIq/
xmWKRbGGpizMZ897eg3QBZjN2ylzpj6BGzLD6BeJz9DA7+cLEGqLuG+A+ftx2ym0
dauqOVN5OmEdV6MQ/ii3w8LKDhhco84g/LfdibKVNQMNA44RgJChH8fCdjxobxM/
nWC7xcA3dJ4gxIZTTGCz0YuHbBcVQ3Y4ecFgDz/LeRmtBVfloLtBb3n+IUBSKRIf
0NsgvXjRBn67bS3v9fPKx//zyE/4uFEhaHiu+cBUTUaSF7frk5CyC8J/IdQ4zQIA
mZHmzb1kOZUjCvP3BrEMHl3cQXqv5pUgMCrfmVzTj1dHrqQVxW3uW6yqFiqb2Ima
CCFa4BL3mwTVzyelxtxoDM0plv4LZu9Y/Q+qiP5vz8PtnDdJBaZ2H4nnAR5CHLvm
Tbf3pLAWSYoAAzkg7WZCE50qLmP7rkRPQX1rJA3IHp1R/caYKkUFKN9Lg5TDgqvG
TECTDq1pFfEXD2TLTgfBFD+DLKEENS702vg0def6BQO47kHLOyUqWCFvfflmUIMF
zblAD9HSTG+eHs71tsm5osK1tMkXdKKN3JI8iKE+L8eTrRjbjIcuCd4XIpd5s88J
IUV7puEMkAJOHU7pIItn1nx/8Z7aaHRqrC4Yq0PLMIqBdX0gQY/+jXscSomCjReE
jz0LLzRLQaMfoHBAbHlLhMTw3iPnvFcOsyKnyZUQVBSQNjNEE48yGeHSrBuW54WZ
9lNnoStKyB0TG/xMOGHbO0CUfr/zT9O4PhKyrd+o2hHLUjgxMWk9rvnpLm5qwQlO
YLlrEwQqBMouftsDQUTRQUcKG5e/nyyg91jtuSeG8dkrDsC99xresMKkFiY6ag8N
lDefpki8Bti7f+zqaOqLSP5yoUdGoODLgnnzOVF98+kWY9nv3NIdrWza7A8DKY0L
+TGzbJfwsdgeFOZsNICm0/BnBaxl0H9LbOtJNl7T+7roXOjgOm1sEa8/xOmS9Age
2StaSi7p1kv3YTfdML9eh1BEsqHCx/UBCQ5P0Dt3pxm9XkabOK1YEF6vyFc+OvFm
SmDi/xcf4dlvibPVfXulCPhtKldio7DMyvtKB8IGvbSm2NyWtRIe7n/mwfaHTxCy
J0s8ewbY+fsrbsfAKPhT/I4KQFcFs4NkmZkrB79Nye+EO/TwSjKvp3NIVincMrou
jcJRvZc8Hqc1q7HBnbtMV5XpM4WPA0Q4PBp0YuYA/YNxa/7TKTV4QxRGZifA/ubl
DafUS/AIu0FpcIAIW00db57DFbUc1+AlOSHKYGzGE5+NJGmPk8X5B1Ur+GTvT5wD
aBLjh2dd+3O73nBcB3DhrSCrygn0rvG5zt6jJh75nL7UchvZhTi8IRrZyC5nGK33
KqHtQecWXGLim1f3Ftzzfa3ouB/ifyapXI+3f8iHpGtf9XFoYgkOVAyoPRME5qUY
TX4cMmHBxmWj4X9svEjbpOPvmjMR931DaXcLwsXiZgzoIhQvs7yq5q+ShLn+n8Zv
of6LAoJoexCQX9+NR0W2eH422ggiSfwM8cz1D9PrCkM3+ZuTPnmAwcMyQm7SGg8e
1FraXjhGDZjYul5Q5+7fXfydd6w7zMrIIOnkdOe3sWw528G2gSSZLkm9uLijQHZE
BqAT5dSUcjpVrk+SZGBSL6YnmnUmxwXnsyc6Db+8umKaF/6f7H9d5xd4IJfu5hcn
QyNVkKab49IRwUoeo97O6Lk63VPyDsakOxJvzHFyC7yJJmdedBczz1HQ/MA7O3b8
M0JF4AXtqqH7wVgf0gD8GBBZk4ATkdo6NT3+ke00CPQkFcodtOYuSclms0CV9koa
AOYtHVjuzJRUecvRFZkkoijZIyTr6gcK8M9XJLY6cLGr866x0fLyp+7sF4X6KETJ
opmQyBTL1n6/82cPM8IEhE4kw+aiblVazxTIGmsEtsFpM9I4JBqM3+Q+xRM1cVAG
7JNMhWfeJ3B/OBR63vCXNrW6mGm0rMwGDqxx3J53QZqJ/8mWc5Xy/RuMpeIcFuRX
5RvDpVjNJ4Hyunf0vbXn6qoySZkI6sZn/auvUzRAVsPdOwx7IrdWsPyr21jmL1Lg
j+NeMCqablZtB1Ahhugajqz1IR6QBHEuECDno7V7seXZBWlv+XTGCwSChzHhSwUs
dr4JX8yLVyQTeOF0/r1IqlpO2GoCtEAPJjyx43dO7CnN8SwXoP3FFAfg9UhAQy+0
pjD/5PuaQstKk766C42KWUpNqoDYH3bF7baOTtqEY7G0s6tUVef30WaSCqmGfGOB
QWahRQeXLLTSzGnyubwatFQVQLWikXqnq4S2r0xYwtJ65xY/O2A+qXXDyym30UNG
MXfK3xhleJxAlEaCi2BOUUjVLm17aO2bTTRrL97Inirq83t9TTXap1W1RK6Mycws
rV78LNUWRZR51EYWfQdC/ZiRS+saSMYy0o2PV4EhluG1U3V4p21I/JJk6j515/Io
tCqiHpoluAn/whT7BZ9AFAF9RYSi5mPGPhQ8XT9bsr8nEP7jbMVI7bk3bANap937
YIeRPJ96Vm630l4VzN9TQ5xfJiS73hciOEUiPx/Zjy89QG+WP5CbXlwDMQqe1dYc
jwoMMGekFK9XqD+En9Uj750WuNnoCQQU5Mf1IIDmh5TZcQussiUpYO+TlrV5j3l9
ZN/lfmqh03cacJkjhQ+Kxnj12mVQ7debDUzbjYOQKGgHg7laqkKEwWJt99H82aPZ
5vBUQL0PSVOlnBGGzw4x2r0RVsfJgcGjiy/Mz7vC9btqz0awWw+v7t/Rn4uPMurW
MHKEWwXh22ZQ33ERuXrW6sq847Ys8vc36M+aFe6QBX81un+VKQbKaZnexrG7CpW9
TW0vjqSIUOdbsu2bVlcBdNstpvO4IEG9qIO3nQMggxarhcsejTboHY7ESlnPM1+N
7qixBD/x7r/cNTKBFX+HfhLMH+YHWz2JFTK80BhEBiE7IvNDW7EZOpozgzuTXDJO
d3tNrxmuoMFSlBpNDbuBq+rSwpqaCN4ygJXyH5OBA6yO5O/Nm5XqK1JNvfc8Em2m
ybiY0o/OGOtAGbNqYqxtKSXGERBb95c/7AQeCsh8EParGFz4CWUbKnPML+upV7Je
6R5XQI3Tk10zmbwQiIUB11SDKZE6WwBrquFvHoaO/XhtJ/sNZA6dU2vBXgkGy1Y8
hg2ywu6HneK5OyTizfm+bAQyOI3cY6j25QxT1rCIH9BchoVadPVhHkYsVXGX1uh/
2P8CkGkGHphmRAs1HofvSQ/sdkFOu+fmaIDDsJfYTmIGE6kRRx+azLih/tH4W/ry
Tp53XT2JcygkoIE9eiCD71BZb59LnJKssKqzqy3nPFzuTah9BxOUY60ftuVubFzZ
9RMoM1FAtm5pUr8xDTE1A6V6r4GDw7y99JJaPT+Hasv7q0EinBauGUuEgni9ace7
quj6CAypWKOtvI7Z4KRyoNiTJFmNz6PluM/LRwOoJC60TKKBfbMRYZWgqCCuVs/t
JtllaoCEOXV4qEuI+WFF2DmBn8s7hDXZZ39u1aZHcccjXQFDfJJM4oVlD3MlKuvF
F7m/fdpNULU0JIurbxLC/WDeU9eFRiXR9nn+HbHoISL0kkf9EVgb6AAHRdMAVVAX
zpLkuFCOXIY0N3qh80AZCkM9lgkUWT2HtL7oXgBKCldsTrUf0ZvQr3sf5fCMTVII
jjKnORS20xKRKTy7hDMNUyOIYc9Mxo2xyF9/qETONA4VeT5oWfyC9K6HKcalirmH
HXExWgzuzRzN5RbzQSR0EeQAki31okTMBwEuC+NO7mmX9Wbc0b9XGWdnE16RUzs1
zoqGN+1wIks8xYorPIfVUhcmNxHODMjL5rfoGavmBBFQtvcL6S/r2Jtsi2uI5n4S
bFqtu/riWKkCUAYHbB8u8pgCNkWOQ2/BR+crrb0tEAGha7pyCFi01aF8mqSGmmL+
HA7rGAF566Y8F7dIfXgIu34aCsRWtaRMB5lRyX1EVfZPg6c2qt15fpK+OJaEonj3
x7uUDjufmRuCfmzj4Cxl6eXBzPRR9VZYqaX2q3ipNrBla5v/LflzIAmZMYE5SJol
iot2hAxYVn0ZEaG7cbVLNT3753NcoapcUUDPyTiUuO4mNYBo4yFetR5qZkGP51yq
P+cgHxV1/ETOuFh5V5FtWFHWkU3eNIRuTxDJubEPq26mvnXZcmB9sJLZ4ElJFexT
GyJgBLo8auyt5hjqxH378MtKbpxhbFgLUpna7YYK0RFJPbus2WYXEk3AVYGV1w4u
u9YtPoMoVFuqManErHbKb8tS16D/ohvO26w7JJNlm6+LFnEaLaqVcchfApXXCRYx
Kh/gR9QJZ1FJJB8y7LPK+omImFit28z3LTUVSkCBx6+eU4OJ1jzbNOT0MhefbglA
xh+dd1Iiwgg275R+34Y0ijmYJ7WOQk5Yu/XXVmV5bHvuUZJfsbUsouHJTIcwmGV0
RCylCWagKC2QcZFCuo+naFQ/0juEmxpmaLCWJNLm0WGHC3TFv/9Bh6b+cT0iahiG
ftpPhh0MShZC/Zp9CyjmRhIAIUybG/YH9EH2KjkCd+8OJi/rEnEny76lGp72OuiS
pS1NUoaj0anOGNHFlSs/tByXlDs/NEvI3Llr61YpmW3kIP6e2/8LEf38mfKZXUcF
vUVS2Pnzhn1TnQLTxqda6W6TgK+oxl8ePxpA20qAx9WmTOD4lFkx/eutunSAOggF
ONR62JmtyfvtSipUMZqS2hkz7kvd6oZ5HCxgCvZtYH/H+Of8vIQEUul+lQ3DFbBI
M47EIrv2XI/qtnmakMxaE64k4IxVcE19xLCjsai+CF9MI6cGl64JYeHRwQQodAMG
BrgNOdeOAPRITi7H9MT2xDkPQXaO1KLcMwrIt8fwYZawhUBuTp/su4V+uQ5vpT7x
3y+yDgBD7bE9GP8K1u/6Q3deooUsxIuvJzJaQzHryd4N1g9xz6pE7MoXdFVf9arj
SSx2+MquCsbsSD5Xp/szfgwiyLN1tF+Z0LwWW+PUuUL1PLD6KdzIJKHKKDQ6iMKS
N+K2sdR3x9vEPt+ZQ5uO12zdpJQ/9Zz4Hgw/eSSlULY80SN9QGFy1zosHz4CJ3mv
L2untbbdWDaIP5KtmOJ8PsPzv6Enpb49mvcEetnkD31R1twgxA6A+4uM/St3VLWc
bbA0KOY4PmJpw9CtjWmIzU6KVvQ21L279MvZJqxpU4PRBOIN4adcgYoyIwYsES+l
QGyCojzEpVESE1SWWxQN7AboNbeD6u9bf6VDqM8oaLwFWWPqU+iclHAWm4bT053B
9ClF1N29xbs486lJoy3JDABkXsbibhJRYD7m0SZYx6NuXRTpej45I53VzfM/aUJE
uXPKaCLedplnuIE0USQ4wo9sJuV5zODCDRaq1qmfba51J7DlLnn6/UbbJ2Mjo2eb
jZBHlK6u185B2xfxsuDRVZk1JN6cT/9wPRqcIUNK9SMFpBvuOi2PLzJrXzyY7o6n
JVnSt21QktudS3grt8Yac4mYHsxW8YUQUq0hZysUNszrO4rY5zu8iEwaddQ5hte2
Pw9DpfexJRmeFSQKA2D2p1PIUsE4mu2EdTadmO+k7iN02XDV260hxe5YHR+dLk0C
3o7Wac7W64wSiyQ4mdwf8pCryXZyKaPi6+8bbuqNYZIivBfQ/LsCXR5j+1dZAI7t
H+xViB2aFVhHtb5aFrHBmPC3f5Fz9AgIu4fqpApUzpE1pvZEA+5M2HsqJogtGiM2
AeaDsk/MkCGC+jj3kcA1dfvs4WGIxXRwEkfk1aAI4hD/BilgTt0ecbkHb3A9Uvgo
1daVA1idWFcnwhlFY69yk/8lCMwh2UceWAUxPNbjCxodlQoctIOTVyYIyG/mq+rl
9WA2OlOD2kzrVwSRLk4vDIZ0tlJi4Xl0/lIb3O3Gg0jSBUGVO9onWDMlCmbN0cy6
rJkNXVeSd2prCXPhREQ8B/U34DwhG2MZk5HzUgUOekx+5eni8vpaRsOa+iXSFbq6
KTT12tK2Vjv69Vn259blcK4o34jDg/+1vOWokICO39+Q+1WIWujwyQGcX7j+Bt04
h3fyhUkmbTsrIT/8vxbjPMRT4eGmFa/lAYoljG7E9OXAhjIU5MNQbjCUlDrZfaoQ
qNxfqyAHYmOVjyF7hpHqJZ5ADaVNWsdxBzFdDYPdsYgacV7t1Lm/5ul2z+VF7ko3
ZzWmLqXbSBeeDSQR+8VWul1W/MT6A0VLGlteBEDS09g8pbnQwaicB8AbQUiCfnnF
3eFof+vif5CLLSq4LSXTMTGVuVdFlSq61yajF0i8PEt1RM7h0/hvMXw1eJO8gibE
OBcr9FF8kBZODqhCSgvD1khOqkkqxicghvuENUzFsy4nWWsIS2fuQDBURkBKBK8H
aKnx3mz3Mb9ADRVT4zlgBKHlxF+wiIQiN9OlYNUAnyhrN7CUL/c5ZD6QL0dz/ELj
VfV8OcyM+R8FyIgn3wXXNJGhCXLc+3Ehtj8P8iB6W2KRnjMm8lhfktglu9HXDhIT
ctzz8zgBESdA9/1Zo4BwPySKhJwg64PeQiPPzgOJsRYo4btjQg/hIK/r6ASN0ApH
jcHo1aaEhcy8z13etwSNpO4vNOa0bUieC/JAqW6JG80v1M+BMdMu6pITxoZp6Ubd
sg17xYdvh8O/OEEB+IHok1CnB3PnVGVn0iVtC/Th25ezuUYrYMdfG+J7TuvOwFLn
NwQqD2s4VrbIpImW6AjdwFSYtZLlhKQ+E5KuE4zxK9E52atfMfqAahb2SNL37Xoj
HSExx1WdWticOML8ItTT5Lo7j/2hWmXoVmuhXxJXpv1nzwp1zFo/9Kr3472BGa8V
KwrZw/IsxkSNUayGQ0y+fv9hZTZJyeHlrweOLnU4ZG+nCBbhJHUentOjprIlx9wr
9n0fzzrkIqVA4L6gfk4tNMjZt+PkhYonmXD5Fev0DluobLF2JZ0iua/CarmoNEIv
DT1q488E+8vK65IkDywKIUgsZZG6QIrMNAzqhjtG1obF2eGgX8S2S5njwv65p8sZ
KxIU9TGj0gADUqgceRu0W0zoAJK8lO0bGokVyWcht4ffvOFdQWb0N0uZXgmIGOqE
1zUBkrX6wS5UdtOAKz1zxk+IrHAnVo0IndupsDhbAOUR6C9oISbpqrWn/fO2VDSO
Hp9WvGtHdIgIRoOY8SuWWjRCabMExb4+2F5uGEFqniN/pdPRL6twKTAX6alfreB5
+yYc9cuZmrDMr8exjoIPPfN7FgOv6nBd0Qr2EdDNRmd29709Glm2gu8+okRpdwyl
EoT1eVIuQs+9+17k/65ShdSRCvt83sd3L+BYbqCIpbQs8in5JQbVm8MoWcacE11I
+gI1rhg0o+zerHmnWVXh9DAJBEb6pPfWefbJm2PfatAnoc2rljME+quazzIZnaNJ
jpNGwtJDTwGm+CzhCkK/7gQ1qB0r+taINNuqwhXcLKrCKcCaq04/V/WrwZB4mNtP
iqvUyo9rh62Lzp+VRRnDzPtEYQBARreSzGu2h6ngu2JFz0M5emxd8FhR31SxS2Bg
0LFtZkN2kRdjI916QT0Wd7Kz3Gdf7fEmxc9Cxc47Oe8gwhhMSIZQiDF63Pu3TYl2
sLjTTNn+agcV1fXDbd6r+/+aVNXWaPSYHqwDIX2UivAxDBIvdHiLHP0wH0JRbReX
B6O6zxrYQQvKpnzrSk26ljScBAt2TbGEYIQFY9k05cprvstHdc7hzfOCdOFzQ17e
fHnskBGbE4CCCEaOzh21UnB5sGWQHGW8dI6CXPbaR6hIxSL+o6Ot+vJDTbSPR2MW
YBujMozvM0VG0CiZBPD8S1kvoKs8mOWDODJh4T59LVaV0djRNX4kaEK7MAIDyhjU
tbpbXfJUMRUap1D6JvDrNNGWpfJ8UIHqg7QWx3ybBhd3D6zTJO452P6p2R3T6htN
uvJPTKAPoo5GpaoDj5TreL/uId9iaJ/aQP5BFjV9jsgBXmy4iFGqqSbQYVSUDKHM
9ma4cvGYAX/0MEZ9U2IqhbFW5eg71MyOb6dyj8v4Mwn/5izY8sHGsmRiebRzPjoz
aqDRLfA4mJAc6KooxKOOulCIjjZTb89gOD5WXKvqImgi9U3gRGFBsU3tMdN8tyOu
oK6To2Rpx75OoJduDxFxZbynrGqVgMF1sPtNasjz3rrgG3F+85zOTE/lkGAxAaBC
i1o667+laEx81k2SNYzQ6tN+nK+j8gPyoJED7xHf23TgaQExwRYaezqkWzgFGbVr
8qklvwLnG8AH2rHYBUBm3SgcBuKTZV4suAqWg0Csc3Lzp7p5xavWbaXnpfQ2yGfR
16vhP+TBm3mOHM9A3pPF9T/hkKfI9InmWAEjvevwdv5eTvKvUK7qQGmMuYuWZcAx
jTWLnRUiQSS3D6C5sr+2ePI3BnCntJdIhBzSRzzSVRh5SKh04BSATmNai8K+0DiW
64Lpv4doG+LLzMsWeo7cO8P+YICbdCc0pLUGJpRR48fxoZ4Tx46dYCmiLzWVl6sP
lGMtvWe42j3qpT729F2AIxI2EhXG4wDmr3y79MxyigqeLC0r56Yoyo8u38LddvL5
S5oEM2eabg8T42GuH2PgXl6D1hBRWqo2csRh8mskcQJU8F6qCd3yt9gvs/E/MptF
tzkJ9vQC24X17J6ezUiZ1St+1YmtoUZn0ALHc7p9/H84bcLgtN4eCVTK2IA6fxhI
h4CyhTDnnTji7JBzK/Yrgu66p1bM6xYK759MXAXuBegkRvln5ZWlTsDRAxX09Hv2
j0xbcpHFpYEmkMlZg56OoPbJnA+4OZe+DyUlp08Y1cglqbqWvBM/VOJyxprPWEMz
ouV5o0Htibs+E1JvwuyrvSBHOHh3XbxwtLUjrvRP1X7qAoQZxKfZf4wpZkjEjytW
dszgPbRbBWqw9guANSWL4Bk9LpNCl8QDEMel3ZkXozj6F5RmANw6aRqpphejT4h5
ANQZlKIkXXs02BliOmRDuKB9wCvmO3navZDcW89R+2ofkpbyMkdtVwipQnS/HYoc
QKrTw/6nRcDe1D2NJr4+PtpVi5sXbqpDI9Rfb1Q4yVtl8gO3KBfDdgpQ1EENrFFd
ryxyFbD5pZDZMMfAXhkcAudDPgwAWVkBlwCQ/kYqIXmIay3O0ITtfIXOliOuIWkE
ErfbIqDgZ947tck+lderID7AJ37rGsGoj31OEUMK1V4ljxrmg4EPEP59oWQlTUk8
s9OjfFQiDF56cxnqmf3TCp7RWW8lDxfrC6MK7hKfm2FcIQalthjqnnkLhgBZHzLx
rRpVZEK8Wgrfy4c5l/Sxf31CyUUvcKsX6DlI83FZKjhX0mU2Ln758m6WBG2ZiIJB
5l1GLzv60SkQ5+Qly6BOrdWsblXS7+EmYgrzkMl6eIgOECiGtpzAsPuXmGZmbknC
tHvXtvItuhpOp/AZczo+TF944006i4VcExSDKZGLjEwbrQG2YtMYIjR523nXUiVs
xE5C46eOAAY5BnDXVW4b54z71cMh2p/aZtd/1SKGmr48da5BhxSdKV1v9L+j2Zqb
wScRNkxdeNBoQEM/BzABz+EN9Xnbdj9/bciEyewOiNoIPVitUC+KFgJs16Uf0Az9
FINzv6pWTmmIBf4GAcual5Ag+lBZV1c/E8URVDc+kNMuzjOsN0gcW3ipRrjgZ7D6
GiZnHwTpavQjlU7/Jo98qMA2Z4IAoHvyEgJm2a0JKRc6pfVvdlY85vMQkQpyUQKb
jO/+FldXmsrTeO4RmQCiGMAiz1GU1dPgxIzefiTpeU/joM6SG9Vx7TS6pbWU+A1d
KfQNnl99NLfloI0+RYejvTyzXIg/KKceUxUYfCDZppX5saC/YX6cdm7ensG8dtub
qhZnt47CPfvS1IhX63rGj9PAP4mC6uTcDsRzvKk6otLJ7b3VtA26QQoh1pv3JT6W
IvoazkleqGaj7cBMR/sMP+WHHBDETHV1kXGjUvzs0w6PuB4noQGbCTd+zJ3QBL0R
zQTf5j92uvOeyr44hTMZS7G3c3G0jRX5D01TOXtG+t9SmJF0i4nBAjVCJlkByu1D
5KMDAi53/7ql3ukh+kTTdWqf+FgSH9lrW3sEe2w7yzxvWnyvu728rxNTPqVuyfe0
f0jSMQ8ODdvzdl9XjfuFAoG1wAbDZCEitsDymDvQHN8vbpPX8Wkwjc+A7ur4e8QC
c4B9H3yeZV+EwYutUWM04h6vkEf81PHXrQO4GxRJlMzY+BT7rIeHQDIAQ0GX+6xW
T+kzVOGJenkSQxxcOdx9jGMTCEwaFjwLYhSArNgW1DhL9sVZIOQf+3hBSbc7yZMu
DFOmZYixDkOR6JiKwFQypxSA0OwN2BRRK3/2KhzbGUGNV9VmpBAaRtlGM0tHzlCR
vDy7ByFG6lNuC7tw0IRm2l5JW7GGE574ZkflXT+ZjulR08TIKlhBqR6rlJKDpHB5
Le0Q7PQWWX3ZqZtq1X1GEsD5KDEeJgRHdUVltLTCkU7KLpZRIudb29Q6woUlqpYi
PqBHGTvi2c/RIZrC+0npfzlqWbn0JPhJhTNLRh8e6ie2OhUFpO24U9t/ub4UKdCu
Kw+qzrfB/mDSNz3nA2LA/HwB8r6aLv6+2Xr9gBJJXcqsoJts7kXFMUNrbbf4Da5Q
PgmJwit25vxHoEyTdz1VErFP4MdOqfkK9KRM+1oTUOxy7PDWlhESk9jjtHI9Cpf1
qs2i/Yfk9dDSeuGct7a3mNZaNw+cvgQUUrcePkjq8pRArjYUtNQM7sne8CvOBI1E
uf3PVUWoOLH5hxH5SWGiLVZCSt79+n6mADUc5GKPP0gr5J0A9WtaK6HD+UuuVupb
OAVPa9DRpIUf88kPR22w8bHT49DtzikeyQz+6l0tPckxVJVz7bKJSGLWNpX9V1GS
lRqyRn5qIPS7aJqdymeCcbiyjtDsxUTtpqpf0ipTQ51VKBPTwKFQzDuwiM7xfDmL
EF621X0ZcTsN734/PWr72m3Ci73g0tkj5ZFG5g6oWB0eUsiVLDpdoKjsv0acjG0i
pVxv41GuX67/EKlPF4mjpWaRULP1RZnBs62DZMiLByesjwpX6K+kzsJh9dwNS12y
QHuao9rkqJdXxLdDCzZJ+9AAqtC6AJyYHPiVLJWpANZrsOsbxrqL4XH4uZ5oo2aE
MxtYHDTAcevI/AGbJsfjWFIqxkhvPRQAUNvS3uO86tB6pwQhAI0w0lGqh5vO8OFx
XrgfonniHayXDU53OJmbO3M7BhDUkDpYiHrH3Xk+2E/352UbJX2f/O0NXxXSYm75
T8801/DSW5HbQNAVBe4Li2Y+wH+CNiSvQY9z6lZce7DSuTNpiLObJDx1GjLorVhN
mTExIOtq1AHVD2rjRUCH+rWO10abJtZfmptWo7vVioiqJ8GDbL+x5akYpDuTpuSL
zVGR8s+uxLSaWDfIegb7/iKGDlvzb+I+ijd6KT2WU1aNobSdq0NlNl9vG6Oiwbk7
skzeDiAhYD0ANLW1KtjS7CCmhmkednmnIZ8mbeypQt2C+B9wLPm28zJSBIOe9Qar
H5IkIajGQyePkA07JZjnkgEMu8iOTUbahmXtlgCzp7kgGCbjDg5uuiLsvnoZNECq
PS1iv7Bzvffk788Z+EyhNOeBNBXUsDKJnA+v0TRi6nHcz64xYHmkfjfndF6XDL/B
GzFGW5SvrJBzJkx9E3xRQzHLldqmsm+NPzZtrNUHIRj0PO9/lDEu+HL9Kf7GCD+a
oQM1xuXUl5WtNa0FlDY0fDJCJf5MHJ+qb+3q77eHLov7jN2Af8Yrb2VPVqMXwhEz
j0UCrcuQbX0qMmPEon1N34iv3Y68+slTpBBkyUzHv18qt3JpdOGXTJiMnywzjjFV
ymOo7LW19d3/xV6JFM0mvGAW3K4fcpI/ux3mmvEIsWTbU0DabM9TlKXSjC1iyea1
yuiuSELN044fuaH5qYCQgjmxZtXjZ7JFw1FOi81iiSQzpCHlvQamlfD6WKrFXAay
5jGqbb/Q75p3PwVU1VW8jjo09mpeUwLHPkq+/Q80+bmYsU/1BD4XA7yVz3SnlmK1
NFwmm986aQvEoxwc2CNvBJj95Om2YphUFfRkXOf4k+YQ6SICSn8ZnutpmVWBg/k0
UhpKpsouZqSSp00wrKMn5kW1uEB9ghHQPlKVkMevQkABj3MHoxM/QO6D3kwSFXu9
Tdej7sWZSBC7AdeMThGk9I3GqwMGj3ZSkUPB2+3DtuxEoJewd2c5CSeezOyFGWlh
m/M3iOyJKwo8RicH9+Nq3V5gtXDrvRSe6N8BzVHRgZTcGUZ6uro02g3TZ70o0fUk
9S+hVUO0rRY3BGXerqHUxNCa9VfUPPQJqRDH+GA6dz+WghPQ/vkc1/l6anBgUhDq
Omef+Lw2GSUQJJ/Ym6+2THDlLhtCzyTxCI2JvwNRtWwGZgDcvuhj8AGETt+Isn10
H0QNzEbO/OVt8VOTePaxEHYzbTjG5W6mmMEEXdiR48HLmNlW7FqAU7SRC87czEfV
zB/KTLTLll4FFdr88hMdSah4xv5N9zzTQRjZVIuT6o+qLdNiLoWSksPBb0ShVIv8
bA6bnNBRGSZZjsitZLIveSBkgrYHO1jt29Dyrwxf5YAxpAB5kgiyRRIAt7HDGQ1H
YaFcEQfYCe3bscdhIqVcNkT3BbMQuSUkMx6qgfIIsPJe5iz/fPgXmEbsWd2y95gw
k9eh+HYNJZXh+nT8tHs16Cp3bbNujRrCHEuedzv2CBUA3Y09uGKrlXXKtSUZFWZ8
ZAtcEu/9cdgvsrgfsAPBLRuLXvXup4ubr6Diyg38kdkRz7t4aHoFYZrf3p/c44Yw
PdZJ+mJqHH0OeOAO7BbIByWqnHIa3esf0wZt9lOyqZC3jk42yF7z6tf2gihplhaD
Y4pE7m6YUznSPWToI9nhe2QaW5vcG0DocH9CbWduPbMRqp87vGbuGiiid/lv8CoM
9ikyA3VdMImKGqKUhz2SEF/Q68SHS2udqgGxBEuCBa5y1L5BHXReQuKV/F+aPE6o
1JLMe6jhrGHeWwAAclr6yFadMv2kZkWJdpMCOCfdpC3RjlpQAOnJyS8OyFmKjDrz
G6SHQJ1eLHT7YqCrGLJ0DXpc3AGJYCRahnC6ZWTVSULF619XefnoKjrrv85p+ZcR
YTNTFnIRumMbHFElt+BP03njv5XRTHV9FfBHHsm14hkjLKymeORmfqa9v6vD2+Sj
b5AV9hieW+4+jqhcxnNvUtMmubO5nyaaPzKoRUbaPD27Xiq/vQRvB2upcOPYTXNR
+uVgdfMP01pLoOSaq+NVjIarvkkT1ZH9ckzE1KgptLIopBl9/f8kZG+kg69j+f3E
uGCv+h3UrGjMdSNwUjADrOK2yzCWwRdrblg0Fj/tjQcKO1FVlVkA6ujhsxE5R0IG
+DAOh5v/6sNY+pCUVhT2Dm0tqFaSohmFMv5erCiJe2l/V2Uqt9ty2xf0/P4+GLmy
Rx/VjL3TGVPu2MYTUn72w5Pu0ZlcVLmu1IfwUKccJ/EG4kt/JAv6/vKHx9kXGUyc
mlKPjrUuhD+EKmdxHmjgGE/dj2cTfl9veBnIi+4QpF0ie9ivjXTca9B9vPQpIUeG
FfvXyPnyRFEIJLgzcu1P0h2yVRAOw2LXUs/3o2V6SAJCZk/cBhIqK48Grb4ase7T
uWX1NHCaiPInmrfi8WVQgj9vPc08znqn6AA4MqnlwmhhFCEmmGo+uQPU8pJdjMem
EjhckM23SoGzhu+FyTqNJ0YhEKHuBlhWixV3Pwx8KCyfx0KnWvP8LI/DNno6oACS
3/QbmcVFU+V/n3OFZoDMSqSlgSPC7VMk7IlLXT7yaaZTsLblH41a194TZLRu1RYK
DW5NrDW4yIpdzuLh41S1AWQjhLFjMQwfMzGDBAbuapmgwmthXA61jNgD0HITSr9I
qqCJfyG1C08k+/X8jvhcbGydK+rPgtO57VErJSjTcgi36ww2E1TUebJGR4KsHrUz
d+9uj/9LretklHZhyLvo2WXXk/SxINBkKxivsVNb8IxBAdI44sKINEs2PAmL8XBy
UG2EH+rvU6RzsVQNYGoJ3C6lfES29z3k8+y0BFnM9m7CvFK9ayUrFQOES03osIWe
g3bZsjDW53QiGpadHljalU7A6zT5PaTv8LT9u2mitLR6fW4N1JmHJuY5oioFwdtW
KmwTdq7HZeTlnBbpquaG5jDS64p+0GJWf7kzUB4Vfq/vqwS50dPREloq1Kk+5L1f
gdkZFYn6csg86IIVdoSGHLGodfKPlAt0mf2iHil6Z2Wb9PF/jPc8nS6d/q8slKkA
HswV9BtslGv2tpuD6+5OK6Z0bIH/OOZ4Dl5g8NfkYcW0XqoZpde4rjH+Rj4ciF7w
BJySFNw7ZBTj8vAwGWA7Oc9xlJnCOXkrTMKXYLH2d87DCzRlkCzOKUF3usWl9qA0
oxPUZ3MJLDkly1xYscmwhQrfZVVVex9sr6TIrnEZr2KiFgE5zjxEvR6MBayO6qO3
HD4YS3JrCcltGUdetyUCwbWft/6SPrGqTYQsBk6Q3f46vMw6yISpJ+sISjKMFq6z
SxdJONF1BBdGpTV1N2R0kDgzBsNzc20DAovMvhdZ2jnXxT+K0HHSUu3Lp71Y/VFk
h7ZjO4ISlF9IFYPdeWW1botb6lOnysHC4PVXa2P5pKFU91d5b2WPb3bqWWE5bedA
L7LULQKUmy2dRZOZdnj4NB4RxAwAsTAXv4KYfrdJxJOUjDg00JzgtMPmKVIFyCvr
q5y2YUW/0Jr30MXVwRQwfraFktbv5VMdhPONiCWjGjbWXeo9vKBTe/MBTQdXeej8
InwVBqgTZ7hLlFAaWB52HgVaXRZqFha/ImAvNemLjq0NpF2gR5eVDv33a2NYgRwT
KD8UuSrBoLsEMlxiFAvwAhcLy0oxmGG/enXE2LKLLffL/yKu4NnQR9SIt/dGiisH
8FaFrESuK6302jJReGGGP2ekua5b40+mXre9O9MLUSPJ3VEcHZqwocNQ1oxeLbFp
C658P2nvife3jZjPAGLXq0xQIHfzvwaGshuv+Mr5TOZcok7uV4DEHG+esumT2jrm
CbgIyusNSahjyJiEVDUNqMI1ox8AjW05nMzcLRvcVuWH3raLDnQrm6INhvp6ZdAM
huibjG044NJK78dCmxZeGuD6ChHMwyXIXy+Hd+CfDJzJ5Cls9jZrjJC1Av8evRLh
MN3kXt44iwHnx33IxZT7w8ngKtK+s3h59gdH4LrC0EbPz+ahLLzEapUJgdFWNvXu
kGV7K/eIXzS8a0PHAqLvOzLuEB8ITUU2hkjst/56+seN3JdqlArcQr+1QrZJMylM
afb8HZ4M07tmUMZMFkjifRdHvuiqkD+2yd53WXfzMu3YQmmD3ugGINTJxmXprdlb
rduK5v7WWkGfldWo2UNIrd1ifINAvAo4v9/2ybR8UfjtiNnIJiQtwTtyYhpE8LHN
mSHeci4XtsatN/6qdhYzSb0IT/PQAxFP3b9jA98Jzyspy/aM8MGcJKUDlZRJ4JrA
1j8s4OG91FAwD/hot9oOU+kXnxB7SRRDzT0W1qzKTtgCTzgLQ/oAE1WOQO/IJtqO
+OI8RHDVG1+cn6g2bFPz21uzB+I5qPy1tHTm7boSr32k5KVBe/ZQk3NG+owKnSA7
/utf4bEU+dAyGJ3FigIjvAWroxB0kjjzeK+crS7B7VqrC/lZ95wvdt3G08z3xSvK
+SZQ7senh7vbuxV4/IHXqtuzsh1w3qB/ABPBvs6jEGVZwa7rTeESaIxe7dWZUoMn
kmD97YYi/7DYUk3dq10xFMhLCL4pu2vw4pM22rAdTJT5ZiKdzPhAAagSLzq9O1Lt
5klqjRYXiIn3H3hm5LtgRkBHvyFQjy7rZBwLe0z2BlAT2efWQJ0tDJQ8FUosCHLh
10v8B+Js2nrhjOQlA8U2cchk70QgMpkVp/s7Wo225GlvYOn196qfV9tHxpd8+d25
XYu3cY6iUig6Om1QcgU7iigoMGcmjEzq1t5EEKRhdZQlHGyDf6EvDr3jX3RBS/Mh
qtp3Zd0c+uFpaqH+5f8zWNl0f6szS1QjHV8dqvpNoRUw8ijmZyvenCYpg03ONgNb
dHMKekjEx+T45TsQB6kcwd31xu8CLZkwjxrNL6Ithbx3lstjDk9q1kgnEW3BDAJx
X9AeSm3y7Q1sGEZwSwkaXjokA6d90UAT3h0oJbwqB3DCJcFgiHMDFgxoKS/duT7E
gOaekZhP2OP7zMBAXMu2KjcMGA0JAtlPnH6q2EhWgExvB8A9r/6fYJ0G4sThOnEh
F9fILNIl9BTkmcoVul+oaGk9tUZLZnYDVGfJq3ND3bgBmVdsqF0faB4+o+O7tPe4
er6zXRaVyXNUB9i/M7jYJBEOLY/Gxfu6kAI5vr/L1LR4rr9ywAuMgYcUjZP1jfoS
zfODgzepH/QxHjmB+PgN5sdYV+wyXRMq2/5lAV96zB8p7Ywq2vxpMZvKEHvQk01i
aQ4e2ba0cAN6hS8/GYkbuDfRpW+jDsnC8uSCQ0fuN4bEC5ufY4eZW2OK5yxaJcpn
35CLH5deHTVXftzGyAyshFKQY6M9Tn/s0RMexzV5snydKSPY2o5JtPPtJuv0LHJ5
xOkJmI4OGXj/t7uyVHTm7dhXE5oiy36WPHneSl/hOWp6KlBWVlMcd00Htihi1EM3
McT3ajpdC8mxFHG+AjaQq70HpJxzRGG2He+JxGTMJk31WXYanhwyrFNqP89SZGLd
kQiHxu+jVXLWBU2fLO9TQYo6KaiGn0V3rVsciPtDemZ4HEWutZAUGfgB1BOoKd/Q
lZxUdXCIfm8BEhHfdcPScnfYcXtTX4c5Vm+plo598wA/TDwCmFMCNNBiK2FsZxU1
jqrsYBaX41D7PUkW+jIYepKQNxeOfXTNvOF1rHe3kT6GoI5ce/6NVmJaBZUjk3F9
C2i0ze00a8RiiMOe8iMqyyK6q+MEodZ1GId057mPNm/f32qRPtTj1Uw5ktdbljLj
qJ4Ka/pSRM2BF7XR98K+JJAA7UjbLEJsLEvpTf5GLMzNwGIloB4X1cvgFAcS4MNV
kk8ILdiAd/nJvuU2LFewqx7iI3p0kdqwJst0bfJkqGCcZ8FUmp33JkfZ3PmFtWuC
/8knnXTf9Hfydc8PFsA8VJDfTSKMXCduyhf1KYi6i/h+SjBCpTAJEjS1PVuL7hV2
ViYvK02ubo7hXcPoTdMG+uXyM+mrOGbzRaUWWFJNt2axNMTAozAL5QInuwG24zjG
v7PjIOseMcOXGdd+lom2I0Qha76xtI0Sj0aCvKhM9XByWvrjf/beA+h4ey2eGtVW
O78zDbWkBdcVkExNrol89oqVZkOyjznagtzLb7CygySLk2o9P095iU176D/MIuPM
/oGrzoeXrQw/JI/0RwG+I0DfFRcJB7tc0lH0xWS/Gz+704lr3waprgGl0NjooBMp
ARohoKpmSNyp2htVnqt03xSmrOKtuo+udQK2Yo8cORKbNTJlL8renc/M/cwjKMdQ
NDxhv8pQIeqdZ85gwXts4tRTtd+AR6ZTmGF8QA/uDvzhJsA4eArZ5hDAxsIjxZsf
6chuLclLTZ9gzfSPMHGVS58UeoBwkP+ez8W+LT233EamoNqtuZv+2bcCbV1uxxIY
ZUQd7AeU3rQjnozOLmz3kdq+0+QB/JHkyDxOr/rF/d5aUdktiXoQbGlweH8BtO/p
kSLldoKI762ZmP+VwjnzfrAybDJRlv8Y5hOXtVdIr2Ipl5JNEbC78uWFj1o994qX
o9tdK8I0xy0ku0z2rVVYDUy7ztnZWqkEgifXTF4XY71KNUsMdmIW98/jSM3fn2fk
w1fOzYvwdIOkIl0KCKLcHSBF74BDdgsc3Gifhh9or0s5lA+WnizQitPvPzVdy4ai
9xZMVx/3aPMfkOnmxFd8ttXhboYASZWeAaTIFdNHSKLcWeKiYJFa3eoSx462Uo8n
cFtb96HHQsOAS6P3QaSN4BT1rhwsHsXDaEFM1nA8Sgd11OY2XkC95gkzd/nD6rYR
D9fVOMVfV4893JMGjdM4Phn0d2RnrUJhV7gvvkIJihY+wIxuLAjP/nguwN9QBV2M
WUDX4ZsiQQOmd1zLzZZTEotOvA7yCc1IZBdDW0CpNNNcLNT5336vEyCF71oCBEgr
IGgZMLzBxLt5ZDWLJplbNIPcpELcqS2zKm8rTCrB5vdnWVgtluSGrUgSVGyGNOE0
W6ObWvc0G37WIm0jKomKxkDCnUnMg5TtT8mmhVfmAW2ra+dJEibmsqAsM0J5fhVU
r2Mlg3xAXul/PyCxBBNo5Cc4U6wVpq1sQwuDbtZE3NGAxsCNhR1R4kTJl9oKP798
Z25I4S6GvoIPCwq4llKZ2Jk6Fl7Zz0Tltn08snLvajypsoayyHUYYYvjSXqOaBYA
ttCsd6k7yq5ssNuOLhFKyE7bGfSqighUYMhK+CwWhR2pW2RwDcgth3ItctjhvFuS
SmrMEGh/l6ohdtUJsn318b8S5l9C4n1MsB91cJvatJ8u5iyb0/LoLTFSx0X1XKK6
L+ZeKVDYO7FugQfsXBpikPbGFsWbGO1qkWwx9A0tvbNPsZ1F+z1pfizDkj1UYyNi
/9TOKurDshJ/We+QRy+dXky8/bWXVSfKGdX8CLI45yJEatgpPP3/YOfnPBC52sev
GHZfIPzYQZusobAJIqBVIrDX1+rtixymoq67sIhVWti/RpU7d8FPH69myyFkIBky
4/1h9MJYMRB8Kn04vaCHlxROiDKvZ0moOjmKpqDao3NJmMF+RCo0UP9eVR2JrY1q
glKvrQKPKNdCrTWf/6gZKQoZz2JAi+WlQoqy5dxiXn1Ti1Mv+8FgFppc8JHK3/HK
jNWy0AN+BpH5Y/33uYWZit6sSdJrAL5xKdOPvJmQu82JhIUxY3v5adz4vebg7irJ
9ZSwi5OK5N+P4X6ExVVKxNLuiCunlq6d0QoZH6+b25kAMS8ulJnTbEqPt0vwv4k3
bDsMT1TbWcoV+bk0VGl5ojD6UM5CfU+wSfSLK5ZUhmmpvJ6fT5YO6M9aGhYCZqp8
Pxb5uFSGOfIxarBAaq3c78EAmY5eIaUBPmXTtn0pzs3PQreeLKbDafRIrL2u9qyy
98QyUmBmFYfBKYrYwOAZ06xa4OxJhb3Lj9y0eTJWvHXSnNH0u1T7VC495FKW7bFE
rHV6nXDFN6TqUXADLMX2wv4saKERxKpkBfk1ufG2hdeeI+TrVG3VmF8yxn0GdfBn
bSKftAbbNPfB7A5GLdgfnfqwm+ek7JAxxX9vp+uG9449UXQimI7eKvMITakwPt74
8FXO5zMPA5HoyelE6Yowm9LMFMfdKpzEvVMPkBhOk7MUAPpcuec3ewicTAs/GKox
4EBdhKitFRdPlYM0R29n++VSmkmNxn0No1ds+EWsLtmOUJEvqIuT52VxYMeeZqTT
RtYD25bxhD4pKVfFL7QWLfLsC0ifHMmCNlZHlTWpBE0EX6Q0SjNtSWeoFZFZmrEQ
reuf3RNs3OoCkIWNvho0M2ViZPib/cCMRkkej6L3L4hJZIibujOI5oYpfJ+4b/5V
QVI4v+yAOVeVK//OWtFnIVdyJqM8mcPmX1RCzpalnnFolPEG2iLiT3KslV1lv0d5
AXSGfTuZz/Zwl3DrbB23l4VQMRYk+DLpJk6ZnlQlQUXaIgKFVd7MOJgNHSC8rCRN
ijFBp2K1yK+OzKLvSUB+yUsBDn5Mx9emYPY3hsHCVoDZkd1d6ELSaH21UtMRUeG1
SmCZnmwQ4xtuq88tCvkqJsltCYzy/Xcdb1Z1GrGzQEowET/fTPjU0nufuhAaiX27
NiSVZhxoNdIxgZEBttbmsFHVehuJyFKaNJWmCfPhYYVv2evSSdWpVcQn8rrF93X8
dkGV/ZabOPsddmTKZ6arIZ1rliGMY3fcJfrClLRzWpCNMaaTgnrREf1VZfiEdN+s
26KFcYZTYghIqWk8G9GU3NPSCr6arzk7JDhegXWWw7StwEt5iGdr7Xqq5lfy39vf
3ubYWjjucfCQeAtLU7YU/rJ8n9uHuJDUQb9YSd6CAGJci1e5YTps89H0IolzlrqI
h4nIN7+4t8vjeuoVbXmq1EeM7cvOMJt1k2lppU5I9VN34imbChB2Kmx6fgu4D4p+
EmL82aFMfpnfsymg01L6sDiOsqXrG5oILKRsPz5pg65JWSl7572Q9QSNJDxwfYdc
ONyTk7h6hSyUHG10hBHx7AdKS9zer9gZs1SLyzRsuxi4+F9moDjYUww5+ZwY+ADX
2SApX7XTAZ4QWLiyYGOUUgxH4D74+FcbCQQLNKNCg1lMLOCuMa6EkqHGmkXYrsuI
gt0PPU7enqGBoebCQn1NkqsCDHR5OQd0tadA3y/0eIUAxxZHNKbz+DXBHba8XVAJ
EoBBkh2aiJf2I0sSz2P6A6mTLSOI3h8Ap4BQiAcUv7jmxuy86mjT2HeSNe7xwCyy
/rPeTjKZBS4uTZEadaqaLhmITSXM7lXbEQlSFdMwF/YwgtPasCFTrgsKHjspbUVC
IyLJWVutKg9mWYgIUdmKI86HklFJW39BV6+UFaFd+rK5Yw7+DLbCngdbkHUkLcN9
uzFMwNf8Y1fTkDi2ikxWoi9zJYW0uU8aCRgsrAUPPwdaeE9brq+qX8boy2n16jyb
eflhHB/piQuRDdp6+dAWx697erGDqd/1rDZEbJ848p8+PzBiPRYuCVrduFEw/NQP
zN2FpPQUK+0HESmICSXLBXqveB5MqLc3Q7QT+Lk1DSw6/Fly52xA9lXw/fx6z1Of
oGbAn/hdrWZVbosZgeZynQlfoLfpqn9VMZ3XJgwjrg+XDauvq1I83FXWy+Qj2UD+
c62sY4YGCNkqciWHX5UrlsdB8Y6OEvIxz1UuYJjflo4B2dQmtk62E06K0mzaTVZ+
Q+3s0fduqE28R+vloa8RUCZZ1uRv2P7vnXwM7+Lh1ucKrhXJw8DTzniG9oObGjKr
K5IUeL8wC2JDsUmg/tojzRaOPefWicRYAadv9aQlQylCU8jSTTpgyIxgvy1+4/80
FsQr1q9YXj/2Ijy3vTjY50ptNpDdaIISMGe84aF8Xm0t8ilFEdtJtsehmDCeuRgy
XJhaVBsZE2BudiJXTgsEBFjII4YZ7/BeCHr/WvM0FAfiTt9AwYfM0zZLCAipcjxt
xbbN6gyTsV6DyvTBq6FQgp9jiN7/SeyzdC0/GVLEEDu5xhWT5CWDSPe/U2SE0z2j
+v/aZ9GwBTVKGlUxe3lJsNU6+wFH0vuoMmT3va0kUeWbSkCrDi18UIzeMIesSuZq
dEa4cboMVFqKkHm3WMnRAQk5Rs4MuATsVmRlDUQ5KZnzUVOXc6zkERBKdzNOGJQ+
zvVXdBaZ9L+Owt7cMFcbXaP54+JMIMGlIjFjzLY16CHKxqVx0UaT64edBWZqrpyf
n7hrSG57WtoFJWhQAUfu4DTZgZWFxD7VrCcwalApaFyXOrwV/5mGcCkQ4A2PArH2
ENYh5B0x0PL8oPKb7tn2gTUiP6vuliq3r4A5ootwmhGGiOEbLCRGM/y33Yjq8mn2
lOS8J64k4iEK3mrHj3/OzkvkO8WtkeM5PWHucYUoIj5p9WItecE0hvhKi2BUdELq
GHHM5opcP/EILauVahfVcX8L8D1cTMmFRQivZZ8QQ1s9BEoEnFnWa0OWTWcfsPIa
yr/7OzQAyToRFSRUB+9SazVClO6IfcpsR4KUMoKPbNy58FOH8zVYko7LK9R6hWPy
m8TEgzvCaq8CXHKPiHSACLfvfpmiVH1WjscVNdWGah108mW/NlrzpVktSXn3u9OJ
kw3VbQ4J54EXbxo67CTE89shB+iTtYeY3x1/H8h2S9/ZyLPArCFIB1n4RsEBPKgH
O4ifCUpbQdPhaF6c4E0ajjbF9EsY6qJWVExMVRfW+Xy0DJ5/XRodD2sR9gV1OEDa
RyhlTYrSb7+qkVr/ym1ROW1dIO66HMr30WCY4BWU8S4XqiEscAVp8/ll4q44hz7k
MndPOyWCzgpLiJOCeQCdpw+RbEiWLjiB/VEb674TCF2LBxvBIUjwlkobyZI6q4Ua
qg/j7KEhoBlbAGjOTkPqdHOhDRe9hsjVchg5ytzqg9qWl0H0OLVPAuPcnkAEjig3
MRvlhUXWTbWfHAgR/kKVslllAPVx2xI34xuV8P3lsqWY8+DekXqziQ9m29qkJKQy
YdO4WcLYdQaHPj6rwINZtAdx4oLNWS8av1gEDtQIHLV2eriot4sDeW0GvXMez4vo
VpM2nZMyDFGkH8UHGFTNn/NvCPRA1pyuOyShqQzVWIEhOb3rM7eE8pSNOwSyA13y
lHUmIPBMZk9wIF6FjOZL38Mnfnu6ai2Xf2pX7Fp8/4MVayQlMOG1rHkEkeqCv4/9
8YXGFT6DnSLZIq1aOLrOMilDAZFGWlnMZhDmaYW37a1xIG0FXHK+2h9BEtGxFUJv
6rnkbW2bQCLmaB6eNn35alw9PVQNzpDTo1wl4SxRZViW0A3gn/nKpPZoGq5UHElY
g/2CV+OGgeal6pnm9La0OmiihTAsp4h8LY8OKw+rapGV0hke7cacHz0FVPiqit4b
1DOxREhtLnXm3LHStqod4gQMBr6hMUdR21yzW0mcaDVydw/biCIrSWe2ypr2w5nf
/SYz4l031LKGDV3EDlk4u1ZEc2W1kGDSGl8HhwW1/A/6kof2R9KTIH+2O5vy1F+f
vgsfU2JcFlwY2oIY/tjJlXy+oc10BAUNr5/OQoGVYgN+kspBNyg0a9reE4Z0atDQ
aOarskflKGOFyYzu3wLKwySJDqiD4y7xNEZS0qkI5eyNKEBvFuo3nhRdSxgU/+bd
TXmoykLttXjblCn9Fdy1pdod60Pg5ooB2KQm3ZpluHfwO0vJNj/n9WRJfmCnUowG
TqWZXwnTbLEMWzHJelUtql3p6QQJon8Qkbcy7okfMfAnxfYpkYG8geiUY8FSbOKo
b1k40ztcCxRgLhl5SdaGzIHdVACFOqMQMtQhMF1u/SiV6XRc9ePukOjalNFgE2aE
l6v8B1UmSOiFVO/g5Ehk/fuMDp2wDajBb1g6Ijt01O8pKD4RqF2RhycWcJ1HzdDY
Q2mzGKyZ9SS2locJmnHHrSpNEICyhg12Oe35EiVcle5oGRV8UtiGbd3Jbk9PsVvQ
1PRdgNcpUmIIookLt6ytqGw6EmVD5c/s0pYmzBTbmg49hZKEB/NNsgtdeGK90RVr
N+y1Kcdnanl5yGHC6MPz7wK3QQQu85wE94A4wjcfZ39nXd31nAtjnrBN+JmCifZG
K7DMgwAZaBH5ZEw8jeGIB+FfPLn6UnI4t0Uv8M/QUFmLwCbFT05lGSPuSsPkq1DJ
YYoJHz+UOJcWIIcnnvwW03uI32NraRB6Vx04Fu4P6RzPUy6C1NBIWqxFm54NI9AR
5iV8SJ9oxLqMFcjdDWQm/1Z4pCO/hTB+A5E949nvX4laeq3flSGTsrUfY8SgPdN6
ooM2xpj1/mnxxa8XzbiBzeT7Shb/h4oGq6ZbrMvCrjJxlSy1Hnpg1p+mMAYjDarV
2EhcifplgUaKzmGC2B/+tEX0r3kSuoa3LPo2J/lX2Mp9i5BFH0IAXkROnir4gDj1
6GcvWVW+Ww8Z53dCq2IKwmaYAUpGIy65KcENRmBRa3uwePqB3b7/sewuP0kBxo7D
uxvhgVxyh50oa1Kxukv+As9zVPGHgoY/z5TcI/sEixvY51BLZc15Zh/WwEJpyb6z
MxBw3hYOg8QqUbsYJCDLmjauEw62WqzKGdlHyOzWXl0KjVHLEh9FePk56WVGe12V
mNuFz2Ymo9japXNhEn0pbrR+yTrtdCGJG3jr0SmPIjAB9ZHIXhnMIhhjlnU23FRL
GGlHrBcITnQsczVubdQHxUjWmeedzbATG4FCsMau0d78oyg1i6PwZsCIUIuIEmj8
OWDHPSAEJkAn+gnjNG7d6eZbILZ5YiZpzoFgTxyuN7/Ny7nEMIhuiSTIB24io8sT
3sr0Akq7yvfs+cIuSO8np5gbu678dLlj4uWMy5e3iVyQ3a3k4LpAihzeU9KsWfIi
deEg0eVxnlb+K0XUcMhwlg8m3mcCkaRvhdt94De3UeCCs1P0glkkHv6kXXP2odom
yufUZuYoE5xZEJsNazorSSxhX0MYavU2D9rQ5JUEJBPPv3HsRI2tQhAu1U7fkguw
9MpUDQ/eH5geoS2oUVJfIjh1vg/vBeOah5f0b1zKvkfrftzz9qIdAx/k9lRBU3pS
G1eqvhvThoViR2LaRkn2QQ05z5hfg8jZTQhKYzglUmnhznIfanOyiIi3Pr1LlikW
ucQOv+5dEVKuuuBWHzIjhDr47hDrA/tEZr+xjbTSAAr6eCWhC8KnLrQbDbrN4akG
GD0E9anfMq4GhHcQnPXx6SRtflVLNMwGgtnWLUL6coiKohMoKTLTPqp1Sm/eu9Df
zi3AELmlp6rY5qhAdMxb8XJOtL7djFXB5IBukvHKuEjcX+VgtG6OkwKQfa99JXcP
2jxo+I4IujPy9YHW6XkKUzfmS8gacYJn9YcKHdBoYO0z4x2Vhkigrcj49FFfFJIG
CjZejbfeBRXKhV3opgfGicFLGjajENZvL39aV7UYWZzHMndtIRxeqpSRuYXue6v8
MiBpWleSyjQKqNfq7gziJ9iaurBq7qpM+l+pybZeoZuMMwB0Nzkcmn+rFdKbOsbv
IlGk11CaFF3SCB5wG4xq8kuJEJvIIUgxsNhBMdFamkKUw7bmQKBhi2XoMbqk9a6j
ZGVReOZ3xPXNVckKU7m+IMVgeoK0Hod90cr4D7CaCsi2GcxqLMrIauEJyBXajbPs
2+PtKTp9XiN8R2ZSaltCCuSKNI3IY0Z3DiZwsr8RwYPP8t0zMcTWrRo7o4T6nwjV
RvmQgcbIvpEcUHFSgG/6bZ6dKV2GKcIMBYXh0U/ccV++qwtea2choRhPYT+5luVl
qaXXJxsnXKDLg6xjSpc6Rnagq6BPgMK0hQrXsCCg3D3IR+DV05ATa9qMLKvZ0J6T
/h7o/3ElsH0Ub6Bgt0VyYEPb+6EMBhSngl1lTFNMIMI/JAX+UgE9q6tYOT5TGscJ
X9X6ELr8TdXyRmM7VFYMi2MvOhK9RB/Uf1+wZtMoKcjohtv/aHEJBfCmsXRuikoz
ZP36ace1qYvqz5N0FFI1EQwI4KN+q0bq2Iuk7/ywmYlzMW9tjXuQ0bT4aLbNUvPb
DyHmIgiaTeoxeqMPwfjbYBYV1mq1eUtVPrBzI8JjehOiGVGOwWhdf/qRtpfoir4L
sp0eWNca23vTorjmqvcACrjSNaEqrHPdDzP6dtvsqlyNjaw8DVJxLqoBFHjUTj7C
YM5N3ZNVb3bfAnEyfLyA20CSFmleGziiA7JciVp6cstzH8eYrSWxB1apBzCRhDtt
HvM+mlohtZs6vo5XdVJZ/E3jKKB6Ibv0ruM/RkA69g5Zys2/+yjP45HNQ4Wc1QLS
nruFrC0hbXya0veSmVqxQNLzXxuQwd87WazWhD/oJwds3M4Wudgv5ns3I1tj1LT1
0pz3XuFfD8lB7MhjxMUCplMduCBnrPVNIqSy50FWS/QmL9quJekGwVDpC5BcNkJu
FIvtYLFuGs9YtvyuQ/ZTrDKbs1aRXbOPb2qzMSb9WYI4aV3hhqdlm+8ACO6VvKjB
ftoTzX/BFzKdm1Hwcf37cx9PsSPRmj/tTlUysoVJR+x4Ns23RiLhG1ybQ404++24
eVyD5aHtYE8/VTts1xCzGPtTrjd2QEPtBHoQXdbS4pc8b1r649fyfoC5rFKx/18+
zBvjNEnmr2qQM6KqGb7FOnI4NQkGX9ceDNVfM1Aiaz1GQj4/YBW1JVNsQtkN1hmc
OdXIzRmVkN8R9d/ZEwPW5B/jE8JMC/UfS9GDuI7UHao+RHRy8sTPBJrCrJM0VKc9
VTrvL/tldp/4EwNDEXh1f8ksv1kfijVg6KpGjCpcENzNPSaUBLvwLdCZ1lVbF4Wt
lE87EMv8vz0nnHVJ6zDwan/iradHUs6gph06hZcpHQGs3E8jZr8779PW9DX0cfhz
Zh7Tdky3N5M7u63wUYhXlHp9g3rFGTW/MAlzT27D8jkRTCvns58e5vkYP5nOBcEn
pyQN5u6RPrTLKEG2+5bnz06iZM5OuJqjbltdTwPYPnRbyXkBb2lLGBkfQi7BGJa4
d2+wbDIKXzX6a7GyIFgIttFT7C2kj9lG4klOl4rEIy5V1eECTgIQ+oLMzHofUYPn
aIoxj1gcUjXmvCyKzkV5wJ4YZwwCjKOc7E+IQc1NCxHhoiCsRHzpN8Av+e93GDy7
7CUXpinL8qw/9gGB/3HsKhas96dU+MI6bJCSGtuGfazP+qE64vz3e2qHnYnYabP4
vh33NUWm12Heu73V6vLV1Jzac+xbq/J/3Y1VffY6pcnA7jI/EAOUChmirHS94mTc
nHzSo6K0kigxOGcXWP7MoJbQwJotSoUIHGHKCLf98SmOLjbsN2EcFV+hi1jVV4UA
+zPRQ99472VB0RhFKpYn5nqnPY3sINcpVoC4zu8tfe+XCCum15tWIVeLHZD37AR0
+cR7wK49N9JhBt129Jbvo8oAqHrvXJoq6J8dfL70LWc2tBWY6fdGjFFL+CTwGsWM
U2iqCu8jKZMQ/SA6HLESx+/LLhO2t99PgqPzDtu6ileQOIpcR3a0vtSKl0Rs1ptO
+VPtIUq5VkMjgFE7PCZhVTBl4VKyOYLGV3tLMG5icCXwSiKMsR4PaNox6Fqu4vqm
OPMtBL6L6KuoWlUQdVfJgh3mT2tHmn64yTgX6xuw8w5EWKT8ymEma/ifADRM1nJL
LVIHi+Y2JeLIWBlUKqzSWyxiEi3ocEPYYchzKqQw39Ja8sJJsigK4Bv/0HbgDqB/
SSIrH/rV4R8aY7/5H+vnJTT6l5lLPLQumAwqwjv/0ikh/qqvJWbKJ4i4vxqFWreB
75j+yiN3yBfwtXqoXy9lkeQ7HiC2zwHktIFIX4AvzrBWgUXSIizeEUTNpmbEGMMF
DpdTjkYLWcFSYzZORlgcV1ifRTU4iQ1Ak3oXwHGsk0SKZykQVaf84dEHBAVtXEzv
PAKHsfTyz21TNr+5rC/AnxjPanWBwSD/ITBiOksb0qKFKG5DeQ+vp54dX2xLhfxF
R3W36/geAcTs626Atg554ftNBY40xiEOHDgLmnvyg/F5N+QSHlTM8VLqDpX8HySq
9fbPJfsVFX/t7gFMr/PMMc19mq/AALPbXotyaXoTt2h7UI4xLqSV5yahMfKHjGKh
28clvKgRUhqHr0NbL+nXMflg80mAhMSjF3l4sSD7NLB5AeODRr1kR/9U14GFRUHe
Ab9fiRVEebxLvKX9JwVoYtl2as09JVzN4Sw+QBv/ETeP8buSZSlZpsNA27SwupHk
NUD5ip+p3tX43hkTmK2nEQhoYkk1cHBK1naf8d9YxlIWBM9EZgnPf6LDcd/NQ1b9
eXQqXrZ7ocJR1wROoDoeAhVIX2zpZ+XHbkeYNzl43TPcOv6FuQTb6PoSCQufrQI1
sA2ujhQWawZ3v9uA6Rr9bmzkxTQmZx/0wV9oyiosCHEOQzhka7NhFCrUDZNbULmV
9VXtHdqKtPt0umQaapytajC0lnvgE8Qlr1QkXrc/n/7aOyZ21KfahAGT3ESRnleW
kGKmKHxHRUlEzX6VqiOYB/yQkPYYGgsS8OHyLwKcUfY67t6P8KDDy9Adn1EX5cwJ
wtsRr5bzco1CDAjtHXHvwJueE4TehTMIsgBvIPE7YnqwfuvTOTiOx4AiWXIPfutV
WD2w+IG85JkWj4bLQSU+7l2Uxi4CylfHkm22IjYvj22J/9pYvVQYk903Uf/ndKj6
55afggjiaJOHo823BBGtLL+X6pJVIJjU08t6i1Of9q6p/mXnEpGybuwnGdd6xJAS
dNiETvDgctUTU6CaysE5TpLx3wcz3EcK7/FAYV+u3UwX7oQ9klW9/2x8GHAZivWj
2GgX7PCKUnIfjvVMn3u43AgegF3WqdgPJgrsFgILmbq+JObY0AYVmWXND6mNSDOF
UcXuPOhPc6W5DfYzKOjOwPx8WMMK8fRXUxXhFln2zedG7SHxKfQtnGApn62KoqLE
tG7QaGEWgbik/qa7I3w/3rTbG0hld1ayWh+JDG8G/weY88UblwXNYM83tHTN8V/H
vclwvutFm1JNv0iBidT/hfD/JycUvKIu2lPh1Kxr3heKB2nGOeTu0XUS/TToaatd
`protect end_protected