`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 12736 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/9huKRhRMtvnNqb3Z+UU7TahEoHV+T8U3P3ufru7l1O
3DlgtZzb9QxCbOjthp9+wDkjygH0eUfDrEl1ovhZG61BwgeO0brwmGAAbfo/yptI
MW10lwV3lwHGTABCg42hCNpfFJ9mxDDRAT2n3MnwO1v1+c1sBM2DOvn4QLRgx5qM
wJPrtq8SYQ2X42WlVtAz9Cl+RHvsazEQ81irykIcmzlyvl4ou5PD6k1GGKiHk76T
YXkaGuJxeIffIYHCHgCcq2evK1vD0Vp53PezZJn69bXYzfoM0d0AD4rAJGI9c/rY
VlOuCTRQDelzTFWsbfRsmlicEPpnzp2OPHwQYlSZpE+ruAfMsemteh2A+xH0vl/H
Zy32CC/8YZUBt9uKkrJcnr59D8itsVV+dG4x6rx1fncnXz3l75EsIJpYUkQOjSv7
K5yMXIkyekuB1su5/k9swlktpbpWlrsRaJTlit0SuDl9QxGqUGqbi+ywz4F83Orm
gnym36fCYregAYtxhc0E14JW1n1qxkyD/edq8AdTKo3P0Jr3PN4YR544b2sYAShI
3nf2r8vS3rT+btKwFGsE/eAxooYz6p9nJUk93F+ZHCuRhLz11oZ1ycq72Z4pyRvI
0AXXTUsWYIhnYrgzGYK9LUbO/9uup50JzYqtdEDtS3+Ni0wlhlpIkhPAVVB/mIKX
UHEe4hm6TU0/NNoCl9Ff8uaI14ufyjTYYaqxM/6GLh5PpUiYGHfcbOVGD4yM4Qlx
hll1n7xkDYeXFmmd1H6p3GuK24mv/gPqEPHFQALo1fBjN49GOZVBWVkPhB22rHFB
0Ma46fcKdzFNgFx+0alVePXCSQAdaziNnGMV1JPKpTGbrnkJHNiKoHQ8xqrBd2hq
w2lQmX2dP+GDK7q/XB5JTQTrIb6E5qTVq9MVRwY7sbkrZd3wI4zH3S/fMBM5QBBx
gIfzfMlcR0YNZhrx53HqL3KTa0qQBQv4CzMDH3QzqshPgp8bXrhXG8bmywHe9o5j
IbJk/H6nvPowpc9gn38VJECF13rcsoakw5dGpR5DG5HN3dhkxxcjr7HUkTUo/2wY
R+PpyuMHTHoFR6+OSf+bg6DIbx6kYzv0mS02AA5NSfTjeWqdS9aD3LhZJDsIjUQT
tEkzf6oPz+U0LPK0H30bs0ro07kDLY8Va5FYp1Y8Jp6dEY1ZjKJhZ6lkMlBLw+p4
hbeGkXG3GV2WV0csUneNAyEAGOnVkdi6e8rr6XnHSO6fXeYAHp6FqadwYtSTdEok
wTcVb28GSyUeVSmuIIFqdXAEvp6OCJqMzXtwV909HeZoyWuSBZt4dIeldVmDeGJA
4T7viGipTbSLSSiy/aR4whjPhoC3zxiNAa0B/jgXoDaRutgF76Q2X8FDmhW38yYl
PiOIbbyOb0FFcXY+sAUGEbIXO2lt3/fO6E0XQ/n2FvflCGEHcsYqWiPR4GPYFR6d
13JVi/Kn4h+JmyS5GX4PjC4dcjgK2pClBU1vDEP4sT84bcOycd+rENjHndXLVBU9
cGnk/VfYsjox1H4TbTBEUC1Bv48JjuyziN7M8otD7WMDP+7SWOO2vlqTaPSFtPgG
oromUIy/3SXn41g/yjcvcG/TtMUj1T8zm4ixpL2+uhzsEuH1zMk5CZt3A3PuC11J
XoScgNxCKt8ESZS2yexFxbfMME2Z2y9/pizRXZQMYEtdHAaGFplsdLdKQIo1ScVg
py1vGThz5EQ2TzPBJeDzKe6CUGaZ2ZbQsM3BCSXDaOFg8Izr/zwCIkuagWLsPWAI
bp7q1NMJO5+lNbuffQ2BRRS8AdZ0sq+jNH/1ToG+yVLNsXccxSBESST+3jtaJiR4
1pS0oBjTrAdXt+8ZAVQQtRf0G9xqoGsLaGLntEHoaOpcCaKjBoNSUT3ip1FPnfF6
KYLucdNl+VoYFP8rgqsiWnaSwJum77DUv5tX7KDavihFcE98mI7hc6/RPFsi52bP
s6Xv0SZ0q07dKsl0x0LW34lgQKF9GdaUw0WOLRn43A5cLob+dAwKO1S4ugD4QpN1
A1L6pKk4zTvF5inIVQkNa8C6rp3EoVqwM9ONCh7UszWasXvZrU0q4ZhCvxpJhcrt
2De+ptZZE2AT7BwOwLo9IF2tjMk3RrpXWT1kTy98GMpe5akndwm2zAZmHDdJ0cKk
7Q+mtUd9ZcuJgKoL1YU27aL/19kHm/f6VGdPhcpOqhvL+JXb9OtnQiDYpEbeTKV8
jsTUN5gyJXrvVCykeQM7tKPkmIxS6K07A3rzvEK4eaCAkDV+LwMlVxR0abVSR+1H
e86KurKU0D130NzBTiRmzWLKTfTbTNKZs6KHCBkgZBiT3Whm1i7rIOhluBT7YYIi
56+mJbJpdQhF1qyg231e6vccaFnjXB9caEcE7MDCjo11MIIffE7u+g4h0l0R9Vh8
0xIqIpjnihubXxliXKB4vPVx0OwKiY/xoHP34ylsBm/WazrzpXjHtnzX3PZ1ABFJ
T+RztCXDjMcU0nE5ImmZPGOo5TuHaDRX0Zw9Yt4L0TucG4Oxj4ovJ1JSN6fZxalp
3fSsVOvWif5leZtM/KWB1BICGcyPBZkAgigbzyalRpNX57giYInd73lYXjZNCwXL
jyyzbcWTO7LFOxGREIi9DIR3vc4a6U6co+X/AAWAb95JuoOGjqGPGW6NACrZo82w
/Yu8ZyDsTRFr/FcIQ/uflYyJq12CcN2JF1YACCNxCULIlZvbIIfDcbWRxkcNlsn3
vUwhagtvd7Ks+f1ISF9S6AGPgy9hozSQZ8+a5CbRcKl60GzrZJoVktyC/sxlL6BW
INnNw6NauL+U9+CsZHxJBNDcGRHUxi5zTsWPoYeoTNsWRmlXDlUrIpthG5tGeSZD
SSmOkpmIh5oFLPZzo1sUUZ6XMzOurmuivbns+DcEeQosBWry9yhg+5k2DgIrA6kY
XvcTGZKqBGatuuYipKeNJMxAWtOC4+vnevx5uuiTbSxN6SHkCIoJI1r3QEM0mhEt
NWZIBLqovRzStF+pUCNVnhGpyd3S3pxgVLJ+l6EY4bMpMsBJH9CnZXSb4bD0QFKx
u1s1m7eDrUOSlEqdSC48p05zZbctGBHkPRYSxSR7pYLBYu1Jugv8JLlDpW7n/+99
6YcyLSjgPXPbo4N7nXFEl+/psy+Y9XxwF/ocW+ZzyQ4u98JpD4JAuUhaUpM36Reu
RUwZDCEETEpKvgpQI2tRPAgrOVmhSD11WeuNvIlV49+4sByJuyY879yFKgP/fS9E
y9wx57oR5DwTgy38vTiOyE2lhKwQaMy6A7WyioqzOaK4ebZWe4SUn85QKwy8Qrr+
F6gt6G8pLLOQnLg/QDHy0laNnZ4c1cMkxeT7nVXRrR3ZL215p9LmfFpn59aPdWDm
kPydNFQ7K41/NOiTzOV4EAK0cDJoIMb+R0kAchHv1SA/MWVuudqYW3451phxBEIX
H5vWsWjobeH3vQ13B05DZrwE4EI/9gB1bVtFY3Em0pMTyzPaA9f8IxiqBMkwGJWx
Z3XVSApE3Ai7NeUqatCTyn3jRqzdfeYTLtjbqaF7S2nCMojvkxMTuMJh5iCXLAnL
gYpxjtB0B8tWzAZgBWeMrC2kXJYeelshVUe2Dwnw5G1hUNaH2zTZyVdyMo2XZLAT
eN027b5nSqxUVhhDmpK93Rw+KyuYUQncURMCQbvYlkQTuVlJfFTcodznBoVLXTcn
0ymJJUwflkMF7+NCMbzFJUtOvvX6yOloyRPKsH3oE8AAs29BrT/N2ZPd4/Z/J9Ep
MSryBzLTo9oKnsNW1p2u5Ap2YVKkvHwPQgtq64dWdipoadq0/LDRbzpWNdSiWZk/
4gfAFdY3veM340367ttnQmk6+SDn07SWN3AM95l4vzamXVF4qmeFTlCB7Voc5Yws
9R5PfaTmH1pWmwrw2We2CVSGCXjhZljn8l69ObIhvkXufzFzuKp0GiGjOlmE3LoD
o6JGwo2VWl13klWV6ZUymPFpg80j6VRMSlNQ6PyfNvZbUGBb/U7Yt3Afcjypz7VC
lE0tVfERi11J/B48qHSXKQm4yu3F9hoN49EGmRGkgu5jsQr56ZTM6sztyBpjHiy3
aYDFeGwZwfhpyt9MnFaHJ4JQjz99XxlBR+erpFsvH0VZLlpOdFWinK1zjBStb0Ca
VjXLsbadahC7rX/OFazJRiqMVUVRvt1fNHyvWGnwnO/x+LU9l0sdG+ghCW9jn8Q5
EhcyJFalH+tIX649+ScfA8fWpSBVLjpCUKVIGq7SZGZSlQK/Q8zyxC13AGm0+pOL
Y6D+ri2wJWLTxvL5qz93jWkejdtE8tlpnQw4ubgR4AeatM4wUdDFpbConyHrJMUG
Gfk+fkSRB0HCwGNZzEW09L8I/GPEpsfRWixRAVp0sFcsOvkKXHHILTJgR+9N6GoW
xfNsfjmihROv9hea3fdhz1DdC3xty8liEo4lii5Rl2hbuzIJv5Fthar7gCGVvEWQ
0JL53yPWD74cBSEDZBmP5t88mcQvvWtPE7M/vK2ur7iu75+QL51PwF6hV9iv+BIY
oAWtSv9eDA0Cm1XbTd7HLzFsiZy85E28wxecGdW1fwGK6Yjb7HeD7pi1ESfAtbiL
vq1GSTCTsQhtP9yMgADPVNhdCR4mTSQPYtAFUzts7KRQBLGHf2JCjKKXCVM9fMq0
C1taemO72VohlEAFhQw08PGta4YRA3YVRkyjeq3kkgXXjjUSYk+1aZCInZ3rYVuj
VIGMcQQAAv2+wB5S2ak9lead8++h18fyq4dTqAyS1T1OWb8mZrIzJZnWYJn5Gyxd
68L+gIyUu6CFMM7aAUJ78s9QduOuS3Se0Bj/QkksZ+vqBDSIDBgfuuXv0Me9+oju
0xs89w1mtD0tOqcBcrhomzmPcY9zBtgiVaqf8UAAmCYzfB9M+RqE98dajn8tEWqA
6t0OHvneTaIliDiWWC1Js1Hsz7iEaZrwQpAjmFgvkKadqvMjkjVDqxJxY74Q1KoV
KV2ixrTZ961gzu0fpTaYY4jmMEN073fiJU7Alpx4qyJYmfiMioCq6RDu7gYS5hH/
3SS0YGPB3ZATiRIZndpL5s06hIZ3nU8CaDOSNpMY7NesK88tk1PunTeQ55wjM1p1
8JofENqhYVnnoBBWJ17eCI1ShQe6fpIw1Gyxwd3UUGd3Equf+7XUR9J6lqhKw4Y5
aVbu4E5niZHVu84VZME1oU0ucGEgC/LBmk8LHmu4DZUr1fkl6dykWzOENZuPPrpt
fuI5zwTCEG+81pkGoo9+zcCsmw3i60UBhytvKysnnVFP6jiu24JcNztQMi/EjAYe
Hy57SGj6JcYlL6IC6CgBWXDd8rhaw8rFpdsvyIUHzoX6TCoUiopqazsYENGEWLRH
Bwls6li80JUR9kM8LPerg/MjpXbpzKBYxkSinBkmAMCLREtaAvk3NWFPvqTMBTjH
R8bBupAigefYqYXpzhD1CbqHDrZNEEejFNCvf8nV8pPBTfAYR5eC3SzRc4VaQQg2
r1AHVaFVgSxULtRUFv+asYQ/Bxoo0/jo5aSUfmz/YskIMecVxDMlcuzqSnGMpRXQ
kCrpQZgPRavKn5YayKMsHUcZrBPsDO8l7soMW8wdG2ewvBh9IrpNHfRQqNFIaeeb
cvkpv9JyOhX69FA2IqhR4jYSs/DppGQ/0F1wKR8Zoz2yNmP50s1bSGWb5/e2DoHa
Oj0WxxWq128sevzqi3EoUCrPPoEzyH5gEzVTJK5kNBUagScFrLwlJtS+R2g+B460
3efBtCUnZq7Xam+jPF+yhw6LNMrluP2RnBN1qcOHajqrJ6bcT+9bBWCMCgQs4xnk
tEhxN5s72Za0UVvUf9vGYG5LwXZTq5GdTRnqMXbEFiawpd3caqMp5iNhSIZKFG9g
o8siNtyEKWDIvZqH4NJqXH79tsDkwyajXH2uwloJz1V6lELuh9FDRrQIud3gtx7c
g9axU+rPHlhpjszBAjOeqq0wvZYlByS7e0fDXG5BwNtKZLK5QTmUoM3mZT1WIRr5
C2mRGiZnfadB2MUy4BlXLB1SGmNUJpz3PjBWMRVnaPEBZyhJddY6M/QvGpfhx6HS
671JphV87KytGiXnW14EUt43PH6Dwf7rxw6YLyfmYlM0C42cO28hIFo8MQV6eFUy
G1HMkZxtS42r1LFpJxAk5todFD7WHzlZq2UbC86q+bSawFPonVDMStYCoS2ARdlk
MY64BopNNi03ZDR41xJYasTb3enFTl1nIEbcD6qt8WsP1o4TPzfyl6RH/xoQJE0o
r7aCM8TX9Z8MpfC8uE2weMtngh8q39ZuTNc6hGoz7sp1Udk8EEgn9d/LGUZM81gV
dTSrRhAB0Qvo4rL9RCSj2GgC2rcPhv1SJXWGjCv7NkVBnQlUWpvSYYVOqq9OFldC
//uyqmIGK033xspTJdaeFg/Rn+nUAoAOMXpcSjGGfB6SlNQfRX+wVY08b3M6ZUOf
fJcZ/TJSvZqIeJC3ts8HLyRzSQ/84EUWL51ifsD+j5bVW4Vh6ySpSNl5VZCN++Wm
ssR7MDncniv2NNnsDd2+Hyee2Ncrj0hlMQ2Nn4ENfqWRR63KnHIuhZEzdB3C8Z1K
x+STgG+JuuAcPv3WMsL3LowoDVD57UO+vsoHZK1DmgTjmpsFOcbb03rkOVLZQoeU
lRhzX8/FL9TnXaYkngQwOCB54834OVmx3edcMM4b3oH5MaoLg8bCu8bfjSdBp1Lx
h/80gzDXySiLPxWDptEmbDpeqUfBE/8WRIH7WBxxS9i0oXw/I/O6IGb88rJROi1i
k1k7jH9HSMiFrIcQRBHqFhsY+p/jJrwA+QSnaP9SSREfoapSKIotn5rhIt9iCAp8
hkDpuYq+y0eDQyRi1OywBDcfakRdIdrdxJXhokUmXI05vC0CSOVIMvmD/sGmICNM
sMfhBM1c2a47z2q1tY90K/n6TmW/qxcdkLFdwkFLiXb7tLLpIVsCuKIqD2YpfH4L
Kotm1fSL0D9ZaiH+weRSjSGrh6az94gETBBBS5vmHjM1/JDVjTLI9NGp41xECubE
MQCo5rKdwiIjiYcE/WZ9JdmUnE0jKko4A149SQFqbAxj8MqNMMtPh8Zt0gxL3Te0
nHVLdNrnKa+xSEs4iVdIVEJVJuab617l563jqOeZY1E1J8YSRV7c9XBLy20BpZb4
ywCY1jvu9qbdU4wQ6nwkic+Daw+xNiYC6MrmxBV7fMZdUysO8NGygbErGGmbO/nZ
BrkoClN3I4l0mOsLUkTVxP8f8plHxh9TSkHVvFtO8Q0o+bCxRuRViVaN1LxQpjdj
8KzKHLmNk/hMMV9Ye5WX1GMqLa+CPZDkJHLVXy1wqaHWlHbsFAc65dwZOznbyakx
wJe8fbO/3qyXVMOlJYgIDnZlqj3T9VBp1f+EmmzIyYF9uQDNgS0Wk2qYMV+vYnHm
eiNxbr2QkTigdAoO5d0k8qG+j/SNToALSm31oqpw/chFNtrZIq9JXififg4ntwz3
88fCNFaLxnvPTCggduCwhBBpjEIM0unUvR1WePYM3HzCEZ650HA2xNPQjNc40mYP
05Vqna7BtiRPI74wTtjwk/Brb/pJGXWIEQoSF3569HPtUNlBXLqQbzt0o5XRH9MA
tTK4xDh+5ZwDTMGTHWVJVvJOgaqw2TtaPqD6dBfnf6nhTdOCHe8hI75pwgOH8uod
1jRyjYv1O9uF34Xofifp0LpkYZzQk6xUylK+hEDM1RCi0AjMnobQuWHwUn2ZsXgI
imKAcDgBQBNEhmfBCcLjrrRl8YHr8UaMeHzfbPj98z0DJvyN30D7MT7jIhDOIL13
Nf4ndIvcAgxIfWSqD8h8l60yeJReL97yS6+fnkEoDm3zrrGmjsNZ2cWvWiHpem5P
SWT4lOQpeJWeSyqwuAd+jL37OfEXaWb6sGVro7uRHVAUl0na0q6UtKpJnu2cpjqg
I/LngMEdYb1d52xX5KU/bFxeHLAPRT48H3eeXRbc7a+g47TIT20RaT1xI74UiwQa
CzPsaj4lPTD6BxZa4SDO/ccUROaWJXFwT2HU90jA2dAdVIDmYRMaYb5PDWAlD5FJ
mSEvH5QnU3b2K176GGlDlaS7uejIZ1rI2r3qTyMAZlBemoLsLmPyux1G2TYAn30M
fU2Nl2+6HHw9+eaQC9bjuvTRGEN7eabEV81Tx82MhRTfPRZRrfIHU9gEUNi/D7jd
KjzuQf1HVbZF8JsFhbZuFzg8TAAhUHbmcYQIjKv2PPfE1rbJ1aM7oBRwV5xp0zus
L7x6UW1VeaZxfglQSAQtOecZCyUFw+WUXGzjqpv9OBW6N+anAQ7iGWneX7gN4ylZ
ca0/XfID//lKm+Ak4PMsm9k2crlj4K8/3wfOq2gF+yuk9/6FniTK3V0xioPttu02
0F/A1mguHJ0t4E2KUiejPJDKRBb75qkI3UX0vFZh3sEocGy66K9jwlTEMS1+jRZG
5mLbdx3OC2KyKgwm7/Nm5W1aKNOCFlyxparnBEBCsPTmEpd+95Qp6gqc60MyBF9K
wO+gSX8M97+KQRFdA8bzwWB68jGUW5v+ulyjprYJhof2SGDvHjVDVeN17jgNDwrH
Amtibui8vmmuxTsaiknEz0fO72nFTxNL4k8wVCqX/ZgV20EVYIYuzewsQuAADpGR
mC/gqiypHwqTIbN5/lzgm0mcn5HQZQkI1ZTaka+bwYEdl199tqic39kEYRlmg7ov
+DGh74l0xJHpCe+z5M5jvkZIhuHcA3KRPOlsa11dNCTOAaWV1eDQKJTmruSV8EWu
JTfst6pgewOGnA6ZFgbjubj1VjTA9rsHD+JrHud5yUa3VxXyGFFvC7c6jaEsIK4V
mhkoUPrOSrO+3H/+dI1ewW8VoXqrZeGxaOb7nV3p2tfK8OGgh2zg1AX4BZ4BeTrE
1slI6Y4WaQ3GBQJLKCNtNoQqBc5ZaO8cI85sjAHkrWIeCgmvejTvCRcas5VT03Kj
hYE9CnOSM9rRCo+TCHCue+mKhbaTkvz1LCapOgfXatoCIQ0mY6xrDGwztRnINcRX
vPyK/121PF1Kd2j8Qn16cfU0p7DwjfM5d06xGzT+9LEcZ3Q8eGnCbCc/j0Va/OMU
PZt4Qiv19r13QgxfJyIDctrT6cvF68Wb7a/LAbcuHZ8u4KtSm4rJun0Q8rBIpihw
pP89FsSN0JFOHPM7/ncItW7Uk+sDO/Pavv9lcxbXgPvs41DLgkfJ9DIdd4gJ8ByN
sU6mxJSfoADpr1zOyIbXYsIsewu2i5kU94Nq8eOMEWoA5ZUdNlA9gull1F//h3Ds
15fhK+TwwXVsLkdhjRkyX0CkJvodSYsE0bglzSzjusULZH2cGXTBr7TJbbjeUC8z
JjEvUUK90BFdEd4Vn2EZBexEDd45yySTieZQqSmUJzaPaMfvhTmrbAQRzmWmTRPs
Qq8xtqxZ8DiwIZYmN6rBfvLDws8sOAR1UZReRDGArxnxj+LZofVCehfBIZhheRLO
QYiKWqQQ6dWb6bMgdZhVxwSlbEupDtRLklCM1rBvYuYjyETgXTo9eED5O+SgbxJl
v+eGCC4+yvaN1koVa4ED3rqKiVGWJi7xhRoWNkL2WVWRXCGV1C+lt+m5xtOaTEoT
w9+3bgvTjzFgVrB1uY4WDqpd1BxiyuTOjSq1R/33P5Z7NfzvLet5rUU4HJYq1yxz
eWzTc/ackngNBTM785RHbdPusBwkS0VNaVMMK3Ys2r0Pb3jHKdZ+5zTCCGJ78tcM
ZHIGETFtw4ZII/MMH0ZtwQkRswuUsVVw/CZ7r/nXqf6fq6EizKSDkUGK3yUQ569A
Mpqmy+jjUlap1Ox6yuLx6I+p1LDshfkr3CIL53u2kLNzHM3vRZNVbRj3YWMsLZXH
ThkJ4+51Ppi8K78F3b849ET1hGrZhwQCnbaZitj9DOFSEn9i165wyy1You1cqMym
ZZ4lQCwoBG+3PdeK0jT7vKsexJVMYJD06t7u6ZYszCUIHmhzV7fK59WGT8YXj4Q9
N8LAl4OSrVS/dSCyELfI60ThYSC6o9pdL37N7BKPIqByKf22Fmhf0Sb8Jmvnm5x7
J4zSvnaFdmkZl/YEYPGCx/xL6oWgvqt8g0pIz/nQ9fKr8yzlgFEl0MX2Uc76qDeq
04/qX6G9smzQHm3ro0WOXz9GSW9ywCSg0wVjiWaADxKdv2nA27+VoNX2WQL8ZIFd
XAL36NLOSC4GkEJt1KHmy6kN2mb/pHm6RHz1TL6DeVOFB1a3fBi4VC5JCAEbNK6Q
4DA7oaLw1uJRk06YUeNGannW6k/HKs7V0tEoV0h/9E7rFwdrMrTR5oBgWDJ3708M
0oY9YtFkXbKH4GRa7ylMT8pMzWg89QgzwTqrIY6lLTTGXsa3cIPr4Vbks0r/Cj4W
3c8ikUrugT+1+a5S35rpC1Wai0FVEL5RODjtru+unctkNuPP5/ywYG0NPU0exNVs
qZb7eCcSawkgfU1k89x4C8hCVB1q4Pg+k3F/K0lLSzdEY5N8rmjTYECeO4HvGXCh
0whn2naaA+RmTeYg+ppJkWpCecY55qbKMJ2UIFH6bNU2KhpvG+t9f56WrwiQvLTF
saIXEkQWlyprdptJHuvTWd5oNGDnLXDEOm3B14YM5J5nqAlizhCQI2KIWmBWkLLQ
JutarjOubh5Y+EfqSyW3Pzu7Oj8f/TMC+3bLxCvrxqqiRHpLkVxM2cLArhx9JpvI
BYwVBUgWqHDjkrL32gmYSaPM5mKA//JeL2mCyKWiJpfKBJUL/RP6HZkRHWJJynKF
gvvUpC+pZXdVqqBRU8GyIn2lah55tpmXXDhQ03U4y0q7L6XGEdM8idxlHIAb/0Hc
v2qbJgPYjEC9m3foSvEo164PrVGEAeqDQUhbk+U4Cl1iKtwyKJDtLnBGTPWUCaSQ
eQe8MS/OT+eoqDbfX5VQI1P1AbZFHefCeUGfIaGfIt2rs/LU8tpe53OT00QWSPOZ
bi1ArPwVxxrlrR8EagbHa/5aILYxUHZlyyqyG7N/kHvStDAXAwDZWCUJlNJr6iww
+vZhl5sDikx+L7cvpk0R+kdT7/fhOupqaTu2mckT9demWwicODim8cVwbD8njV3j
cgpExlB/VbPgCfbUecO0fXBDPAkk3WHa3o45KxZQQvQbnVClThQpfwrd9O6BZHlq
SfUjuKwzFyG95nq4XVrXBFTz3ubcLUYhDQdxX2hHUnHEBrcz4BrhwsHkTrtzV5E8
Pvr6NTYJTidFZqrj2Il3cjCh6caJxQZQ8oAFDHodxaH62rEA3Zhq4NboV1S6Ir/0
NJyRX1WV/vManoln1t1kjaH1NsDZMSawQLBUbMhrlxjSVB53d4aZl4tdYuLd8s8t
Orl7NPdj8XeiviYmKrcSGHx4rLiuUUWb9A+bN3yO7jw1C7Iy+NZYOGXao8sjwEg6
OqfZQR8rRcUCsfMCxkYl0tUz24FY1gB4gjHbSq6R2WlPOlf+8lZAeLWu6vJtQvuq
xO+nlB8Lw471zU+Aak7I6I38i1gG0dgVV564og5HBHvYdLzBSa9wPXmeSWZK7lTk
DRTiQMtwP5Ly0Fwy8VcgsLBCfkFITkyIiZq2lnfVOOpVkeG+S5YAJPjX/7LSM56n
KeAdYFSddIDR8bBSBIqIuBBdx1BXYqAKTgHmYXV/mECrvNk/+IxpJ06VhZR404Yc
3o26Hw1KhdLybVW4D2+d/5TF4r5QxBLG7GUGAp/pHY16zSKgKZcz+i9Yd2DkBq+I
JMT5IokgXqtQ2J6HBoEMDGsZRs8OPt1d3U4qFRqfhXC/t42dzTEj7aU6JaqSbcqy
tVTA7EJqGP7PugfnUXyN6Q1+/QOuuHR6SjhbSQy854AbbEyAnmtwkXJaZy1UBip1
8xql34NEQV1VkiHmYMpmFDf7EoW7+ep5coO0XG7Is8W6Ht+B7ZD1102O9eWzd07S
mtVboLYCeeHKOwZaz4meEITB0L7nc0H4JquO7cPaawtTJgTMt4K1uIOt8vt6WguP
ypKe49AR53EfwShHFLPU4UWdxeWN/DWHqCO88Km3+D+q6zpL7AAMjE8jZ+ftx4YR
cbpXTPexpMq7uwaICy2VjZYRJ461J0vkkpMKFhFUV/BgWJUXhTKwHDAboj66V66B
hlHYGzuLlSc3ciUazlZAJlLGOskBGK1pzNW+qbbzHrDaJbC07cquHsod93YLNUjf
FbGd4ws+Po//aGW7NsJg9sm3DPOrXwh48EB0GsrZVIsrCGNB7CYS62oI6w0g7Y60
yugcP1e+JEenHSzdSQzCn5vX4h+duRLHaiDFMUehMGfC6kePbcWk5iHcffKLPKQ3
5JV2hcfj2aa+JXo5E6DAT2EgcUlWdGt15dggmWXP6kGVgVA5Mey2rnl6hhJw12NK
E1ozSUZlWqjaTfok5amDEYDO4R+B7L9zSsH2IgGg0m/8dytyS7RczSbx4zg6s30l
lMQ5MsHPheZ79JvxMstQpHJGxtcmJ5agwvdDAlOjh2f8jL1b6FQx7b4yAMD0SqJI
BUTpjnGalx/dIcf/WTE50kR/cgd+ys0hZ1EQjPephPn67Ztbw7QCL+L9IjjnzmB3
hmRfovKBy961OM0LVtitVOemOoY+YT9OhZGDKG5AQXuOHvgISb19qC1DZ3O8DhcM
ilRe/G0i8OQrmHGRRcHAdqbDrNm32HGy8ugHvle2qsenes9GuSHtjod2ACLuvIqz
AOsHRTMEnuiSqHprA8Y/gs65htzHLHkdXFjRiZ9IOAxZluYBAr1psSmBwNOIKcvC
KAA9MFkBXXqxLnYw4MglT+H8lNzz19IkyKvM3oSmwVItwIQaINZOIg38AcY+S5/x
s73iJQySaSUEGFToEdSxNbga8H1/IcLqn0oY+he9lu4XT6u80aTfrdKsc9Xxb+kl
9i9upC3v7NvZCUAbuG5OMOv8NC/IWCMOeCZOoSjUu6tOrLwXIGMr5kPe8fXGI09k
Zmr17r1dFB38IAv5U0F99njHPYdPykfKHMLAVj8Gznb+/1P6SUDyh1kSb28ATViH
H96uIRMfRYCrS60yw77/fSk63Itv4wQrCfu4ZbyG3/KztlUy0R1iV9oM81iXsqJe
4f36qRwiabI+a5GqipcHT7zqZF2XbZ4zH9nEXKzzzcH6dAQMkWMKZ5faW5EhkHFy
Yho1LZ+HmT2Da8ChG5P6W3KcOzC4URhDyl/2qqrJ3HEAnfugg9n9qKqQDBXKzS50
teNz8aq1MT6Y5ak38a6sIBaQ3duwP0Ov6Jcr3CuSOnGcUXvW2SCCF6l8aCNyjCGC
sc2yPdxI4wJzcVQTdlw4ngis8655f76H864FuFTXE0MWqCj9OXe5W4jlkE7/OXFD
G6/Od8HUlL3ClQZVWZRYtNo3oPZ+xyXTXentzw5TIVoRoeYHzLVN52NQXaarOwGU
PHaZeAH6ptn8uxdqY0UbCuPvn9gKNtOG9Ue7WZ+zHvlJ4jDd1XbuUim1c71RXUev
xlJmRqDrjY3uSk78w+bEhJANWiOz8XhXFbG/feaJOkqvMuCB4TKr4OCxK4zr/tQ+
s21lQFmTE7g3dPpoJbFhaNQqZe0bGUCjCLz3MV0XbY1nheSuYRGy9KnGn+NzbuCp
kScNX+JoldiAEf19X6wfENdiiM+QF7TF/2ikKkiNuRILyq2CjEvPpPtIco9FDU5a
6Y8H2dXFayVPwe3Z7dpSeY5Le/doFewiyP4V6znFkAYm0uq/r5qqxgaMueuK+efT
tuBgDyXs9mZEmJJof9BD4BRnIQI1nel43y2DMk6LYgBTwCkly0njh9fCuZ+nqy7O
wVIZ3SVnMIHrclMpQyeNzoRYcJ+GN1ssR54if4iGyVXWy/qfGiwaRFp3T0az+9WU
ZTcjiMBmoZYt8Q60HWyoG1ZEcP000KUctZ7Gh796wA8C0lFbIQg2GAtAXp78d8sf
UX+qXyIKhRAwu44Llm4lO5wQAVK+5j38EtpUlmRh/GOSDoMK7E61CFQ1LNHPuYeW
8imRlA7fI4XVKrn+d0/X9rfau7kF/54uV2kiAxhfdT+hE2jIh3v2xZohJSPi5Dfs
8qYXSxfvn72inmW0Jbp62Z7dzrrfD5hbvLzzYuzY9sNqFoIcVfmz1YzuQusPnDmc
1rJfQh4kCUb6auW1XqwPSt+34QQPtTUwYHJZikZMZMLi7bx7uabpRgyny/+781AQ
EZr9PgNZgc3do43BRakrkpmyZOUYliidDcz74KDTmF1ByZza/xlsqqt4xO00rewu
D4Erh/wfS02GZbGBp44exuOPOJ43jMxFIV4fMe2FuXxOtalEWmVzyYf57Vhg0K9W
t0AL8qz/LDzv9BvqMWBQiKTz/1g+n/ZyPMyDmC49sKEWddfd4e9GeEshPX8p8L6G
PTJ7ZW6HCqjzafAtQS79AS9YQ1G4uI8NXpVCOY1q4wQa0ZOItJuVj5O4UwjZet8I
obX+x6B3ELD5apRmvu+lFQ6HQETF2rr040UpNYEKUgV+qKFQmTEoAqDVaeZZf5fS
H09S9LBxCGHRnXzORdUsoi3maK+WBLL/GeAINyQAVVVZOZLcaDfv96K0yk4PNAN3
lomp1RhBbOvCRG5hT0iJK3PeRXVbbK77Te/OpDQNZReSeUect/ZnVMrB/iRGbw/f
l8RCBdFySLvYhkWQRezkt/ZumCmWZOM/E/7ZD7PqsdcdYIwwdSBuXG/5aU6qhREi
bSvNwuFnbFU87W89lUSZa4useKz/UTTAYu16XBYYwgd0TvuNZA+C3OKczr77Piqa
VpCnU+F8smDQ16zE4X/N68Mx/vjzYiFq6/N5NvmglXGTD0jwWEMEBOMjgZk7m6DM
1hxS87it1iDg9uSuhltXERItUdWzsSozyjhqACmgbAXOMoq0Z3EKv9hJtYWxxzc1
wiI/3eVmj+UI7/QByhnshdPdGInvZajGLRXo3Cnqn7F0rv9cIfR2SOI4nF0FXXCF
cxAHdMpOnbKplc/BJtYZL5cPG0j4gDeJhIMQR2BCE1KcFSvJDBsfcOkn+oihgnGK
xy7Ol/T89v4dy1Mu7fYfTYlmaODtKxNi7iAct1QQn3AX3hjs9DYXZ3X54gKZZfez
uyKEw0XmcLqh1wfaenw6vjL6t5In1KD1i3DMRHUfLUJUAWCC5A1aFcFKo90cmF6m
sAS970/7Lb4prwPnUGBwY/RpwH+ABzqEALsVEpzejzwJLnHWrKBU4qT9ksv3A3XC
Y+bTBJfYW0oV9zm4FzeE/KsOuc7Z2AWt3zPCTm2bI/91OOmyxZy2duAZgWukzmtD
CKgJ9Dszu8vYmC0XacM0MHhafrCfKts2XTHchlUvMnsKWyUwHIhXFNiRI0UG2x+o
JGn8SftQqe70YV+b/fKTAJO8NYzMSa+HEUkeQsElvDvMSNZo9gzJ2qnq1+3qDjZO
Rqe27do7pddVNDP5PRmBnvPwEC/N5yDmiczV/7Ow/A9WGxJczw5JzrQ01p9gQVSG
MTppVeFEeAQzgTGlUL3ySWsMf+usw+L29o5hPFo+i7bxrNL6VSQ1uIGzp5cJEzlG
e7NKluu0+lehmE873idXyJs6mhSdgXGiex0icW7gZ7D+o+6ZorGTdxpBV+2mw9YE
ocsQ6FHasoMLEcJjifQ53mzJV6IrYMtRlrcCjoJBMk0bvwqxBm2qYkhY+MNWy5bl
e/LmdLl+FtjIpRp1Tq6V8+ajJNg2CwRDunxfaQhNpxzHuuYmfAuye24WVexNK/4Z
cd+IwcDp05G8KVEkhZH3hOY+GMAbJpfFGLD2h3vEC0UnPR6azmHU0eSriGYcKnCR
uH0cnqsDHtYQYyVRH32KlDJiITMvSoU9iDAbikz2R0vzRPzjSZjjsAfuUwJWczs3
Ggko6m6OJitkRPjyeo4jwGVE5GyGzyAbDU+PdLTEzqMd/ukKkXCEZ1SWwl/uFkrH
CSVGKNwUTzFvGGWFfAhbeZf1heQEM4Jak0taxf7zDg3Yyd4JLZ23yg/eTl0pEovg
QqVweCSYbla2qF4SAHKT9Mjuv+ix0tzT4femTvIhn2/kqCGHlBPXI/PcYEPm5Ts5
dXOHGnDBdmyjBECAB8DB0MZqRJfcKxGftoZJ7kUs0TtdJ8BMLeVGIYxDMP6+6gu0
Vf+E6+z49A/L09LUQv1ypZ0YjWMuuBovdJXVP3Y9qr5gHh7nd1phQnJ4mGEYzja0
URez6nRiGJVf+0o0g1LUW1ltuH61/SVV7M6YS04byTItK+34wgFX6SiKqL4fojY9
P1gdMLr5xIGNgEsiH6kp9YUJDQ3JPWokcIbRRCtjj+C5BZt0SW+KbedXC8Z/xGF5
WBlk2L/o3O9vra4e+qWE5gIqrUuD4CM+OogbWcv266yXBxIb9+1K63IgLRVFfCuI
7KrthY6yTQC+7BwLULQIJKCcx6CkFjXngsI/96GMCS/QySLln+jvpR7J+On50To1
ZyfPoW6+tFjOOI2O2l75wt4VdnOlG69WqSi0wq+xoZTAasBYnJV/Th9Xa2WDKeUC
q166XtstJ76fH5nTfXDLI2hSUhuKMgpr5afqNIoe93k9i5RcokLq7/rQKo+E/A8F
tXl4nvaZtcJPF84J65jCbTQ4MeWej7o29aNYFd1VoSvW/kKmbJRM9P6CqGNv0w6N
w1qiusQD7gVFTNSvAyQtmC6TLeZiD0XaO943F+0qvPvZsKIQsv1aRrC6uoo+57Rh
ctJxL1HYPm/HLjxyNG+CLi1dvxBxSEW2stezhyrgTUrlZHaxkiQNmDhThgmUWu3w
TSInjadg1MWG3puqRISoAjNwPCZKjW6e7Sou32WXc1901F2X20p0j8HfKgNtxBRj
F1QMLkjiiPv6DM3tmrG/50jPpaC4qCaNBbHHISNpVpxMYsYEEruVRG1wtKARjgv2
Y8SlqSsUdb1/DZuDszaFVOeFQNZZHAoz9fpolzhZI+giQ+U7WqVMFATMGU6+muSA
l0xAl8vkPAibHKiy6Zs8mPUFUw2Sy/QgSiruAYvROyGjf4EaHF/D8uk3G8BCw16T
o+kuhYY/do0t3pBaEJRwQQ==
`protect end_protected