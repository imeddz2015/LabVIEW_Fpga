`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 9392 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/9huKRhRMtvnNqb3Z+UU7TahEoHV+T8U3P3ufru7l1O
3DlgtZzb9QxCbOjthp9+wDkjygH0eUfDrEl1ovhZG632Qni8vZGO2IDZjJbx/uW6
z6QC0pUt4BbbO5Jdrxc4NQ8D6xSgyhjIOVglCS2/0Agi6MH2rKsMkhx0uRBXtdTE
zcMqGyvIyyPk0yDR1BTqR8rp5wb7PHrTqMk4++WjSDl+hVmH3qiw8fyHGJHKALI8
FbCPao7jgK1JmSlzZD3EG8LATL1EKHaH4PfmzCUU0NY6jVhpg5bDpGWDC/GnluDE
hvoqbhGahFfx9CDTFv6cFQqYCTjd4AeIrrrYo4ISReFnYO0fppduVqjVgFxI2lbF
FVcuQhXBxVHIYaL29o+IHJuBsv1iY1jOMs2qMoAJ983rK6tHGuERRsG+PKptNCvN
17vg4FSa0kxBhX5F7+aLcTo4qhkzEWOoPjdyg8eSkd4or4kUMk56UO/jXINgVNEr
KORBjr3vCE+/RQbnutOJdnbrpux8uwgtR3mCD4MJOyDap5fpEw46CVHztHPXKp7V
OVjhaiw1AtH/uJcg1O06MMzgKby/yKup7SEbles5QU6gO5/0cO5iA1Cgve9Z6Cav
kPMG9Kc4rFRRlkK7R0opGTQyEvBmO2P8hkY3qOSrTiYVej2obYiGqMLzwN3brVG4
UbFVzEPxVRwXzIhYbMrfLa8XXrqpxjKFFfaxDCeyZDx6yRO3gZRGAefY9p71N1Ae
yxjxL8iYEQzXbSoHYpmlJgyf7g3gGibRNl07iKu0kzWWrD8NML9QKLxgEpVabCdP
8269YJAs9q2elgxiZ1ISMEZhKbVzmkI8ZUB83HARR/u3SNSOprKZw1Jnf0ZFOqxH
NY+lBLYqLv6qaUi46hsLOlT7qdqxni5p92ZxhAZN67hD1QcjYXhedEn6lhEra9Ay
OHj3siBEHHGb8/p0HwG3f4DvCR9mXrybaPgwebBfl3HDgcy3H+CDlLkdxqCsI2hM
YFnVKEzccSlh9bVBuXXeUjOxLSN/G+2SZw2kHDDyRY30Fs7rwXJ37PlDYMtlq2dg
0Jrk1ANSw9OY4SnxxH8NyJiHzqRNGBdLX+is+fazxzS+QoTiTo3X+rtwxV9B4LGa
Uy/WR0gbr41Z9i++B9nnRVYjjLs+L1yJes7KJF+YkL+o6GnotCGMzeRaYNF37dp9
7gfpWFgGXhSpH3mG9ZqIhFD+cG8pnltbfuNxVRCN3UgAlk3cxNIIRNERbNnKA2yH
P2HPPZjV4OLHZPC1s1TNjYO6Z63dfibCQ7h58L63GVAJNOYbxXx+eTjgMD60Es5u
WEWFgZPOoiOpu+ZLKCef9QgOeerJXdBL0RLfCQXCnVrk/rCHeOU0Q8FT3IJv55GK
HQFHNmnjDk6dx9QsweAuRuPwiY184RQbQ+rD1NJW6LU3LyBTPCCqBpsoWoux4kka
jvH9uB5O7qkohFJsf0R+TWuIrc13NEqb8EjzxllNNcjHViGa7h16aW9G74DesmHh
xVPVmtc6tCGmJvAjhs4l/kJeYJry7cuhuX07FD4vPUi6L/JBzivewLimB+tTCJSX
3nlo3S6zCGfX1FfHZNap6Z4gZrGIuytQBPb8CIzQNidHNOnYZlznzWqKjigTtGeG
fQVz69TVUtBPRjFTI3gHlM6Jmp6YAywDbDYCP9wBhw0afJAK83Xhrrn2eUIZyBiu
SsTvBx8IwqA91AXKihtZceiTP5TYVV01q546P/9t6fXQlDqTrkOiflzhDBhLXWrP
NzqShKqQ8jUbQOdUXPNNjpDSOXFNzeDSb+1DlFes1/9XIkkrZ/ophA00XjeGfW59
yjEhyvUL1+nzVFP6csBhjvl+EeoFvC5R3I9jGQeAMhb61XnYUCYQ71XFBFlH6iu2
CjwGslIDl44gmR0OpvcQ1vNfyXSVYkq2jqSYuK1IvPe7/CVL7NhLsV5ltJbReU58
d8HIJH8h7HNEmcpn6q3m35Gg6ec6EiCobtF2DEct3JcpAl9zbyQ326a9kPxyfw9x
NN5+n3AYAc1BYXirfHFeoKu6Z1FGDlIkwGQuSL5y9KIY/EcKT3AMZbWi1W5rWyqT
D+WOlKQANu6w6dQY6CAr48JoOmbnP7937nM0YgSXICoqwh3nW4piLXxPZ3Pv3DBs
sRZWBMAFLFYiN4qly0a55sbzH9c0Mn8MkXWVq5HLyDgWYSUoj12Vh3ZddedAYpLP
JRRyv+OBRKOFx5k9Br5N/1v/m4e9MbO2C1Dbo01NC/xL53OZ6D3PIhrDITYdVv/5
jh081IIoxwVfGSooCNWkRwrwTjtSf0G3Q35sN5fOt4IBNhpoFmZ1ayvl0n9AOG2v
0KSSfcvs73xAw//CUsU9vG+3QovlF4dRWOJQ2Wp3yubEcrRfpM4Zge+oLRQ/X7/5
NS05faooHoX5ickkdaWYAgVHX3hmKXGsGyQLVZPXWxDKR7G/1/qZQgko16nE2y0x
xoxD2emt2W/H18UYRK25XgF/EsGz71acA+lE5CpQRvdivfvZzXTEqE6fHL7hjLMm
92EJiQ4Er1xvsKBuF/TZfnTDZMnJ0xo10UFlNjAio5OxJsm4nFQJVfZmnJqO0omR
Sqa/pK0DQkWl72PC0Pga+LA6Z/3YBGH1dzStbb1mglTEDInUF2llOL5QVIBX39ea
F+XlBFmv/XcaUq31J6dF6AgfbuelRLWCdhfaixGm4n7dZsYxiU5NU3eBi8GPchen
u1AZ8jYXAT9D2rGhBBqPck1EKBLxS7tpMo5Oio98gVjSNYQBaCfXOLN0ErM+RybP
B54NrIqEgAEaVxAcm4xgw7IFy5I6XSf95bdhw0c7h3ALtlACUeAp4zxSgZDqIiQu
+Eqyw7EwDX7xmwikcHfI+XZgffyniHCFhrINdV9qfl3O/BGvu4QTEacwqPjc69MI
P/SjBT7vrm47wYwJbCag9HttAO0pVpp9XZ4yFVEHqnCZ5xo+5qqsKv4bVvOMV+TZ
QJDVsY0KTY2L/o2XQl7JerS2Gvhcai7IzfDcTCbKm2SpDYT9wwFmZwtyWQVgm7f3
SkJgnPULa8jPgbi6kiW9djkMx9rPVFxssAWWwpxR1kAQNgOSRBFiZCaP6RLZ9txa
YpuqZUmJSKR14W7urkY9jnnf9t9WaFnoSL3H+g5BxTQAtuv88JOq5jqTnomgTIHM
iXypEyw+TsgdlP/F7G5j0eauL/F4zRSHuZ0+1a9YwFuJnrEMhx6/ucXnDJc6Hujj
Ii2gbOh9KQOB+aP7MPy/f5L7X4VPPyXHrdbiMtpic0OpNS9dQdBtX4UgaR+pAcE6
UaYW5M4fi8E+KWQIrHHWpFwUu+p0eAM2YL/QfhZZwxq7IBLXueRNvPHADByXNN8A
Abr2We8+G/xZsa6vFqwnDHxWCA5GqseviVXsIeIJcEtFqLyMheqeRGE7P4tqkSbE
jxrJpLQn8CKfmzuoIAK9LnwQ8FrIgArd6xl6Yy02Lw09yMLGT2Fys6TqYkODP3xb
gR78Nt1gSOMTOfL+eOHvE0ifrsBvBB+CBnBHbkTqHD+CFT9ZIZtPGj1tPMOE+JEG
j5Yom5D1qDtF7aynd15znYuapRqE7M8sOue4if1hpH6AP/vxRMU0Vpp1fi8Rj2oB
WjZ207p4BcIWx0fSwNrpC2JAGURz8WOaocO0bW6ThINNSv6WiTGoAgFjP/2nZhJV
r8xSxn9T7RVtKB5x7K0E1Oq0fM5sMvC/wt+cyhYcoY3lmDKYk302dVtzUkB0Yc3E
ANdboE3YAClosRboZ0g1i+edHdlZSUe6X+AOSkrBSPRcDJjQB9Wh0cr6I2w5vGYV
gtedNexdWcz1pR8U4vZFONjG03G2amk+bwPBAdBqu6QdWxm9QD56MmylISYf/+Pc
n5p9OlAZFMgvG+UxvY5y9EBFbAXxgdPjXSqkYRVPQXy3S3aes9jqdxniY/1CMptg
h2crx2XlA0vlU0KzlQMw8iKBJPd1T3g8SMmG7Z+tZmo9Qkf63F6canYWK2jLoJjK
hsaBCzNTEA1cQzSgY42QRqpvdy1Lm+SJhk1Fsp0NTfjrPzrYsC+IJ/IIpRVUVqQG
xIeWP2CVv/c8khm5SMB6X59OGiloAPgNDuw28Cy3eBtZD71KgRaX3KE919zi8LNI
lgMFDGyYjB4xT+aY3zd3GBlTE13XCyW74IQrRIzARLjnfl2axGM5NXtQ2URf00PZ
ZvfBU5zWWNuCnMhB5c6W9bXTd/LgGK3zOEaw34ZpXldoJoNvBlo+aqSnt2yfBJ10
OAzcXrmZQLBmA8IGv7rD+LAtU8Vq5H9LDuoq6o5Sd473KqnBmL2Ti01DFyPp5rMN
Lp+wqxrI171oSLWk4UPIT9iZbIp10VUIIFeM4aL6D8CZInSdX3dp34Xad2sJoxYN
rWDBnVkg8QpdVwl5u2Iz88Fy3ZuhEUl3izMUtaYsAHD374klzIiBfo3Ei5bj4t9g
vePcDriEfovFiNRHbFpePEy+eNTib/kWDPi52fc6rEN7RhIHyKK3N8oeaWHRWb22
GsltHOeVaR7MYlarhu+ki3JyRu2yb8V4nAWUoChWX5pwsQ15BMZLPpcXYHqxNosP
/cu8qVR2dBnSwMY6glZhXMxxZS1VeCqTcs1AkRUTnb5Z/+eJiYQJ+N9iM9tf1Es5
QjxCoewCGmxf0BsykoQQ0ziAdwvMhdIacd68Z1WeRVShnpO9Y+2sma891/mEORrM
Uz49yQ42g/6dIIEP9D8YpZyF2IsC579NnOADPBhi+G0l4NQqdjmtI6HM4oGZTSrz
ig1tWnMedg6iCwUcGmlvoHJfb63cwteKrG3+y3lB1MjUpTL38ZnDjVHX0ZkgAnvP
kxTHa7RodFwGM8aRWU1P9uvaRfGxd0vuCh5kt8FBYISbxkoiZD4zWzXsk6oBOR2M
TbdzE82SLBoZmxjjr6SKKPymp+DRw2HY+GtPjzJITT5d/yR0QexafJzLpqDFBzR8
reqQ75RW4ED5r1GAp3fstXZxd7BUDARiigevCMYTTqhP1NHCXYBvNezWlaJC1sna
LkFE+EmChG41breOqpPiVz01Z0WhWd3lX5LlKQRQ0+Dfvxl7HCCb1q7stL4L/zoO
IgKHWGLVBiVJP5xqI9JHpK2i/cuHaBwDld9f27wRv1zSWZAG/nu1oMLoSfB6jrSZ
1JGAuI3twMSJkTpmZQP8V1mUZyQvKfi9whsqao7212yfEHqVW1T5BjUv1EzJTYXS
WfggBdR2rc/6C5HJUhS2SZKAqViAtn1CyZxwGa8nAVG9FBloRONirmdfRJAN5pUr
M8XlikVVr02ubBnjiIAqoE1KyjAT7k5LTHXXU0uqntp7gk/dZ2kq/hvjs5j//LZt
YaIHdU07RwRpEPz9Fcdy3Yz3wRJr7oWlA/rKGKTXP4nMUBjU/otl7zeFfxKC93xZ
P9ScpfeRJS0x1gAYuRooqRaQm0Uremxn+WtFczP3mkT5ZZyO4NhL7QzhXa1mEFVN
mylLoAmL79dkyoaivQmIkisH6FVNbTmuqbuut8xVkVo0t6wZTsriSRzAbO9Tub+t
puvqqpEA1xdsRQq1I1yga+3Ffay5m399a3EC3xr3cI+onj/2+ty7xmD0UKNJDgVX
t5U/KZxEvlJyFZ4MsCwXaZh+xE7hqM+oAcrYGtPT3Y9u+NO3r4Lg/7pc0TR9nokO
xAD5Km/wPqJNhy8q1gemaEchcHmf1VMxcncx8lYcW8e0OicGAfOE73l7kR9t0WoK
vr5rnQ47xfXkljjAxzSfkxdOfuRsFwLIlEt63MqnFfjWn+VIniNgHW9HZHvic0nY
7pL1ppYlHnLcw+1WMaIBOIuOCL0NuADWRgx7fGUXxeGTJBQEBO2IE8i3ifC4SjyS
w1pbjbIxmB1CYGJkQ8bNN25Xn9Z6VlhdeDLHUzgiFmVrhDkENg1JUY2+kyKlEJEX
GGa8BiTmjZMX6/THisgYukk7CEEzDTXpZcOOEn6gEPacPEY3EoVXvti8VsEi9TC1
dLjLnd7sZAfQW00U8fI/sm4nahzpvP9d5heJIdIAhOZWrGDs91T5kOxX6ZkwXlR3
5sZDSO22BuAL4+SLjdtDZNY+83cr7S006q+YGxT7s+cC8ZSoGyy11EKadbmGPIWp
VkEdSSo5u1gZ5/SGotcbImoz/nZ8U9QZpS0l0Ldic/PHKS0iUZNXOhffRty8TsY4
lzy031jSWNiVIQm73rGWQv3XAV2PH1W9TzaWNaOtoWzsXZ2io3rx13ZwS/jADo3H
TH3zcXYw1upHr3p500gl7FSZVVDdxt0Apa4ALQzsB2s178/LqUxkRZ15cKeChMA2
cbGKRql5xywO2oBKPQRv+o7NmQM9Jj1yB6ALGv8FX3K4Waqig1xIuL7b9RJsfo01
mhqKUBo8BLmxADTuktFXNmmJr8JZeUtr4juW4vuwE55bE1rrG5fajZY9jAIvHlLG
YuVnmahepltLjLeALhFPxlcL6e8hcWg4O7OQ/ou4y2nHM6p0C7JV5dTVQfnfuqVV
/rziEMfPtpUuWJj4NxnVFfA1Q0kB40uNVdC9L8aTyXRg/aViArrh079r4Zxmchne
Kz1L4ows7xcTIXpKggVD74I4VdtEr0AEUyB9jQfglRSHquMNgWhOwEaKi/mF/cof
xlQDTQoccmKz+sCjEgVCsHudscos1KMO9P2dDpxzNCKqvxPMFANbOxXv/YKsDfVS
2ePXF9PDRM8h9vmpW8Y738KrkIFKMEHM4X+O+u2MA/VlSdTKy3xZFV2FHdMYl50f
DS5wU7tOykzkVfqCg/8dq/2eQUJ8/wEt4/qvxX5Z2VCqw0cqsfCqW55I9gGsYmwZ
q4OGwmGm6Nh04+Mj+LrYwhCXsxji/mu+VFo2WA24eYI/vGs2TK32KzZ4R6VMqQEF
Q4bVkK39WhtiUhXz/VVzoRFnlN0cxMggn8EAAFXksB5+LXXYu9eTPlSnN/Ei/Ebv
yCCu4pMpjVlTa3hWpdC22SyMBPFXHElDrDekymJSFmGZ9OWMD6dPScZvb3QP2G63
AFjsdScOuqGdiZS1djkOGCQy/NbYnP+FXE8JYP4GrCzZYVgSKhqkFhBj/h9Oiq9K
ywwT6rB9tj0iC+y/sMh50ftMzxMzJlgMZ+gA+IOoPcMcvoc1QyhX2vUx4m5OEaFx
MyHO9NCtlucpkkep4rioVC2S7MR4p5CUJRpNUgmsYRFzMGCG72CewPGfQelafwiS
4h664j40l3ILUWdOI+VK8mmUVnGfaoym+nRbnmL1ET1Jqdafo177qBE43bcU0vb5
4E+Bch9nGe7BMLGTlvDDU5WSRCOKdqc4lSeuhZJK50l3ZMyQTVU7W/La06GBfeg/
OG9p1gakDQ1cFoXBWPJHhqBrbUkvDk3yGVaYq4Pbxy521pXabXeVhF8u4v/CJV+h
KwOibBgBKbMNIWI3cYjMquzAl+hPe5jGtW5OT002/liWpBvKWy9jX70nRmKBIRah
Y5ie9Pbb7QW40QKn4jqjG86DP1E7X/ObZtkYZMczBoskeKPZfNnfTuvrqBeFQug4
AvPliYajjuLkWYIAALv7TcWdggqWu7ceZpLuIpVPhqYw3xVik0ZY/KHMmqxfy1to
kD5k0eJ2WdSlfaR7OGTRfBWazlTfDNg1Ap0lmQSkg1Jql/Go4fO1l6zZL944GTp9
oKFtGdbgMwsqNfbzEwJkjOAuOO3eTua9ofk0S8Cv/lhAoF/2W859mwfoz2Xp/qEJ
+ngjkD2PoIzfgC/V5Sgy3VyILawDOmyD//GTfG5BPAXhRM+Oy1KSxODByydzmHGZ
U/yUwgF0XhhqqJsSl9u9SDlBpLBmuYpg0yEehsiaQRQeIX2sy5S9deiYIySoMjgC
AScVLErKBtBScqCkpQzEhREXAAKbxX7TBEw6BuZjp1OnQwyAc4dGQRfqUQYp5qgi
c3u/W0WZIyjrfgT3N1vt3B2jjvy8RXhvGjUZy1MW1i5vVg23i5T2XzgN9WFveK3Q
j+0Crhj6B6ryHtUcPrFRcNPTAbauYcS6d2W2egvI+A+kPAImp/O7bEO9iecl/2RG
NKe8h39mzx6NDxg3F+uBYC9LKAEArXSln3iNeeAcTjXg0xOSr1CLECnTUNBUIEuL
zbc45O25ji1eN5Mbo2mKhY9AHVNz3XQ8ynd/kvQFjv1sCYCz4q56M/FWVuW2tgyI
zI7RfvmvAJtzGC5CSeHYGO2KbOGTRAhmARBgUemUELfhnOk2cUgebQg+KSM0Jb0j
zZhBt1raYsdZ/x191sP2Np8W8xaWN7Dq1IewR86LL+UNXQ69sAcY3dcWvp0/ZVVo
GjRzTR+3N88bEsJW10vhtS2LcwjZBrTPK2T/s5EmNPLB5ssHvQ2FhW+rxBCF95DV
+JQOXacN5PmCrJ0hpV1oL4XkxvqcO9cvzQIrfr+6pNYB5BRPkp50ubTwnr1vNc9M
Es8PoHH0cc4XTnAkmZoKkPLV0cpmcmciTK5mPsK/+5cC+ygb+GhXQ7VyiXr35dea
GQBYjxvaT5RyLvrw+EK0a0Lxe22dx0vJZf/R0i3pcxcPDc50yZu6hydzrtq0F3pa
7ze/aNcNcy27QquGjdfCbHUoWfZBhIswCXqSoMCrsHi2FXR23rKTiu78TwWkqjfk
k50PsgEPoamTrhFWwAEjbpxvdYbvT5Z/DmKK1Fez5lOWVffDdJtS/7xXmlUmSxQ5
SOm0iDoVo2YXr/kiPCe1MOTG55v+oNlQrr+Q0S/dolukA4OHTrWf4jzogA+LBf1O
s3f3gtl/gInCdxGKcMu8/zHcyaQGGT5EB8cC2z+1T+bt9mhiCljoIgpwjb1cLSrE
HRqKAvUTyk9rySVhQN869udgVtVMo9gFuWEScrjCtvisFDeRmGAVHCpbXC9ichbm
62BpXuVNLPqd+q19uzrQAVSAYHYmdy4/ZWzovXYt9ixmmQC8KUCDPWsS6KG8tZtf
Sq0KaL00ZysMAi6AbG/ozmEDB/RLjT7IbCENwK7/v5Dv0Jyq9EjWhlQyHAXERaOa
sGTZwEu8nWyBonAjMe9d9xLZG56jvYrHndeo2mYB45SzeOgeEJKTHtRuIKjhvFji
CgfwcRkB5qYSGL/DfiFzVaw1i0oRl7KEMa0Sn/o22gCRp03X6yBH70XBlx9b0ATU
+M6Kzptn68laSOTQ9QnVurDfD/miTMpX4SH5Fj414BBb+M9RcWkITHNscJt8e6jC
AP8lkeNagqvCpMo44pTau0XER0vDAdncs7z2xogKp49SFTgXtPpQ7XjlmWfbS8fh
z+6VJxMteH7hHib49RAl0kl8QsEnHzaR4oKjW8Amn9cYqK8ZiPPpcdWwi9TTZMI1
zNtlKVgBjr3UD6vTXiMxajrYcMZS3jS38j5OuCnfqRDqTiimiQ9tq2bDMTFUbypN
yhmjQPZMk+ULlJLcmhQFs72QNAzEZpvC0V1SX1yJE5uR9r/B7q3L65mFoRXhmJuT
9ktvr/oqt6b3/PrgxWewAWch7tp0B0A2EEoDyZx3my7+5Wn7EcZYlPHu4DbwKVpp
OvM6e8luEqMJbs52TD9K4guLhfM8jJsfnG0us4MUYMTfaor/JsXXBxKETeyJrxRM
miWIkC6nlrQmX2jeoKr6tFxSw5SEcZyfPk3XMOtTLYKVfVOiPEDVa2G9NieTZttC
HgMFsZPhW1eEhUeXvmOVbOb7VN57bXMfgbvauA21J8u1KVbMQkPaQi1cfxaVrZvh
WntQCKxNxc1Qh8kKWb2BWz13qI1pzaBlnKfHVr4Idb7R9S1acir28Rh2p7Ett137
QOYaJ6P/mZFwMua2sDqno3p9UNGon8zZ3tlBh0IolkELpW8P3bgz1aM3Azj/STlx
vRfyRcxfVlpoTvlS46nurShkYlPU3BICuRpR8LxsiZ1hdhL6NcXDiGoyEFhr8mev
9ZAkPyiPA4aUetayq8Aa+zjZIWlstptd6rZUui0EtrYhg9oiNfS1afT3OucmAqGx
zZOGXc2/qf4muvjyvCfy6NIrGSRWgbFgBeVWmYfGzcBQ9QjvT7PCLvVi4NzBD8i+
iTJpRsC1x6sAEsNEUGuuTFA+jGgLlQDZhLTnwAlYMEFQ53n24S1g29S5BTSq5p1W
yuPA+kme8Y+P4+g1N/G+h5QfLE1lemRo1rBrvD4yuyMQfOUzNUJoYIF0rP8Pb98n
zoRsHV/3IL98xFSC61a/xqtnHbGiLNlaeKKvORuwn5fJAJ/PSCTMIWhdOhOl6Y6N
LKE+Hf6SGFbjPHS8mIwoSp45dv59f6jLrPCIMaSxMxQUOWAEyKC78kGt31YRQ6Oe
/sMgbO6KKFxooD72Q6GYVDaziFxbc3qCSB7cUS0V+GmPXT87dPo7mbl757IWpG+9
sg0Dk1WCkwIe41tD/CXcOGkmsdHDyu2msD8c45jtuiQMrwFnYjRk9SWUJonipbJ8
RKXZRAZQ3Ib97kuoOTSYxqnCfyGbOOHz3rghbNDzXL32uIMAlLB4vWK1TK37cKm9
1n+lZsmskI1tKEctXPGYEUwDDkB7x1jtX2opnpHGSnq+y0M86sX14RqV68T8CRDn
nfaI2mgmJ4feU9CbtI37b0MSve8WbMIrGifyBc8bS4PLzwK/UXX4VBBwVt/GfA9N
7zV7jCW0l2SwZQ6sni3TQXkA1uka9cHlqC7nf5PvxElFabTOerCgIOMf9EAe1x8R
LamOqBqtZ9CfLUhgytbgOKPwMW8aO9mfRaroajnIObcb45vJHTVE8tGxMkK7aXp2
wtaqmLHbOfODETZJIUy9XsEj8upBNh44zokfEe2e5TyMeVNwolGDrdCDOdpAEovl
ArfR27zJbY2Oqyt+tUc2LQkLTw0c5UicEV4sIbxBoRBkdTLNUw6Lf/Swdx1XwIV6
Rr+KWpcqlqcgRmaSXrSJEQHyMRk0i6LX5JUtkN21NA3Gu0F6tndDX14b1i4ZMsvD
rUE8flZVpS9qUXUaVW298ojhYuZKY5ZWOt1fxi8qQi2l/ivlY95wzwMZDBV7KKFg
yCFmy0CctrALjkcviRVRfOWwVDtfqVByYmgfHiw93E2w5Ht38ZC1notL0174NMdg
nnN61UboJ1nXjtuMnbhpjJt88ROyI5/67Ty9juJXHJx6JsrMffI3U57kDPqnoNC/
yKvl9MIiErYP3VEOOWMVbWqGnTBA3Szbrq42JSib5Fa2SK2F2VQFFgVcUosmJ/1c
YZbLsQZxjwiDUtGTqmSwcvDhyz5BPETvAc4eGBijFMp6BBCQCo7i+DoYdpMhHaQI
OeVhhOuYecMemdSvkLjiHcKGOkPP8kzE7KNo7ZwdW1tFyvYkAufgvwWC3XmC5urr
JpmSHrRisLQ4T0RYTzCvbtyMxhUZK9EB4thGt/08Ngl899ueQTS2qiBA5EKXc5cx
itIPLz+YtDSp1Lh+seShhnrQA7Ei3oORm7tRivobZQxQWTE0Bm2Tyd2LzNrKmT1+
MFUlD349Efh5QSNaV+rqlEhIs70/Qy/7DYTcygIBySlUvtDngAw0y+JPfuyh1Dvr
4vYfaIt9OU1fkAcVcKLgG0gr1S6vgDgzgPWggM4SAOtYlVEP/M8e4KmMtzZHBtK8
CJT3H8SxeCRM3oZCMp6Zyl2q3okUqPGu3xbRL3cU75+lKpLekPKljMI1sowZC30s
ogTI83RfrKLcqwYkHH0467SKQS5aUhNgVFi8FKEJalEx9EEQvDQiNFnlTVJipSoA
LSCa20fxBjJWzeuD6UqHmHn38ViGok1Bc6iayw3SkzcmYftZkmem1AFHhxytf33S
PkYDN8ekhpyOPRcEy72ggA+FS3g1RBVkwfKe6QaffT1DwNBPAmocU30slagwShYM
9zMNWH5uomRAnyxaQDX5vu9CwmHgbxny/zbVz27o6nsGPlYlvuS57hUW9QigKnHO
nL1O/ssrrUjpG7SgAr01124MkVb23cGN913EYcEb41z7yv8Bp+zwvuo2E2D1RmWc
eraAD+kMooSayXu3MyoY9iNY4sbr1ERz38sdf+JDbYAtlsp7b7HnhHqZu5C2qCWR
L+whAxBXt4bE9GzB3PP3Ay/ffdk77ncQArux3iM7RQFL12+87fkGEm773bDFVPsE
MpM9nHKHOqTue6QGAPvVydFxnrDhwVkXaPeS9EMonM2Oj3slNRrr1NggrWlyoQBG
tkErrSUl4zr6N8vsujjhT/jWJRyQabGOrPoHCBtyyiK+P1vvItuJrLwdS4K8AA36
G4tBFwiJrg51icqon+IXo1YqR35+nbtuLPusptsI8wLxyeG9GeV4JsC/ihxA8URj
3BSW7O2vAHXeiSDVhbLFbOBIMDqBkK8WM2H5Ep5ESkrD59sZkbUGd2nTU5usrnDF
gPJna9UQtJmRBPybTlTfocCedMZCnrWhijcYWezRTb5cZrqtx5U+kcZUlRSiMWwO
9i119U0Qnk74JkOjCyBSh1zSgN8gtrH5TN8lL+FD0gvpNVwQsH3hm+hl47Mp83SP
aSpVUzAS1/hVOoXdMYoQLTWryYgxFy1nPP0Hu65G7mE=
`protect end_protected