`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 2800 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/9huKRhRMtvnNqb3Z+UU7TahEoHV+T8U3P3ufru7l1O
3DlgtZzb9QxCbOjthp9+wDkjygH0eUfDrEl1ovhZG61RQ3QgeWgro9W/wJKB5reL
B11y7JOR+9lNh84rxPaNL3tI74fKVH6d6C14ci4Lo4bgv4A/SXqc1J6Gu1C355IC
ESvfjHwD4/cz0yQynffoMgYPxLIxxQ2Ah4sDml6lp9m8XogNnprukCIwtO3hqlwm
Y8la2yvFWhwrzoFvz70msxZj/5v4tqpUbbdUKZI+PUgsippNuIYmn8ngciIQQQ40
RPjITwpBGB3Ut203E2oIaNqvv28wZP99J1Sb6V/q7ENQw4lI0mlrofuUXsgUJ04G
Yr8F5bYqqMsBuHkSX11gQL4U9NOFzVd4MVTE7pZgUIeUGLCGT5wnISsRNLA1H3Tn
inHELoi+QjyOdhGM6kFIOO1lfg/RdaIab6DDwuJO1l1XyyfpKZgDv0Qa+7Znwtqp
FJC0jO3b4+dvsiS7v6mdDu9GUEugxD/gch88QVPSYMqRO5xg/aeQcMy43rDpAzVr
+7UsKA1zzMo3jbr5QnwPTwtcTanzIpYPbiydQMFhhGztc0tCYVgcrrcYdNQ9TCYS
tKtob8xor9RNLQN1ckVNNUt69FwKh/+ZCSlLfPAIIcpM5WIG5yB/nv3amdRGmuKm
XuPqzPYnShA1BhdgsDXUgFYr6tRM6+KsJQFLGiMBioS4Vp9W/9ky6ud1j/dKhItl
+muB3q62s1+NkfA0i9hc9+vTF/KgZv0aetaQEn6T1KN78cnOhVt997/dfNiEDaK0
oaSb9LRcKLcK6TSk4Vp8KsPbWWx6Qcu+XDu58BGA6ZiDv5l/jSikvLzBpY4Eit7m
VJMdQT5AIDILpsBfbFFq+PuLO+yft0yqvCP43i307LzH7jQeEINFIbNyM12L/okw
ZN8SCAJPZON4Qc6XETiT+a60CrIYXKpu4Nf+XP5CGherhXggB5D1SGNF7zuIhGHh
omF1J1GfoRsW7678ahgu7HxsjGDyW4dTK9V2BqoRJzusexjXufkzIr8vfNFE7hHY
GorzLLJGi5uP5W1wYbya4y598hRt7aF52uF6/AfMdKL+qLCoPy0UWSY7kPJ7PGR6
nLzYgWJZ8FQ9T7Y/VcMH+GnktFbIGjncC8F3HnULN19IiO27+c9yCudo9dty2mza
UUWJKP0WH01yT9kD9iPbA8B9pwhwunOgLF+3bjGM0POXkg2j1zg0cf1uuQxtyv+J
TNBdAqHmtKyk1Wb4+jnOQZtkdVV6RFfVaOxj5bzyeITqhMKuD9CpMs81N1C0b6lC
ZQ+SEbQagBLE/xe6wtzty1hsHHzHh66dsD0Dt3Ztt/3grG7/lNUGiAoeC9N/DS0C
jBylgsMprMXQ1A5Qsm3R9kuAeUISihaDpyeamMQ1PTGTZbbwVxwSr8ShKbUn22pe
FioEuAufuyjFKDYVs3WQXzN+jDmPSvfI7FgsyIHQwvHfB1kX4E1+9hqbAKG6tuHi
YpEoEIFpolHggHrob+pk1pIbfgACarQHD62IapfL9DOh/Z7nt/rIlKR4K9HQgaeh
hVd12HnvnKWWkscQgLB2+TcEm3ONZZ3TktoF7EXOBgngyAJVU1G2aV8QcomOeNrn
HQLjvOOJncl4xUZ/xh4tEz9QCyUbMq9mVFDEUOKI7HAukw1CKqyySRN0GZoXI4RS
PTvq5hAhfFld+IVNBlYE1gRJwG083dCyrtB/o4z8Kj4jZpG52+BUNM7EC7bMb0iq
r7iLJx+GNg/2wO9+5kSdo6YAByQGbbXd7lAPYcWdNc50mvgHl6SDQWRF0wNvIhbm
waS7gk2D15PX8AlnX6sCr1mu+KrCdvnLo3LEbCQRVf0JXnmWaQf9n4pHv9Eb63O/
XhfCxNDo1KkHsjRxjTYUKsgX/HPOBiIlQ7Ab8UEAuVuT1LHFUyI9ZCyNG9Z/hlmk
T5kGXVjAp+DZX+5XSkphMp8N15R9w5lkrb31mT7Z0Ibf/m8t3Eej/BvycBk2q2bk
oAPbvtTzFCodiuW5TI1MMREta2xC/uJ77O8kXdD9AZDBhQ29IZhipLH/nlr5yh7F
BHQkATCj/OMuTa67XLsiVb6aEYqcOqBDwkwuHqMXswQASKjw4/sA919dyCQeA5QX
Amyndqc/mgG94JgA/pF4iUWw5SqVekPaldVwFeGWyTUAzqqUgX0ZpYhalg/5GMST
5bfDrdlDWr8jKSV0+S1xZ6ulmveSgEwpZODDBVg1pZlXQSMVKsOvX2CJXwIFxQGS
lBXQPppL/0z3hR/VxGal5zjFkPwyQmG56yTttNN77g91GLP0OenhrJUh4UDj8djN
LDUuk2ifIa/6CJWHMEoajqaFl0lOELP9tGF78k29l/Jv+5WwGR6T646yBPy/HGu3
w7Bim+y6heCm9IcGUoagJj4i9K48r06wwMwk1QM0bmYYGu8VMcnewVqxBw1pOaJ+
fCg9viE+7TuDoGsHb53XyQdkjSQMOCOhqL+ivToSWfBK1FuYaWRuRgpob3CADRSw
vzbGywRh3IOi7m3QCVA1cmfvY0dUQdpLMad+oIFlR2PT1Db0WP0UBkI4rHm2LT8p
eCx+3eyXJMLUqop0hWlXaDlv1NujiuIhuCtqcjOE3JTIy2OlRvafRHcB2aVnmhsT
U6YMTYgbq6//izzL9nGHB8y7axmgE6MdzYsNilqQ4h8RTaBlE33Nh7rSGW2jR6Gj
JpeclbV+zh8W/j1iRzUMeTjuc33P4swpk2oa90Q2LMB5WtOsiQf6vrqBik/YXeRr
fDzVvP7LoMAFizvaPhh/cfGoUoIakl0zORKakKhWz+f962mYQXpTWyJjoFNS8vhH
OJtcD7PzSEFyER/4ytuGboZ0+LPLl3sPJ6ce152WT0ZaAGuQ3vRlvotevE49iWUa
jot50Oe0sengmJB2JwfRgLi7qzSqUuWBfLyaiLtIPyMYoEEJDpAyQjh8K25QSSRG
N8VTb19CJiRGaQqx4e9+whQwbV1VBAAsrQNRHvuq8K4zeW6asdBZWlSeetfNEbah
7l2qB8pvBLiK+6jHJAULwbKkX6U3LGXJpXp60Sgk9Wa/bh2fhGzvqGb8ZFy3vxxD
s3g/o8joVdtDXGjZz/RGkaiL/zGOorE931GkO4zPjogr4g09KboPO4Pq/2qEH/hK
84EAbYxUR5T8HD29AMibZzhechCInm77BGuEHBp2o1OrrpxMxgAfS6iBGHGFd673
OG8bfn2soc3lL00dDgelJ36T2IdbhHx3gH0VMJqTq+lgsk2u69JsUUjYkfzf0eAM
OJaodXAUlybUcTsOaGWu7wCc22KKhJfY3uDNnRKBufz8eOuE97/umCV1cAup78pL
Nsx3rwowMizGJns6Qwb059IQGB+7yjkJMIShzQ9o1APwWNCb8ZuSbZPzUIdh3fWk
r2KAvov9eUqnzuTk0sghAWj9eRv49difWEOG1CGLssvo4DwOftZphVVw1bn9kakY
7lj4wfA+SkT8bqnrixbsZZsHrDaFj4NqiCQahauY8Ikk01C59yQCMFsp1ZGS+tuS
uIqAlrOoqows2lhTAGLaBkhuWZCWbZSTnNlU0NygRdODQRPYA+OLmx8n87KCCa9p
DNxds1AfMGnsHqvceu3GyjERNTW7ZV9qgLxqUgPqjJTkbUsQT5ZpNlygMkA8ddQs
a++9pTc5Zqi9Tx8DtRnaDg==
`protect end_protected