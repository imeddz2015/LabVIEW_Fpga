`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 13584 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/59UwEX+aE7FohaWu0/8IpTj7mav863zUNIsgIH2BWb
Abd9opeuBjbGF/waQMI2vMJTwD1ie1YueHc3nSNpEh4OXp8P5ybZFY89uyGz3ztU
W1EsuUnchJoQgbHZ/sLbgtGRgsrAFn+ZoIeGN1d6RAF2wAESJmYP8zw+p00RvjZ5
g/irlrcvR5923+bWtjXsf9FIiH2yETDkZPKxXPvX6Bzbh4ySNswhyi8nLp8SgpFX
zS9w+wnw1WW4nNh0Jp+GoaPbQ+RMDg5F2EPIU3bBJmHN01AA+q3DA0mxYDzIiDyE
H1uyAtXUTn1SSvBQrxnK0xZb5s6Zn6YwFF0tFyLdJ8pKp90He8Cokm6o0yDWpFqv
v16F+ue9GuXP/BC+xyRqqh21ak+T4bmo0LrdiLX4C8W6oW52gh3mn4mwKG6B/w4H
mIvEXPAqiDija52kS8KefkmmwzxmdoNb2ZA9vYhl4zVzWFnVbN82HX95x65ckCR6
5pNkCgFcUFiaTt14Kfmt6N4PLEntmn3ADvXTJyLbgpyiIaA2hb/Ihxzj5K+KeaeE
ekJj5rCC9mwV38CI5xbpxwoqyCS3AIum7y716T2ZVsCOx3B0zFamKgOSjP8jJ/oa
fYWAgqZHRbKmRsXEld6FefSflifnIuNyJaGjnwhOPSA9aefUPFUS6zP/Y9hol4Do
tKfpNvU8B0vkhjkj02YHYXngwhv7YTVgP45tVX4PbcmlVy9Y/U4uqIVaMHpbyCuz
D+L3WoQJR4pcUYk7/vVXoI7M6VYoMEO1AKg8n1KMqB1pNb+7dopqXWjYtUzIEGpk
Wsrq+jVQ3oOGU2KsuiFF9raSPKsUZjX2CiB8MVqAAFLZNGywUlp4sEETqCBIHaUp
KWRGe0Zcz9TuzC57floKnZ6bP/+pVHWIKCqFAsokcV97biEccYqgj7GwxrOKCU1Q
LG1gZei5AgH0pmddyS3Gl90+imDHY5yU8k+dC/iZnEmKEiGTATs1zqoY9AFqx7+F
NhkmLuJaaVj6HUiOKLvlPRO1z6qY+KpBxuIp90Vmqc8e79qljMPUVJp1z1v6nfAb
9WA2anTY58vIhvl0M9zNmYrXU4xp5Xu4bW3pEINTDg4vZ1g4Po5VhNetXNkxBUz/
q91cwtketX5zC2XZ/al4VHT78wFg0nptwVCWwhdAJmMGr/v/mK6o+A6qsvyfoxwg
Q/dd3pqgrqvu2+VwHbdTnqiBU6iHDpvOZAItrEX2Nc2mzEktZ8G+SiAxi9RuSfX5
gJyJNeaHn1q1CPiQgh23Twj38Phm7IMtwYqd3mw7WE96vHAzGYOxN0jeLqt8O/a9
8TARUfBLghSrt9cBvdx4cIbJAlQqc7GxrvSA+wqPVLooaPhvOOm4K9XmL6++OZHb
JQakjDpoCaXA1slNxS3KD8w1RoD616Q+GuU8FndzOrDl12YB3ZBrR1s141A4bzkS
UO9q2dBoblD9aP8F8qhGBpUwlPnrXaQAR4ALAfQQufxS5pO+qHDS6uZeTCWAaXgA
gobWXTDBIsw6Ob9dwEuMdiKuwrR5I8hIJXqpPQ7qIlzkNe7oEMOJn+zUjyd0LZvC
VVtuxeaPyO2Hk7E552lDhO2DYI0fbdAZDaIopOzdpHVlMPwEY7kX9ho1117TTrHU
uoz8RQ2zRL7Q0SQP+VyVTuUY/aRIys6fS+dly8bGY6gpj5Dww3yPZim0ryTeiH9G
MJb7vwnqVGA4B9QUDbmBGwjpLJ1rtkqCoa2BnIfs9V/swVJwrTWQOexzZCFpgZhg
yM9GdpPeDLG8rAFz1hfweyIVPMUZf8wZDibUBzXc7fai2cYzbAxqOwVM8/pXkzaC
Z8dVWIFCe3S+9Aap2jQGU2mmNGPT1bn/qw7GVpypdbexhFa6pP5RY67H+o00lGtu
MQTNhoMmJyeAnzbQZ5tE8VA37LlM4FR5EJplOkv8ZLGcwVCbUoA5mtVrbgmxE5rd
68lhEfJpVvFT95QfhpimHGYVtGo47s6oEA1q1dpADUkc4T4+nEvAKsHLLFzHi9VT
WUpSyvCE3HyHHhrkCJexdVx/y6vT06RxFGkNopJDnlmx77INmEHP/CpAEUxjeo9Y
jDCU8rGo5ADzGp+3LYyPct875KKhEknkUmK0d2aU/nVoH8xsLigA8gR0873/pPG7
vjNAwBYkVNi7a3q/lmn+ZjT9eV781qCQcZhaFXzB/HmHXHokf5+G5GGF9Uw+M0bW
+7PKDGzNgc3gXP5oV333CZgi3SQNxFPi3qmhNZWUKoRm7LD8Lx13xsKtri/Rxp4X
M2tPJ01e/5NrIovbMvvJCE2Jt4bzo05v8Ulz+pUHVv2ia87RfDqiGCTZMQQWVYe9
db1aI2pEHjp7N3l9YkQUOCyezCMjop4Zgxq9hYFRT+DfchsJMKHyOFEd4ix2Uz0E
opPkDcsCsmX+PtLB6swyJizeWpt3Cq1EpVLXsb0cHDEtHsuZuux1v/0/6tL2lMYq
0jmoep4oIw7lu4hUe2UVvJABlyw9f/LsOGhhCspkGcM8IKronYt9O+WyQ6wmeU4j
eNrnHyRjb24GI/rwoF24QjrqfpbqJ3lwSgKxmc+oqwUjJHjh9zLqhI3CnhR4D7gY
0IRgMN6RcH9gDWaHVRQ4iXLZgl4/fQL8TOFWeijOYlzcXngy2y8UKsodQX22+S81
nNdjwqHQYiO6SJJIbR4HjmJ/727PdOqP7maYeK8wY+mVIFHZxChiidxSrDRd9K0d
Rh5/fl90hYyq7UZhfLLFYe7RcBehn5Z0+/JkDcO/LspPFN+MhJchaYhNRcE619vJ
WP+frhi4lU9iCuHVYYaqWPamBOEMwX2MRFpQz0fuIz3ECVg46sBq/2SHQfeAZRvK
7JZOX6Kqz54KdFXf3v02dJOK3bmc+wdQmyzDrhZd/i3UFSFm1o4q3K22BoGd3bb+
4so9pjukxGbp1mCUeHSIAWh6tvnIGrT6fNquv9Wvv9a/tzfl5B2luEcakmOGc69O
hpNfs0jYwyFfhBoDLevlKGgjKa5AXbMWj0gFmL5dSkX7QwnpswpDeWULnFYiQpkB
mYDCMRavqlFxbidYjhx1QygvpiQ1roJLhO+KmoA+JiuItoHbtKJxCfuWR5O+p08h
0J8zF4dpGBLU5dgc8kbB5xpjurX3Uz29pxAu6+nvVHx4VPubiLwNWeZuiEs24IC+
fraj2kK9vejCikyZfuBE3hmBJGoKqgdB+OQHs6JU6YDsJYRmrdugTDy/Ay4oLhyh
TL2DFfnyneqZyRaRSWHF8Xu4KSP2I4RKyaGuXgWgQK4rNGSYvLMDwH9e0lwrEHLH
B7wtJ6o/oVecKkRniJoLP1k6pSvxXIjlRWktBBaJEXN3hLCXMbeI8s34cvlfzQbM
BbHfQm5jjw6FeyxKfcRt1V8jSNh80wWYKTJUUYmd4r2Vr0YuKNZq52EWEfhAqBju
Nr2VmyzD3wdWUKlnoncq+w6PAwZOhZ4xHWHMAjbTTQ8PND5i1gBRJqWezqXgjfwb
06pfKq/819ojsjSRlEXB+cXy8pEvm7fkAWlK9PwiwTwHar0xefgPZJdb41k1b1+U
vlZl3fz5zi3tT+VoY/D8x+nuo5QXZmv82rC4iSsMZQn62rUWNDw9LT1hNXvEOck3
qA4IkmqGUADTEAs7MYnLIzuCyYaT5p4kkqbUchmyPuzR3YFX9C/FdGBYgJgia7mx
Ofcreq8WO1ftqEAeMhR4scl92UKmVgL2i378rFztXBfvtxQJhuzYZ6OPk4sX62bR
+ZL96HlrT7H+O+tgMZIIYYjeDaehBx9eQCHDnyKb2GYK4YTmiZfQbm7WbN//+o0p
E0CxCHnuxJqvXlZSGzmy9/IBCUhMgOG+iWeVhCoZfxEateox1qZk3a8ZUOZvpztD
HJjROaS1COubgXKHURmpKr0NRvtHEMnXb+6C62XEGipQXojqyphHdyv/5uWc/Nyj
CHatLxpzOafVOb/qAnZIs8VyA7ews84oIhn8wM3OB2gHRTOrbqOWflwyAh2yDhac
P6Xt+6Zt0ivK3f/4LsEOgJPXLF7FXGi/tKr4s76AjZ/LyYlU88utGSrVeTYnvo2C
jo/btRWvKoT8gtgD79GPtuu92/T9JuSFcZ7Pyt+2Mw5xo0r6sUWNycRwrdnLZJRq
+7oxhBf0z4W2yJwTCjizsPTGN/C0PEt1Ww5Ok2+ZB2VP+2c22Jh3CyQtWd2nZRyX
/Trqx5gEEpgKV+9szgd5M9clEPwjNq9xV0eIEmbYxK6MCmbnOfc/So4J7MgUdiYq
SrAn9mRLF34zLn7isETTPF0ekWWEWto+LPhcmdetUuLlmEPi3IguGAXHl2jIKP44
9L49pdEbUhZsXju7V8m9kdLZLTLkSyXWks+Iv+oS8gx4o4ImnwjyV2PT/gGzPdcO
CH7isC1YVHOjOHV7Zk8RatNqBNAXy9+ROUSwAnEyDRZK1zRIckT6nJcrmKXatLzv
0vjpyAuB5Dgf7YmlXW+vWz13tzBZcfoI0r6FcZiQ/eWFmZEtRDwQkEGJb6nERaXF
HhNFTROgLP99NJo8imfvUkr9x8jkbRpQCbSX3+lDtVWgEPS5hK5sMdH3lvvTmBA/
8vJnG0PbfszyvnFhFeOm3UDbaeClgSYQXox+yC5T1IZCWEkwGxCxmVLd/SfMgjeF
czhkYDAldcHRtcX/TfX/imWZgD03nfU7LX4ddtRJcUSxAUxKow43+vYcwBmiKVpF
VHvU3Iey6K+PAoAhTCy+2EOnCFAtZ6TvzVdcMh7kYipuTebLUW3KufLBoED+f8/x
+V1AgmCErNy/M0ORK+/Lo3aaeKtQpT96goimglQxafZgdUkmAMlypJbHAMqoouMV
9Q/7NbgpySBYlO/E/GREFXnSsrTLLD3uFNeyfPkm2q96dY0s0YggyaKwyMMGopKN
0LInJ4De0jJusIH3beWKUQZm4POW+UOGbhrg/CUrg31V1bBhnaOV61bxHxpDGjEO
8lsk4b2Gvyrgz2Qb7cB5aiS9Xmov8wVh2tg5LiUJD7vnIdGGJdBfuHn/8hKdsYqi
v3DetXKbmR+MZ7IPqKML/B7DAfNVSKzXEdfMGhPGfTJlOmrhnz8WD+9qa/aRwzaP
kQEjBLHfytbr8pzSKyBoTq1Ie7elYWB6YnuD2NdKgT+AxjSzoS2jx0CuN/Unxhim
2aOxxdFyQ8OiOt4d8lcgF5YfzKyTnPXKXdncxc0uUN/CE/6VWSWg0gfzF/Zh5b5d
q/Mtei0ANLwJL4vAwqj35meug2gEXlfaGB20jmgGWwR9uCgYMXQG2c20BKwEXlEm
h4BZd7z98PAwtBaUie11dtqDuBqlQQiPsrR+kdfBKBcIbeYzYpUHF5hEr7T2QrBm
7PTWxhGT85MJ+g7845zqsXZVoYbobgh6r5BcgX2ffH8nNLTPMtv5wWsbBS0hhcU8
VAT9QjdY1tJNvr4M8XbUBPMk2C1emrKvAqk8uuDaxzF2e5iVh9312REHztO129P1
+KfeB1FksYH0pEOk2ULkHVNOCDUDx8sFcN2v9qtGD60AR4bcluMLKHo9a6VbbWwY
xrVtBOG61Um8hBDHSuUTs2E9lXQ+Ank6Eo2KTG3gcuOUa3J4R47uLfCAChhsi18o
4a8PW6IxGHTKZnmkzuLd5CEGfvNO9vHnNtQ3nDFivgVpG1jjKduP/ASZTpKdwjKy
OOxajnjXj4zHq1Sob1Q10dwlMwXi0jOG3UnJnZeC/mKJ/a2wWObXJVTSYJSkc3bP
oSkIJorHNpJrfFZm5A3R0IS3sBTC2fxDSsc8aHEh8az3NYFbmpxFU0IeVOuQ5Gjf
zvPqZCkMCluR/Y31OoWZm6KIm1q3lXLUn/akzhsBQzhX+4Hf2yGfYzjxB4e1SJUG
2BXqplPoygC/5hnwnFdzs1smXiYePaCESZt8d8UD+2F8HGb7ieP7xMEQoLwuJxfd
O9tjnrGKIskjEd8CS8BN1+Buh0tDGq94yp6LWYzgEvDHX5jQ3/tcEFei2kze99ci
ydkefFqtfhQ/twAauMFpenP1evdzKkv+I0+iM4pYgvempkXIE/tWowI8GQF4kV/H
ctEsfjzZqMb/VwCAN8CAosbWrD1H2guSP6NuDig6Y48J1rS1/mA28EYE9U4F6y9p
O14z2F1g9giFblfxYtHGG5gP+0YzflhUrVoY78mJr6Iw5fOgtt8FzijnyS60g5dr
ANBq+4gVBr/jCv1QIXmsVKfz4Si8MHc1tdxGkTFE7G69X9hMy28Dd5j+K4ClGLmY
fSdTuSFbCNHjHmGMFYPmH46a2WXAeUhE5mFXYwFP3ORl9HBPgrIA1SE7TBeT3Skv
Gr223Y3hUA1DnF8M7BKO1m6gVm1sMz7FrIjxk8Ep7IQjNLjEFk2spj5ziWPwFU80
ZOYUmorMp79BakCFnTGBL3wGYgsn2O+s6Yw6vnHwH1cBndxx1QoPiU1Rj/z8b6Rf
6x22F1H4iAwwp3DpKIMmAafYtczO3EZBg0fD1sapwYYLU3Qz0PTqKp8BWaLaA3m6
aude9IH3SwPGHthQFPOGxYoJj+Rlja0RO+6niSMaxOQ0G0LtKakOlok8vZqUHVNi
miWE/aqdpzA/9hU/C3Scje3VED+GRGDHcCdZADDO972D3fsmInr75n0KEd79OSM1
kQUCMbpxu3CKbs7QMQ052cYxyRgbBfLd8bmR0EdjyqW4F4LdMECDwESxaaauajmg
tMgGJ1p24RY7cQdc24q+Vv9PyOayS+LEEOpjA2G99MZhl6fF/y7eXHl45MQ/Qekz
G+2SVseZo0+KTbnJ3G4gp9DE6v3Kbkb2LVdqPRQDq551PHmNBF8NmaYq/nNfw826
KqCwyhiz+1aLB11Zs/j/Abv/SiQN+rXgNywANO7XQgq7yZ0la2/K3a+XIZtWIOvK
N3flq1xKIoST5opZgxMXfWwn6pEXFruKAzFZAqBhofGfbmjo4Qjw4QqJBxj4ObYr
cAdZqTMzLkDhomWkyKjJlgYgOsyTSXyqNX+eNa/YDALk+zfVAwSc55wg4mm/t85r
49+gEbdMf5EgEgGUDEOER+MaZL8hnVZSDcIgOTB9fUy1562lu06CliAZKcJZ2BVl
icyceEdwr4JvLAcCrGza3xRGcSl59KiIfXtcEsgn3a4TKiYsvF4oQ6lBQxyEoZoE
mdWmdWwv8dPUgxEg+R3/IYcI8CJbMgud1ddFveB6tiBsV/adh77uMXF6+zHZAWb2
ia4e6jwnuJMtg1O7hCmEIeAZMrik+gtlRj+poTY76eolY8YNo5zOa03Ge+TaG1oQ
0dYupSfQkuLHeURLgosuSE9i1cN/wd9jf5AA5TAMt1O5x4LVWlUWYZt0mUONlSjw
UPtvFORZWbgcnt5vTdK5mLwgoAFHWAqmiGBXW3EcIke0d6h+Q105/KlP/Mt3AOxM
aUE22ntJ1My2dk4nzwI+H6KU112in2kVG2JuDqpmwJSdpdV7lR6iumkJ7BoizGxA
eG8O3xg5CmoPUTh3jabmK3uc2ic111ZDkdWmsl0cBshAjQa8+7b//rwdiL9al+yC
PgfYzptOA2VmlclicEWRWJe3MDp3b3+Ov3cBS44NBOgstdKiMzgHPwIul5DnLFO4
7fl5PUwC/0PDGzw9m5xXc008l+bdRAjoAGWaP6D0p2WjpBNGAyVSOyfEKNKiYabT
AmJWMRBd1DR7xqY4FGJRuwU5Ts80fau1ePqWJ3/+AHKNERQkVDjZlDV2GUnxF1In
CODmxxJJ8dP4o40Vu+hdlsjR5w8dwL0WYuqh4/nonBpQRfeBvVyjLYwVHhg8hJcd
KS5nGnE7/vneuAuHd5ITFZNMalHKz2XURiKqvMGMpu3KbOjJlmR+I9DnGRSelWz2
zoUqiBeRCmwsk/GdU/j3qhCPNL2c4SXO3optXj8BO22rBM6bSwr0ZmdZeFj2EpHB
3jlw1n9HMshKY7DfLjK38QBGmiVYEyGsAIinmUHZlBBLmzWUbZiMOzTtcUsv0ktT
4rvslcle2Vj7X7kI9evqDgPIKirF6+yRYS0FsHrdX8YXBczi1ZT4Z5TdYGwe+4oz
35//tk17gUNakw+H1PKjtkwAthoBmj4xafeYKa9hIY9JILMY5yP77WywhYhP2oW3
NSsRtKFLaxkuDycsg0492u2GSZVWmaxSzW0W5yQeC3gJ2YCM3Ihz22iUnypmzpkT
/WYAvFQm9h5RH77dWlqBnpShWEKmJarmUjjcIJz1kieZK8zmWhMUmV/cH269eapG
smhNr9GVSDTc2W9FUXoDZwyaGJXBu4iko7OAnhFQ0+KX+NOqdGbka39GnRUQ3Bgu
t67LBlD6moTeninYB2zJllQzzNNo3GfxYDHCnvHcFV4q8RJ9vswCAbtq528qFCrA
14t7MyZgbd+7EeJsrgsPw92SEa1s7q7RkhJVbxV6uOPJMm6hbV0fQspQ9g/AbEBs
yYHX5ihQaCUgWQwnyBPkXg3mDyRX4kxvnLLpfS+3u4ZQQHEB62RghsjnmU207vdt
NdF9RH4SNA3jMhU6cVWAc9Rc6VCZ8nBP38R9HMiiDCZ57fEPonLVioxBqlpE7+F5
z1qiFby97YIvY55Jb+5AMYBfYbEsAGr3kXMm/VfuDhis/n+NeOdXoYTXPYwKYSjI
1jnb3RRrPf32StOpQu3iw5XqXbmMtjnged4G9dlqoubQJocS0eyVHAjfbtDYAgGt
bh+vnfvKAdKNVhYHzQFJp3Z2I6rNvS3y2PZOCDkj9ZLZ/rFtp33bDX8tXzvoIpEW
8RskIYUf108QjxHCdqaZSXNiMZgfE0VMo5rUop8arsSka7O7BIUccOvQFit5k6AX
Pf4seFK5hLjHsU5MUgCHkI2WDVfeSqoO4IujecnjmtFYpyeDMkebhb/lQT4n0W/X
lDn9HjRO8jHKBC3E1UzZ2wTcQzNUn1HJL4JJ17LfD3gs1z7F/u27TuJTSYMZC7MZ
+LSo0NzaIv5oup/Xw0ySk2A4+6Mu/030ot6bbnbJ+hwaD4a3XaFxMJBfwzD00GG1
bgSwDZ7Cw/X0yiBUSVYvMJUiSIv92+c4dBe60kPWywBoMPUYqIS5On+7dr9DNrAG
Do/Gm7tePuWVLN+x4bYGzvkMDJaNsi6wuFDCXZScDplmDzCD/rm+PRTdzQnZs1PH
KRp1bQT8+DbZcKu9kCoiBk5CpIWhixYt6urRtRFOOk5vAi+X2Vy7YIGK8ExE9F9+
74tnf4xHYHIopCdIlnviEWXQc/anSoYy0rvilN62Fh7I037mdpLdUds4bT6zP/0K
yTIX6F9bi9ss0EU2NpmeEoNoMVzpmpLOBBJHz9Gl/cQSNGLUKvJ+OzjkqLHl2LxK
GnMVrHPIX/+DjPPrr9FItAlhtd7rU2b+FOwnA0awfXMx5q9JCULcGyNDrMPQ+WmI
WdqC5ztRdASG7Iz+95VPYgI3GsopAMQLEDDZDIz/f3rDwOY56jqKYIUC46LndGa+
mVjAOGNnXRWchuwnBBakyysmcA9+3eL6ooWeFeP+0xMuxZNLy2T6YWelBPTgZoxb
4LbixGnoPCZCVtFNzkayofTfQ8DEScrdTIJDjxfbyJd5pOp+4ddTxdMEDIGNwwKT
8s0uyzW2OHa421XCBxxMxBOa6996x5uQmCNrYFPu9Urpbr8FLhCnVrLdCnqsF6Uz
4ppVCGH3DN5UA3plG86u4Ru3837JvtYgyRzwQomV8zwQT6G5PdBMEvlMIhEZ50/z
ZNRxPxFaDViMWD9nz7o5R2X6D8BE8RpoA8CZh54HXl8DMAnLEl0W5v3gAOXrRd6u
ySUqVopMgWH6lC9EoBbDpq09rbemtjzZaJLFpWizykjvDgA9TTuPWvIIGhcD62Nx
+vm30+Yxwguhm/o80FqP5hcAGsetvRwPC/ZGKEEI/X4YhBRWWoqopYTObrUdLpKq
VEKbw6IguQ1thwa6fjAKIU9N6YKnrcaLr/KA4cxb7JAwGT7uS8PLLyZ33kJCZTlf
WDxl23kBjxAKsULnxHEDj8tgYtIWlKPuCwyLh683rYCWuwqEU86RQZFA3vSXo6SN
B4PC0S9kVnItWvHASM6NWynnJZIsyYaA7KZn1TfXrscEkCvpqzHPsp/KIicql4mo
pLOvnK5hQEmWniNCB67v0Y5kNOcILUTzy36NnCZxVkuJyIDXvKQEelVWiPulA56l
dDKWMruZRNMJzipAVC0AmhfCGwBUPRrhL2EUUpRQX9cYP4IWanU4plRFnXSS98YW
gwSu0LCMk2n5sRoHUeMnindI6quoLNrsAyf6+VjqA/ipd9mRHHqd/M9bmm6KBE9l
RRlJ+1JI7lOPygMz3RivQf60piJ8dzvh53q8VXN3ODAjs1arYCYXbmg6SgI+dlQi
6jmxRaTX1BfSV+fCxp6zFPlndOd+GJ/E4OIpQa5HDhj6wmiwGjBa6+BqD/0j69Tp
zId2WrfVLIpbtIi87SwsITTkfj/zUmJLDYn9Al+XsLgLE3EkpjY8lLhXKISdRpGf
pEJLBCNYWKrGKnH1UikgXReWrQ0FAegTaorHB9f8Ir0TJLZq8MPifbglkwMAmzcQ
qrIZlwQ2dlj0VXegMT4+MK3q7wia6csZ+yjZp2suKFIuL3LAJ21qYBBaXJ+6SwPS
ZXioYos8c+L6EwL4goa1PB0V6Fme4Z3hj49yZg7EL+DFYG4z+4f3oJ4cwDYZpo2d
DsJrShhYZJp7uxVe6v63tMu8IWutSgROdh0Si9KHPa8DCuA11SsKNu9OuFETDIj1
JVw0cdNLoLr3vNfnixe3++zBZT3hHhEUiu5QTc6tmzHcyAodqZrgv0687FXhMJKg
0a8Ek99meLmXxB79MCHU7OjN/g6JbruZkTnt/98x4gIKke74kKlMkmxYB+RrSa+c
0RNCXVH9p7QsxG1kgRwvNuWT53l6xUh/yH/wC8BzPysqREX1MatqqbUVVe5c3g7L
RqSM0Uef1jj7zFu2R2W3t4/66Hc+tyLsrXq4NYJhXP0sUxENJ1Y8JI2yMN2EWRZn
cxglVv8mfCniglnl7VTtDUYljiF8qtdH69gpEbmZUiLvZ7t2E8htdODbudTy8Cto
r40pCW6vvRhAwz2T/LS35zXcC2yVS8OH0nlIPkOzXAUn4Xb/F7jDUK0ViJc5AE+i
cjYUu14va2EIO+k5+qY8KBw1r9w6Tv3CpA8yevzGR5fxOsBtmUyI31xuDyvNknMc
9ah7dR6IWbFWd848AOjh45YVZt7zerVz9Snb3B0NVeoQnqZXo6tmnsimYMhZaagN
vUaPlh1ym0ZOUzGM9tpLYJod2WGuUAhbm4VtOpoPZ4vQINKZHBEa4dSZp6e1JYVT
+kB4Ol6/ZnoJwZYebLN/jpyqmH/HXvuYIU6is6WerYmBgNCWcH+bljXBXBVxFt9d
wsQPb0uTccfYTw/HZ05JK8TBS20asCJja+6JfE43JPlVOBYtlDDvgCm3vSxOi5Mw
yR8oWgZAccnguvSj2aNZ1ob36Dfr7wSWCA8YDLleMWtJCb6l+aCmrEmiqdLGoHx1
1kXcfFXDbyHuBo88y6lwN/+Z8FaTm862NE6FVYGmxt+YJSXA1BCDjyC+VTcmvaW1
6Cwii1m3CwrdXhIIBzFY8VR5D030Yk1RB31wjiuinC6d7O/y0LfIYRBSnG+cLTqK
3C5JGYeTcF4G2emBZSF4R9H3Ht16DqO4nszBZQWc192MLmiDjlflYbGbzSXIuje9
CJR7cGRICukvepiWlJ2yBc9HdFtK87WuWGH6m9cEIbGmcWf+PKwGLHe6fVsNz8IT
CivzZ2040eAWO8sbZ2UEeYM+017hFpKz0w1RlvK77zzbddfcdJlmpgVtPzAaaz7o
WYiHdX6QpDDdqL6ElGcVunycQdzPCx/SkEASH2X6tUMVzVxX0BNDT7f6fyWHDeg2
uwc6B0+rny2MVTW7qm1UzuGXvG5IMbnfjaxpH6cycixrzto4yOlO6n9AYVpDVhLD
AovUQc+0a10Xam0avCuuUpcHuS6yhVwhTdewi0dPgYBTam78n3eYAtLuqhFS/a8s
72wi7j/HB+DPCHsKqedV30HzRbiFo3LwR1BKsoUVwi41uSVJM4JryQrjK0W/yoeX
JdS262W84ju5FAnaC/IeUMkh2kbRNFzsrpVE42M6p7l7tnrKshFTLa5+N69kzQZj
j7uRW/UleE8Kadj5rWf5gQc+V5QSl6ujDoMgSLnskhFOrncLelNd5g1dRrX+++2L
b+zL46pXMOaID9+58Oa62DKcgt7OO6gSX+QjJo44xPtIup5aKJ0w/S30aQFQZes4
dKBkmIyCmXNHi40R07ajYCwRFXiO9u3LBzHnLEvt1vJiDNx9bQqy+k9FaGE9CKXT
eMKEi0kHlc1CfA0uBss7CWS6O4tTMJ9PAjFyjkS2G+BmLk1xoKw8OL+mpv+bM4Yg
Pmuq4lcSo0thXzkfZzePIZFjKqwIYUBY4l+AU2+ybmdNDyxcq7tq4rURmRIoaXoo
whbJxTtZQH2SV7r5S31JSfHV8bIHEEF5yFVTFajEg5wYUoSSsEV57uXrYeUUl+60
E/kM8TAM0RZyDs6uhEsg1L0KxHulX29QNR7MMvD8w3AHZr9/biC/H6k+mh8/JpN5
ZsjraQXXCiP3en5hsGQ/k4gKvuKMHotW0iUhwBccGtQh7eG3VCvB8kCuWeMf+0Gh
wEr66xYt7lbWhx9ZhgbOrfAroX9JypnYETaCbhmlbSbd9VBWapwTdayh2WuCic9r
pBTqn8NibOO+6/fvI9Vhc1JY8Yd7JFeH2ulKtIBZANL4M7WuSk6auhvwfKtrQBaN
hHUMpxzoexF67r4zAcmAPY4WdSgOwk1XHFNy/tsw8TmO9c4xqjrbcM6So6g5h5Lj
5Ot4GauZcoxBbjQfSfUANc8Vvhi4AwB+wKmL89ID6v84FzfdKD20qDFiS9ncYWUG
d/2jqDYCRDjaDWqURUYRqtoqrrvzRGlDdooOY+UkGvs2uJgaob3/B2RGLi3OxlH7
KBOq0uRB+VaNoLSAZ7hRCD455Eqy6/QArG9bO7irprH0F1Y4ny4IgYp1DJMAuJHW
TkJYI21vpKKlk0qlugxhsrC0rqGHZ8NitXhq8ZBVbe3iwDJrTB+zP1+KWKYKvgHa
6t2UVij8JFrjwbToDdx6Ri6JRBdHL2yo2S+8lYjiUs2Q+UeoAGJmDEbCinE/8BEU
Kco+PsJKIlhodqtPU0S+LNxO1TiRH7VBQS3MXIjrxuI3VCzTscaGKwyL72g+6+Mo
Gve61iRbIVAbqRAuo6mo7GqMqfRGyrGsrb3PDqpRCSWoCuvXBeMRW7DQ0GPz3U0q
CtyzWdXzRFdCO9l2JGlkHI+Tt9mcFj8noDN9qSZuXJA/mDiDrqJdFWHm01NuaSVU
zB+78OXxLK01Go8sKOIq0UeJuncPPqmKCxTcYwASuAO7CuBiusP68ZcK5zFm5d4g
X1tCUD3mrX1e2AnecfXX1dKaOcYXyYS7KnpDcX6bQnoy3ZLYVOfTHgW/YdLME/eD
oncRIH87gzg7L5nATMctIdtY34NJCmq9vId3ZuMUMAzf8oO/ry2AuQcaNJRUDtKI
iHQOWVP5fhCdPyjXjhIowyxhn/bDVAmsI6owSilVHl0gqzym4oZI2i6ZtLIvkBfn
pWOwIKQ7J4XzMb/u1Oq8sWi95t3zfctjpChVq/mseKGkbowqjFw+EkmLQbqowQ2f
Ya+E+VuAGw1D/TcGVsSiUWbKiB9iuHMgtOj0uJ65+TVoY1NZnBgR9JYdhpARn0A3
xFXr4+KI9ruDwB/zzq1OCnyoEKuHYVibos4QAbqGlzyTdDy11zjeUlwXB1KRReyy
i1Qdy404uZE2vwk2eIaxBANUefpx2k4SQ9Ve8V77G4jxx88LoDQrOXjNvJSI64+5
Ebl4XZTmHw7LzuSejA9/pKSlGhQkiydSFdcbBoRXiw8ahNCkkaNVeSwDFBh84YxO
tRv9Gjy55hUtYa5PAe25kxqbOkZ4TMZJ5TLh5jxCCb763Na9NJYT71IdhsrdiXc1
UZnFF1AmSlldxRv0HqU/j0qkk/LGr5+aDwweWXw8fPNA31rgKUf4eweP3z/TmMVL
sj2jLcm8sDCZyEt1AHQ94TlglAGV0E2Cgev8vrMwVQ28dniv7xeoLc+DZbMv6Wg7
LzETaobRYu5V7q4p59Wv4T+WMgLN8V3thkvIWu2kcTlGMVtJwwPrmcaZuV/XyTRh
7KVJQJPpfixDQ9+OflayZs6PGjpHi3QGo9FCC0GnugDh5ceHFbyuxrTKiFYtE1lF
5KrDXDT+/xMOppA2ux5Ix+gcQtRuvOgBXcAIHSY/KwQiG0qd2ccwSzkuKjuQC03+
kJqJfe9CZZsqBW69H2CGG7Z+oX1SMymzAUSIhSNueOGSJRz2L9pqcjK3ZzW/lSWJ
1YVGTHJd1Epj8cgr2apkD0XCOzZB0z22g7qnhHmoGdWNHLcEjxZpDXvLpXxCG9w1
kJDdDDlnAzdvh3Hf4kjR5CKopXqSlMNdvlFeSAYNSH50r7fE/+zNZeskaRCwpt0Z
e+2E0O4fSOvrOVpKmuQs/lZGtkrktzR4AtZXs+Jq4p/XM2/ovlWbDFlpY6+p/ekh
Mjg5zighEO/Wm9gSW0TGaW3RJSOXdiWRuYchEWhht5u5X8g6DIJfuXyCz6z1WW3h
5ZIodS+y5LjFWh5MISKkk5rQJGESRnCjXSGWHZ0oxV8chQE+S8QL4y6hQPvZ5KZR
ffTjA/8zO2Dmoj68Ofey3bzP3xXUL5zXApQ1WoMRBvbRQOwceFbL+8sAZIr+DCAd
pc15230ql1vfzgm345csDNyMDHm237f4UpWXX3EogaKLvSbB4n/VUEQXbqmie0Td
RhX0GnPlalzNJoW21fiwCoKRqviSPHZ0/BZ82wqwVWEjHnhDyIFNX/hPvwb5fW3R
fHXX1MmdYvJfRmV62Ep2BAKUfPxhhrjDnOwVIr6v2NWUD5hJFRj676daOJXNwt9s
xBZmcMjSJvhblB1QrhVlDXC1gshHuOk2SsA/H/RlqJO24Vigm8F1SRUiQUGBYiFd
1z0OOkt9lvePnJ3ERPXUamNkLOAMHkhIj2gnkXD9/gVpzPSvZE96ArrAYVoe1MsW
IWGscmT0PZEfJaVnYw51OmHwWpYCLkCRY7j/AuhfhwCS+aYNWUOd6Sa2SP1CJ6yh
szAHO6xFd31QryW98f/0iT4OSQT562luxTwrdvW9CZbqMkUKLkOuf/aUCy0kaIv8
l0lFVxmgxWY5z6A+0aK4Amfrkgjeu0CvaCClCz54FExB78EXzMav9yjZfJeXBI+3
ebDaj+W2ZWgouhb0mfVI5EgnrxI+cJN2WNkJbKTj0oO1zFg7UgeyxoAJVaBUIYV/
zfh8lDjPk583erSVNYC8ZKV+LYOl/kCZDtMWwu0sNX8OditIrjFXk7Q1PSYjEpUU
TVUaQlziKHxDxFYB2q0pISSKCLWzIa4VlkVfmBdsBV6jobXbNZd/4h3gK+MVvXRP
WZ1bbFIN6R7a2UvKVBIuA0rSTcH6xgBfCPR4azha5m3VI4ZfrPzHAKGx0czjvqSo
RiX6jeZcPQcOdItIuTfXDsLZj4MwlS576NjqhJQsvkJ1sinDFbdzS44m+N8gfAQN
RzGTQZWSM+Zota1r1Kynex+BUCsd8RL2iV0Gyw8ELM8dlS6MlyjkPR9wvEGjFDSr
woNj8j+8dtkfmy7iRN3JQhRaJlK2/ifmhw1tkLsgMjCnYKSXJgu/xhEMkesFgeUy
odg0Pk5DTBQsd9aVPi5+AdZxiU8PsQEfkRsUG7Mc4i6D9VenmCCDkt5rnsIIFj+w
Fk88y7qa2PGdApb0EZvSPnsHIjQTbTVUfmINPOLOWHdQigXKgQ3pVlDl7XQv3BA+
/rk4ci6Q/VNKpCDGmj42KO7mjxVQIeF6Hm4tO1YrezORVxHIW8fNkUMU/eOJtSNW
VeUdNT4x2wos+R2/YDB8OteDvn84hgg/WPCvyT9zwYXEP0hsphuP9ltIXWFt2poQ
HOoY1wXGbWTeSIR9Pxv/Th3AZp+O2rOEQ3SNAsWNaUXVj43aFPX9EukS9R+mxbdz
4Fl4Solglbn7HUM9Hn6ICPHJXsAB+skzFPBHgofwlcFZRTW9aCoXEsQ2PUWkYYMD
o62iXsNe6lSqSBbVSfsGRKRoi59l+9MXLE94ItRifUhgDFWfMa4VAuM5sejka3yK
6VR5KLYAdCvIEpIlNYdgqIqa/8TuwieBqmY5btXiHu4r/7/bBCsZAatXBIk8GV8v
7Mxu53U6PRWQ+DeC5Z4+q9vdyCAwOJX60ActnPh6pKJT0RTWKtc1Uc9bBbOqyl7+
HmEt+gXoqPikZepyIH7i1oXvTWbTZ+AO+l+JV1RNfDH33wqKcqbbksLHFbxmj81A
MJRv5oRQAZu0bm7/DtVP6Eo+XnovFx7Qb0Pmt9cxysAoWARGh+cHHhCqExW9TYgX
GoBclOYb7NPmPcndw+WlyNHBXNbvie+78TYIiuoL5uNC2Mm3O+xfy+vg+dwPFFSQ
3Vh/JEh9Ih/oeOpT3rnwTlsr12zOKZs7eLBtxBUkD2vWiZXkhE4MVmCcZ4Cozs/O
xsZodYqSDWl7LG+einMjxwUaRhiFXKTNETYIG0x9TXdWTB5VdFBu1/nAsYXZqiVj
Ou6ytfcpabwlNrSgPcQuseK9YHpcfJ8XFKob0Y4PMMJJ+IQ4iQ+rIMZyA9GjIAW+
qK0hTniuVego2az9fUyxDqE8mFVouBg3G9Qs4RrFBPaTILmpq4IB4IwddWJekRrU
rnOBYfPEDMMhh2YlkdZ6la5M5Y0l5D4xcAg5HMKyUOIBLGoKG+PIuo8yS8yVSj8I
YcXtKiKViYsrYt9wJEqTBblEdyF4ULRkhsnU8iEtTpS0FqHUtlPIAO5S8DwSsiGU
pCtrKsD1GWl27BnvatZzQdA0miOBLrPJwSXu8X+Jydhz3q6YiXgxG4O+cKl1eVhz
2lPIGYbGo86X+8GeCWemdN4IZ5OEc9AXtKMsFZIztMqMIfc+8v5gi7GZjjxpBjS0
xWxHITGcUc4pf1bRYZJQVxbcNa0c88CsvRRJj+LMQu4hf7Mt18/HWU6AeBD4k5wE
34HW+LwDwa0xQROHfkmqConccTfis+p65tusXqEtm+mZGIps9I2YKRRvcHTCaA1W
7TGXp6KIqTKRSSdxVLHKDAX/vWJAcczKudixjSo08p/Y7pWrmMctQlIyU/mNRLqB
HbtAY/nq3NohquZ7i0hEF7W8t65MES+OQ3lVBnVd7sgv4SjPTpmOOOYxNywHq6Sc
LcdwWZ0bFckmlUnB5u6FQS59aVVUJqsoBBLXxQSQCyZ8uzi04BsxeqGwKbyMdxfW
HajsG6wgoO72YsCr/LohYLK3kP9R4TOZPjDGVfDg01jz3SnzoBVoLkPObFdMhrJY
X+PeZQ9iYMyMfho3OJpsnqlqpN7oxG5rq8IyCrwFIeAt7QDjpzVM89fky0o7BHtK
KqvzLWUxWLnmrWmpEL1dFKflO1VPj1M/Xp9dIl3QM6c8D4L2iUOr8HgD29yQHFbn
NIpN10TEjOTC/nCjRAPfZe0uUdo2OFE7TztAijSmL0IWYZoGSebbjzBg674tasUg
D44dszJE/1LdeCsixIsTIE0n3cuyYVgOrL7b7FCaSrQlYLCv7xr4UAaDn4q/fGLD
eFAqwZ9r2VLRbMiA6wPf7iYzJc2eEq9xVz92ATEq7blXmUcREczHU7C/wm54MbSq
Bb2yHTg+ddMwlf3OWLT7XEmKie8dGOxeLxIFYT1mSX8zOMCjdT5rT6y1HcQcyhma
FKEcp1kDcYVjbd3wYNciZ+eFVw5bh/8fZn8raloR728f4bzu7NWvgGWTo7ucZW4k
zHZBz1WcD2LupDQ6gfg09GxYBtpXdll61D0ZjByYAlHoSb9QfqIBqwyvC/GTwK20
PFw4BhrgcbinEdHZg4Qgrji6o8VJgXQiszy2jUWRjSPT6T7WhDoqMmM6M6JdG3RK
NrdB4QMbJvLgsDnJozx8C+uN5Gi+CoyBIp1MlQ3793JOwKlEtqo8VPbf5JnCimXg
dQ7E6DSWSc0m6P2f6lOqUI3zFbNIYSW0v85/+0G6PRrh7ZBYS5/5k72yaR+yujB+
`protect end_protected