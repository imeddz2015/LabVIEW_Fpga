`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 12400 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/59UwEX+aE7FohaWu0/8IpTj7mav863zUNIsgIH2BWb
Abd9opeuBjbGF/waQMI2vMJTwD1ie1YueHc3nSNpEh4OXp8P5ybZFY89uyGz3ztU
W1EsuUnchJoQgbHZ/sLbgtGRgsrAFn+ZoIeGN1d6RAF2wAESJmYP8zw+p00RvjZ5
G2ATm2jrAjm+J6bPpiDE3+5ef4YRS0a0vxKZXEx1MJvxc5FryocM+YAf5b05O79o
Rhb+/a2iD12CMKG2AvGJillXWCQQ2qHmq/KSUeEF+2J3k0W8q5tvF1djQFY97b54
E39OB5c58mZEHBVSWY/qphfV1gqGvpDwGt3hJ1tkb3d6KfNda/MSCRqPGkGblQZZ
C587/afzvWr1Nmu1AfJQS0x4Dg5XqTdNNgiIaqpISbFOwrzBb7rxmdbF6h9fpA1U
a++2uAfqRX3LNVZ/rkU8l3u+vw9kszB2UtrT7Uwic6wvb908j35v6kFlLLGl+54z
eeoB5euh2+Fa8KgpNFD08hCDuVJF+5gBHsR4CR7Q1bLfpXBGvl8bMgjGGcSVo7XE
Ck+6+uFvFLDjrFqpdWVYOIue7ZtgTxU9lP/cZ/qSoR0RTblfthfvQxOtOoNzKrkP
xihyghS4f91WfzAhXOe4F1YsKSWLWkfnYJSPSA8Sh/gE9j1/78g08EMUZT+nZUgP
mFHwlogmw/TYFWiYWwrT1j5BeZE/iuz+Aq+jRm1nBV2e7cYwDw4XtswEnl8ePISW
bA9ho7612w3FTX3fUpV1JePCDZ160mux4hjAvR0HM0QsH3Xnn/TQAS7qJEv/dbY3
K5YzWaMJJgTTjQpyTOYGAFRJ6DZ/W4jKtgAD+sO967t2RMkaM+AzZyc2IXgYcdIW
YMEbNi5qzhNTnL6+S6ianQ2Ou3LW/3H/1AlXm4O6Sfxn5c5iqdlWq05jAcbNtddi
IfcpBXABscjU6rc7+96RZDQmKHF9QvB31CaQcVakaMfyuy/IeN4e40V5KRkKRjHr
LWeM0c+bV97WPtCfu+AlpVDMjy9bfD4iVj7aemsTvQG2iQ3NGqVmMRxLS/OSdP0L
A4OhgO3QqL/uTh8Gxc/KkBIT02yfC9Mm9AXK+PSJ2SO8jD0g2XKPJDL/A8I07zUo
qT82g811Vnz0XaW+xNsUMA4oNEk4n3QFz3buoJlk++QG28mTv4Ft+EkYdtvQXtOY
OQHwChrk//QIJ/5oA+C2/nv1FlYX4dfJW8t1ywHe9/bMElbYJDIdYt40l7kSDHAm
m6O/GJ7yXRAyC3SVGSrA/3ER/2zkNYg5qFX6e/ay+clc03h3iUxrvjB3HUrJoP0X
mpS2pQMDSah9S53KSLxV/unjgtpeis+vbtpqbUZ25DeKKV1BeVsytQ0wF9vDbgVY
7yM7+vuKC1CZkHEF4hSGpsyaLVaZNXXz3S7etmBgaJa0ijcwKiGQZN+rIaxHgPoF
e1mWIm7tdAyB9TIUjh6f7H1s0dBMbqrWwPJSeLEnapyOcyqN+vc681mLg/7l9g6x
asFxJs/oMI8nec6WGDV7UvipQDUWF6nbdbZTjcTPe/t6OET8YSXh7VrJ4Ztoidsa
y5Sx/5XiDftce/Xzff4fP7mnlyRIgd+9oAJOn0CPQH2AZTmN/5isYpExEOsTxpji
4GtLvX14K4OqlD1UTltMIdxDlcvLts8emzUGtcGqGrWz5Scbkn2jgIc1VQ1ZDubD
3z+Yr4qvkfLBDxs2n9+4ZQfrXXseD8PS43j6fi4zK08e4qXKzZM+lk9t9FKGZpzm
ecys0NhJ/jb1iadp1ZvbGc7eo6Zypk1g0sAKHAOdcyC9dAqngWkfWTweMqYk5fVV
UCqAs6/rROg34Q8TiRwNRkxK3UYPrspBCznuVrY4QeWqaKszazjsbiAnVe+pQvpJ
umvri8LOnC2vHLdrt2Odunu3X7QtmvhFlVpowkNjdIrxcvxemHYmh1y+TgIsITgx
014F2gG87EDZY4klN0IGSkSEMS6sxKWF5sbwELoTHFuZFKPawX0VqUzhKbhEyyyg
zlZ13wSCZZZoA6YwCiQRKwE4sOROa+NHB2QarZZH8915C4ZCQ0UH69rPR0DJ1uKH
VOQ7YnAjv1YIzm7+52Kl9nvH1sjgoLIe+RtTAgAhZMC5bqPBH4011yRo5GAKoad9
MDfsr4qiwTHTyvJfUKDeoVEcE5vQSrmKYwjmY76cwebB+9oWZhrZULUI9ZXunG4e
goAnuvuTTyVQNxgtKKHzCZ55ttcb6njO+WQ+d0su+QlTUXIW+DiH3HMPP4Q2SA3X
5/A8OagtcYUBdvymYJGnXC0CiLrKbo62yXudDZK73+k/kloefX+hj3Nsih1yqkkE
NFK74tEqDrGlm33pO0fCdDJ3BGUMz6G29Enw7jn1Ru2TMeAozgutD3dQ9V//MFQn
KTdeFQUu1qBbRDYb42TRUBPzBR+hPmcLAtDw3aT7ygOhs+eDFSOCzI0RQjij4Bcg
tH4a3swRpNCgQUCQulvktNiK0muS3iFiE5GZquMbbvQw2TMjAMdvd2Z+QgeodC4U
3PNeCqYFoVL3T7GUKKrezLw60rNEvNh1M0b8pKYO9UwfG/2XfnzGZmVX09zita5q
BSIK1nf64sq8a9+7Q7HOQYriPDgR6T8fLxeEYTuN+dmSmMsBfJ8ua3FyE7TdraqJ
x3H50EoneQgPdTfs5EOJtuF+485bId2CCmJLVRyR0Co4NgHl9aoSSzUyWJz45fmA
2pMmE9tUafIH7EMB8NMPIY2098exO2N/9/dJ8gWht8QpqZSFbumVgZhlxFPzdPSQ
LrQypAOvU2wYDKIdevGFvIbH/Xh9De9s4emOQBjLacUnlPW/I+R0r85FczanV42J
bwIVxZqhbs5lBuJs3A8kOn/a2shH0gzzgVzg2kzcoKaHpEeuWU41qaVE6xtBw3xl
llLzL/+E1HoSo2+h1VB8USPWlbFCi9F6gllRpojFBV2q9iELVgfkE7huxNiz1Nea
dd5KJ4/lyvZv7W6wqviT6lDiHLn9947448m3QNNPkMcjLYl+IbgYf9cNwhb/wpxw
qAp7AXBiR63U0v1N53NznaF7yLUkiXOHWLTYW9hfptbORcLlwM0uTnghlobvBy2m
js7sRq0IBrol4pILKyFJujxu0H6yCcNvpdJMWR20U8Z8nlowof1VQPOHaP/lUOhe
6kjvayotq6U7E7qczwToQNvJMmAhj3UfVTk3AQjk3VkEDTCtFa8feEflsIdx4asW
jKPUAK5zQVrdC0PXiO/uc5aZZpu/iv8MYZDCplDuv2+PtfwR5mYozSBB+AM6XI+a
7AXGcHkhp+1KRTxFdkyX/qbK/CEtPyU/GVw0A+ny7ncVtB5BhvbCQ137/leiradc
cQlPl6vt314/kq5V2Ho8/PG46fw9fUHSKI6kT8U5GQHdwKMWSRjnKnRPZuPLigE7
T3q53+fqByTXctMWTl81valoNw0hiKmusKe9aLGJzFcVgbKksuGNDtc+HNENbAij
sndhWdru8RMvXcLm5gRV46wrXdKBPOv7pm3TZnWftR5CLIR6aAXYyTC+w6IHQkza
C0lbyN7UjUOL1zk35REAvqEncw+RkXQR0BgbivATG0VSZw/mI3PlyaEC1n1in9l3
Rp4VIwt2AGY0LKlH2T0rFXgX5WGUmthZmlqmCIswtYcqhYDoQjdHex8pIC4P2V1l
kMCxooeDatlbyxlo3yUIkqV4vhI/oC7cZmSRUeFYzG/OZl9F7B4q3DpvY+O3O0j7
8u+YhGGUggJUUQc6Auk7XohJ59Pk5vPm9QwHdgY0VrqQfLjdJi2/VGMY+uBkymRw
+YQHdnJX1t0WrPhekaWBthXyolVMpSEYVEjJLMPV+MMJT6H7GCpn751G/N2serNz
6z6fP6t9bDMnMMluoJkqD5lJvXyrX1R/MqLe4wNjpr/xaXw7vRrIAkhoBJOgVE6G
v0E1hwMCbR5Wy00eE0jOuHXTJRLhyuW+GKESeu1kiGhdk2Z0JhKNbV2h2M78X0vu
GNQkZnD9prXgN/4PKv1lzVHLFg/dbDi/CJnAxvQKIMN/IH5FZaa6GiAm3RZmdk+t
KBSQe1P35kWH3ubJ8p9dtQ6H58IhH/J1+oVdsQ5f10izBr7JISXISkxANwKFpu+e
ltnjnZEryVH9FZAl1ZlpFn9x8wIkZ0Rdqh0BkrbxmwhAQB/sVn5nLwyI9FRYtdf9
ynLsCfQ/pfvmAfQNK6ItUpxiYGuBzZ/rmZDl6Ge4xY8BWvI3yGqxMZxS43BosWPA
W8ckv2IhVG01R56d8uQaGfvBYE31OvBhr1IhEg8RWpAooooIMPMTTMP47aFB7EK1
6cJkhBjFMfqnYWg5nK0doZ3VydhWbeJF6gehgr114kl9YPwOTcnkWIeYTTlGim5t
vxzAdTZOBkvZNJ89YPPOEA7AfwD+jOhu+MB/482jbYrGLMEjy7NTIZP7nS9V19Vj
vrsJZhsfBcIwWjqE7fAIimd+q52X6mHcCbVZhWp0IQtsz8T+BsOlXml1IEGo6GzF
JlouzRKSzfuWTZlDhXIC0BVyo2KhIky9bQvsbVyhHIP0PMd7CxPxaaosoukC9vzK
ss/DFpwfnkBfDStyCaPO7hc0MIX50wUZDWbyCAwtUFS6lW0RoBpH4/LQHKxbYfU3
tLxYRgHfTRKQX23zTp93/etoK2TkQ1cE2G+gxOy9av4H/XGe5qk/8X3+crmyrZju
jzNHnaYq1E1Xokit6bupana1b+VOjiTtdrzNdeYbMwdrufNwKV5vWf8RxJaJ9PJg
KwhjJXwQATbMzbe1nHEbTnIt2yjfc2USWDYO5wgE+Dfj+5O6Ou+Tn2GSniFqsXnp
1fZyyRHxrYNiO0br2XYy5C8jTkJub8Ij+h+6OK+xQg7PZJJHPqHVKJUoe2oSvqV8
XWYgYvzVpyJcW/e0GbhaAJtklcLq2Mioa2GLH3GOv0sB5IGjoDTNSEAh8IhHRwJN
eIuygooUCJ07LKieJ6j2EjiNsdhT5AZgBdiEl8590U2/NQcNEhrlNcApRBtRKBZs
Ye7K2gPAgudLHUUEjRlNVQeU9bL+S6IkuCW2uss8IJOnbN+cv5nWQC3As6OtxN0R
sazjHykeC5y00gS5+fGjQjdotSBuObuH58ffn2zq3u8WAh7NDoORtpc54n1MeDCS
9Hwq6wd5ntNEtAXqy5dgAJv+yslQoPFciOMqyjT73MWxjCnGBaYjYjTFAC1K31Ju
X90CEiMB412AXU+ujbnlFe+3wNrTtNLat8mhivw4MXO/lQFAjIKY5HXN9gwRk1m7
pU7f4/lWCPnztLDsfrZlmx2Hy9CH0WRiQ0pOQjZeP6odY8/ZATKtsWg3CFRtsDu5
RjdQBSjOOOQzvcC3D3+0zKrHPnC13Ml+/odB2rwYDTbAobYDdlrZAnby7AF9nqIN
j9hpmsOHXhd/TVrpI1jNHu5JfjNZEi+SkdFB5V8A6NS2VfbBFHqDIlFkCu9S8Bba
U9FfI/Y3+TwpkwKO0CHy5aHd2UShibzEsgVtXQLW8SORVJEFqM7DAz1XHuf5Tex0
Hallq6Tsm+9f9cyiz/TQ4YxhrAHfOUcb8C7bkLxEWvrpAXWU/IXhN8NIqucABuVj
rlba76eYlw9NGAPZ0z5Iqa5NJ/9fSXChOBNwbZYElcp75w2WxOq0zjk687wg/qOp
hxrK13tC0BmcNrdo1ivTswwq2M/Djsdz7RNSR2BUjJM3spaH2FEU3JHCVyfLJjv3
dxdfjMFLuASrfhO3BFZx5WTgyFrhGK8vPLzi2WdpgY2dXmd12deMshIl4Tepunfs
B68u9BsUr8bg2NfTBMkKLoWtQsoR6nXxBuprjCRLj9brgh/6SVWXWBmo01GWVHAX
+NkiwQ/9DTv6GPsN0FXadEqaI4SyBscJ8lynJ0YQHJ//8y4cfIgffbdlV2K8f/VV
EG5IIV8Cv8ASSj+3IuivuxKbGbIZC4L3lbyzbSNZfox8UUcYGtX4pSz7+aAQZ/wx
Y2vf0sL7RaiyCFMC83Pn+kSEVSs0JTv+g+8MjGtgm/Os2VYK+MES2mzUlS/tKBF8
mbNFWB/E0QXenHVQ7cpg3UEGnftgXE74r1VufUhnWryZxObqWckgT137AyHqHfp/
iqCjjIlPecRDtMHRMN+ncKOEn0izowNMulaDb6BU7av6bdKSYzBRmBaSgpQ+hTaL
iBzze4wAlxsXx31N4nb+SlaGI9gx9q7349vpF0CAqmHwaI5pY2IJ/LKZ8X1A8SXA
DXrKTmrlo+830CJ4VNAwLIyd+tfj+ijRvXTdNxDJMuGM3Eqxv8zMBWOccGdcZ4Sl
Gq4Ht0qwRROTV9IcJbBgKoxi/S3igvX4nuCXw7qJNAYi/9fPzDrwbRiWwNv0SlgV
V20PHnOliiifmzqQUXXKHKFA1bOr54RuNIRbFW1rIStjq8eigUQDuk4ryd+9ck6N
on2DZFUULJdPTd7Uloa4HQjV7jZBRh3CQE2MXiDTo52992jolOil/h9sTLmSBTFP
cKMJ0giExPjUsu6u2k5ijJItCXAyC7zLDfz6ZsGsKOFA0j5HpaJuf7XtxiuSiD1r
VNAn35EWLwvEr7GojrZYQDk1kbeTyxmzTucb0qA2EeKGC1K5+rSvaWPdF9ABMDKO
rr8BAPEwyuH8469VWOpyP1dRofxBKtedzz6YZyGkm7AL1TTBBF8tkCNqgcqiteWI
xplLWHGKeMM8+cTgjgFKaR3n4zZjU5u/y6y7iMwT2q2mcjrNTNN81VvAy4dIdNmw
bwYYUZGck1VpEyPD79fVuCuAmF7vY7vsY7cZeyD4+8bBbwTjNsLW4W6tJaanibTx
suJBAWONXAT4WegqpAMVCa/SUrEx5grKg35udTsYP6KlXv++Eh7wPp8VpOljk4Cw
Z6EpHNh5M1h11QLOTq6vgPXCciSRO/ZprWsC1R5SlZAHqItLp22JN3bFu3DnWOcF
0Eq6yqQBmhrKQ3Rfkp1WBGh1XhByXBn3Nc2vEEfv0zRSeE+a/GO6VdSgdTbFAebt
iPZ6E/wsODtYnHYqyA7BwniA83c4eqOJAnzFSLSk+Agxe0q1KfVZYa/xQTNFrqGS
t5V3mZwzEg9k+g4bs+JdrR40tlVoxNVp8eT1ELz2AGVzJzPkDNQ6c3KBKX+MFlgT
nyqT7wbolIFO7ugnEl7eeeY7UQRGmG09VvhiX8Hu5osjsOsP7vXnZ3e4fb73yF53
Mjesft0AadoUHGN9jXGl660wO+GFl3MZWzJPFjzyg0QXOiZefbtmmdOtINXPCWe7
sLjPnycF+cZw+Aulj6PLAikMLf8ml37052jHMdgTGkh+kp3hWaEoI9nKzQ9jQpO8
YiAoPrjB0HfzH2GoePjBfgFYZiyWCh+noPOAvemvYWSF95l4luYvaq18foJuCFaW
my5WH8bpMMNrvPyuuBMEV/hFDTmQ0YQWk38jtX2Q1FWylGe6+njqAhSHe7ex/z6V
Td4XB3mnNDshvaqCyCI+wk7hyonWhSvZZsSXRDE7KMUYTVNlKKBz0ftRwsSsWcm1
Y0SQsQmqIFGpwGK3YNBkh79VeaaWEuFZsuWA0MGlqtu0BRS+KVj0uiCDP0s2FQYI
jN4zIIdS9TM4G1Edp8UMK0KhfyMBUFVPmiBxzv5x6UH9V2rvL0QpqSNNikNechf4
SmqecamLgrpPhlEoHipueicWQqzoKxeqwrXZko5Iv4ZdHFfFRQNHfd/kwVmjYkn3
4XM5Lj8HWBxwL1G6+6YSkQ4oRMGc7/fJQqJFIhqt71Uz88re7qMlRERwULRpNMxy
K8nW1nwvQZo0G37BwEwKZmvIC+z3hCkiZ4vr/jwK6tH97u9BmVIAY1V+FUFUlY4v
tiXZnIRBCATzYMCJoiSrVPffJFQYX3cgQXbnoCDVvSa7juQr+6bQS3q379IXBliU
+6Em28/u/b49dnnNa1Qfl3BG3OyODAhYGaXBdaM9Qkp3Psn2vEtPm9dpf5NYD+pI
SAMUgByVZH0nYXpwN87knXhpberJh6GQxh4OfzT+1DnuM1gpTnPQORP8WqiTdBYj
J3OQLzo6AbPNUxJJGwEA0ALzlCwMWvyrqih+gHZsifwOSJBCFHqVi2Zu9iTZl2BC
4QUrb51FW7tNo2u2fucpClS4b9zknRdDxx0H4E7RoAkvj7MNbtP/SgtyFVQTyLEU
6L+11ThIi6V90i2FzGgT2Mk4h4h0Q/CPPUFCQP8MRY9I2z1Z1QXnsXIzMQFU7Uuq
NT+tq7w3Htkb2v95nrbULD/7IQGY0oH4L+IM3BJWw3xlgJK6I7ySBvusKXmBeeH/
KCSdMIikTUANHuIJZ22p2DJ8m8M7KeIqe8oR9fMWu7LXEHIq29N0/SGJE7+buSgY
GTrLNu84KHmrC3QXvD+jdO1Nvm6Ilh9zhy9+myyKS7E5ZooYSgOGMnOdkr0dtGJc
ZkK4VdSKAYdXy4tvU+dmoxtI50qpRvaS3wkVfFnz4IurNLM59qi21JFz5+Ef/hQr
2cVDhuk4y6Ep19di39CuL7mD/72ZAOESrXyFdohAFYxoMIBNPq/di6LCZwUw9XSm
VROCakT6Cl4TwvwsRVe9j7EHLyoFWt0jOWu5zSy5iLKiih/0PQ+3pjHw39YRCqsy
4qpUD3xo97s4Z123EuanFJjucXQjZemrSBrVeJS1y0eDPaKgE7iaIihs9uspfA7c
UUXjul5pMPXTPg4QfQ+nhZ9bvt/149mGwhoMWyOwdl68Ewn7hLKw9zd5Vm3vKnDB
ek/nXd2hbsbxElidiieboWEmWM8/dT8XZ41iGm705nAC1q9Jfv87Nt8XpbckAKwD
n/fQkfMiC/2B9RwKw+gkwCVMtNWbUtaqn4yuEI++XscZdQs84R/glEpyeNc+lqH2
N1nHRjdaRyYDoQ/QlCAhNUYbyvAR3JMmTAYfD+0tC2+XIughBNCYK6WqOHRxeNkB
BbLkrQnojmJhUDS1KavIhds+L2iO8Phb1u+wF7HdUTYQ7K36KKnMpSpN30+qMai4
pbCH2iVyeBQn/Kxtj1WBdpa/dIAI0JYmNU5Us2vTVPplm4wHDTB7LfynLKOvwkRL
WP/9SrlZJlKsSiLH7jbhI8fTOauzReJVTAnSks0xuxX9M9+B7YK1PsXvSoMTJqeB
SJ0BmdZQCnp1s+Q0Em+5gb3Zu8Hv6AE8j4GEgyflsthCSgmIDt8d0C/9UVGiZKC0
N7Dqd0gKjHsQxT12qDb7tU2D+Ki/DxWRyhmv8Fsz1qXVFKc4PmAqAQdodtvaM/Rk
qF0DWjpaTPE7zjCyR5EyGB5pBpOP68dyrTmIWEcUxX2Ij94t3rsEDxDFQvKvEsjD
giuAcALyChGiIROOocUh4l50GtoHZtYST2zjVTcG+tswLUe6DqF5jKCsAPsyKIV9
Hm245lV0i9jP1WnrpYY+56McQXwNT0W7oymKldUrqgc1Q9NJ09DIPb2hMs7Rg/rI
pLQt24pukM10zLMNcpY0zok5gTLIcCXobO23GE0WJTQ5Nz9YLCezoVJ+j95R6tpL
DwreJMFN0ZgAINiIevkekwraJmGUYQvf9Nusb3bQu81uJkZt+qKYA3z9T7kGiAPA
MGXil5Fnx+SUoUwoMSf7hrJj4nJakunyINzG+hVJNvFV1UujX1e0ZVN+dV82r3XY
hMnF0MR4U5JiY/pGCx2dtSV1W3vN28tu9vpJ7eHs0+c+6sQAPi7mI0xPT3YSa+7U
FEg8yAKPc7LU4+7Ywytymkdh3Zvw/4xE36MXC+XcDgyh8Dv0O0Ac6JNbvIQesAjk
TisRb9YbcUdtr5II+L6n/yXVj+ureRwmomRqIdkfcOAH7ZMbb6FRW30z5TCLrjmn
YF1FmYGFyplmKE81CHXo4rcuVMxoeawFIrxbjpbJvz3bSL/REamQn0dwuGS3rPRd
lQrD8lUkfdOrQ4sRvbEcrNrmV6KVMMz+az1why5f48xyycj3uvW/8bbgmybjtfOQ
RGIEpOJdWr/AdfK8pRwSMQeD5MHV3Ag5uCDcAl3v/K/Ivldf76Z4Q3SBMNbKfRc5
uyQRKTEmwNMO/9t05Gbsr2AYkqJo1pALIhHzTXvkwr1MZuv43KKE/Qtw1szBXaTy
6S3GrNUIorQDBI2JbZn1TS3luoE/XNrZnlsABRQQ4uknbmu2QItEsHD/bL84DUPf
+aUy5Qre4OVzhhdmjxqScRImSIyTGM4LPq9dEImFho1waHg6N2u8g1+T8J7lI8yA
1FrIH0KXVUfz2AWg/m6YFj5wwXZJYq17SjZ9vUQJWPMTxKw3Cwb2kmYTc2dh/g0h
4ekK1vfSAaphnN/hjKoywWIgU1pmfjC2NK1mu66Hrq/Ujf+U7PeT8K4C220wf8oO
oof0BLn0Xqut26Ptr3Vny6Z1s1jqmOY1ouxs5JCfhRvBQVZC2o/YIzMP+GoKXJN6
DZRTvi9oKQnWlyPQFHUjxNeaqboDPdKjMEtomSCaUQ+Qu7Sog9Tfn8vACSwP9N9S
XshLPmanV2od8nE9aMr0Y/R6rzJfOf4kRpil712u/P7gLwL567OjW/hjqa4wFfF9
XnNIKzNq+3E527Jw6k0IED2qWgu9kpYYPNcxXVHTAkFqMpo53QI8w4RJfrvwWetI
bHhAEcAPt+yL0FYyC9AuABnv0YFUuACD2DygMrMqyMxuXvkmNbMnKSaZLuCI5K5M
4cn5Q9ZejTDcZtsi9/FbeQ5tCBVN2TfVzNJliLdcf5Ycz4Lit1W9zxRC3nPvAV5E
yJ6xUqo/InLW09Lt0amh1s7SenTLT4fucb6zeSbT26uuUHBe1n/Mt5yyuXz1cKRd
NkIDebQlBylA4zgcnsffJ5xdf5jTQHDukpGVkR04fPODVdM/ZOLl1Q77rlX4tKpT
SVyd7aiwc4H+YBupENiyuEtKMJWstQogrC5Rq8yGVIZTTX+cOto5GMOvg4zkIIGI
LLKdFGVESCOJQkcu4FjYL3s1gUfeotIvnk5haSxNaJhII/fZjPO2dGTgVkAPco0k
3W8NFlueFh/JGKpWrLmGcKP2gCUqhN+jvBCOf/9PdJcvsepWUYBzfv32XRQ4e6j/
rIj/tAtlHg8b0C4pp81voSG0cGu+3danVhuFhHn1Y0dqMxTeoAEg9iKz2zuensBs
qOjiK580BOV/ni2HJJXtmFmO1x1W16NGmi0BSoKfOo2NW6nTwvXqvYofTQsSg+kv
tG7m5MyJ1QX23O0LgzlZUJghME8WBzQ770erS/SUoY+CUwZVsgE1rsdC9B2cr1dZ
HLVn6zaL8gxKwP8woFOb20Iksi+pPpEIYm8pmO9uXGhh5CHoUSI6nw7YWdF1YpRj
7nwUxs+7aVwOXWUgZuh9NIHSEJHJIodrkUU62v3H9ibeIpHKF4b1TZmuve2qrcZq
i1uemqefDlrhM0eD25YbouuK1bVN6NajlOlnNC95Z5IIQ5dVMdW9ko9yZqfJ5+4/
C9tZbynPgwHOjQR9ss6n78CueMWKctsJAk/hW1SbaSIfdiJxYsiHdv1FB3MnlSRD
4g2+hJVdjyEPosxnFz5mm04iwNBmD4v3ZWQojFzOue5MGFM0oTSMR/TeyQ4Yd2ds
JmSAkiJDHudh2UHvwwyLWaGtpuTcjIaW9t2+MnSwm65Gfo0IcWbBnWf0rmWcG0cv
CSTuNnC51Agr7yGVe+54BMAPQMggphPw7XKZZD1vDh8k+gYXnLGzaRzLbjB6KMl8
abosKyVHL9ofomqCccjMRUSmJeuZvV5VZlGqyuGB/HIPJutLIDAxzFmkCvZTQDKt
l6TpzePPGf2mJOh8ekfOVnz0rbIn5IX/o/MrtoyFtrAnzAAJMUWr0kAwWUSnw3Qh
26v43Bmcph7QXgYMo8evRP+wfjT76/+2yZqSKPDCuL28Bcg5pqNpWf6I/GGKQ81B
wb23sbmsEn65EbTf4Qb22L6X/pizhtegGAMFzpj9DaZtgKKgWQa2pk5G0k5uPd1q
3tb4SIqQI912VojnMRh0EyqqxzbGT9G1YNewF32dWLL8QgN6SuRopDpZCYnucGpZ
iOtjQze5SrnpdhLvItdLKuIk0tm5x8iOQmTppoA/OhE8OXDTOP1zvVD306jNqQf5
aEpFf4cJ7xER/fG4OcqJVOmbdM3/yDvppA829e6CJWapW68WbHx2tQYWDxNHLhkU
CJLVzzaPIb+l4OZ6n2qNIRI+EMJAILUhcqb2fICMYY7BMO23i+s62iLck/nIcMb0
Cos8Emhuc/AbTl39YdZDDviRdgoxqjSwSdzidwrOBjdOC/+8QUOwi5gkmPthefny
tDiaGTaENGjDRvPJ908xhMAZl80wLKOdJRiAiBI+eYpsZAxJa+7qttcyL80HIDhF
k4F1TSZhVgYecGYLbBiWwluMf007BBWNxzcxJyd3YooKqdc7UKRYpSyVFDX4dK0u
3wRTXGYcXLwSa9oEFnUaSFhuGimHAvUw3V7w5jHFD+SK4dLremttRHPac0YzB0b2
n5N0pwo8lVv5c4RaGOfysyxAsayDqM7txN19neVoBFffmL+mp+p+6NKd/5yCLYCe
YBApi5eTBojHnpxi3rATgT0vOYJR4xrJaeQDmifU8PzeTM1KgUpllyd44zZ3FJ+I
gGK9aa+eks900xzCjFI3w8sENYjV2jNHgA8KCfoihYoQshK4vcRsMtIhVMiA2zCR
EssT+RVWXanO6EwwgcHhCkEEwSbo/DVf4GAY25GVeGLX3KBYP+yRKtg0SLeclVHN
0ZiUgicwxFsaMlbF2hsOdknyGXu4vSU7Gkqpq7KGNXAvAyjPm53M24zCF8rLmpt1
/z8elGW7q2eIBQ4TYWqQhRHZMRBxPI3ONKSl4OpEX/UPDYhsBmJdnUO61swiGWzG
WpYieiTamKdNsKjqep3bWvxRGcHgA0uqddeQtEyZ6tEgDv/IYZn7HfTMuoWnOA5B
tJs9yuT1olsPGwa127FfU7EPbuckynCU62TrSZIqo4AoJN4zay+iYYYBAXDhR5jv
YTctV2sdf/0ASuZeij2DzuiXfHetUFNcFart3cTmoZwMmDGWJn363xbyVoGsEfDg
gUvzCWOAYZiLPy7A6i2kub5sWOex2odOEOHI+yplJPI0SvjMYN5uCtbaW0iTVSD6
69gVGGqAza4rbc3/bC75fVC+3/mSygQGJHoYHRTER6eALI+4e7mcSofgbv3cmI5h
NubFdmUL+A2wWreC+8AdjVACG9aQb++a6SoqGqOoyRiBHY7wTTOnVc2HdiJH5kf4
sm7RFftybn8hYjmpJf4seE4STCC2hdPQyu1i3j/CgBNOzplJQqe8/8dhSr42H5UH
Oz+CaE//Gm9EgOSoVwG94Ju3GSenJ9VF0byf5Q8HqWqR3iJYDsDr9AvxUd2r8Rqk
DtbT/CCSFE7I7f466wHhOty1Ea+6zBwzOWFY9JFI7rZc1aM9jdFn2gbMEvAExP9D
lyQhbgoIt7FDyTtLKjcwo4TddjaMj/vxkwTttSFrOu6zfbkUtQGeAZqDRp9gF+Gj
jBkpIqhWnRQPNJfP21YFNp8kVP1q/kRWinyh+ocJZbuE0grAiTSXnEn3KPkzimbv
/RQh+T8oeaQv+HgwUlHLBP5hE21q2SNZdkWSSMuF2lXfdfhHcP3/aUp834lSTpt/
bllam+XbiEhrNbrFYvKYDMGANwvHLaAgVaCYjoKFASI8H9N4rZb7O2d0IKmJ3lFk
kc+A7UDjT5sTkOy+NnKJg6L3YEaEVwaC8U7v/0h9vddJp2HsC+J0DYzRzpltMrBm
TsvZjtgnROMMZeJO8TwVva1XCz+aIk+u9Tqijl1nk/gY/+cP2EJfGQI77YnSAvbY
Wk7BvqVYS39heK3ojqSnA+nYt2kc3VHBf7AsoHKdE+HLchfakyLmLaBCwOVyPuUh
dexttzR1phvp8n3AJVDGiLtXh7A/vfKnBG/gEQGKC6jds4qQf0Plf7DECCsbLmM0
YV4F17BMhGMvV0h/TFuODMnPY8Bax6gC7ha/iZ4X7LzmFZIghyata/vb85paJDV7
F2zrjemPRZd4sUF/waQg/7QT/iMCQdlTTyBf6WqbzVyiKMk5tSGtWkWq+u+uFDbD
z9B8VC1lzfdQyt5M7QKOd37hdcT2PttjvjKzUKfkZ7e/qesllebrQwCEZh/6OPj5
yCYN5o3NlgSEG+pzY7Alm7S7j/fKvpXv8vjJphAiF25AhNPE41wFXpO4YedI1zgM
JtOYbAi9q/PrwwjR1U6HwZsQrj5HwQCqeNm0zfIwE54QnLylcZssKybhdVgbK2yz
/X8yLk4SXhJ2OZxW8B2y440eW1mF+Fu8496nVaU+nqxnuHTjKucORc39kE9NIzk+
JHGZ3KtduWgzgK1JRIslckchDT5zGtFimo6H89lE0BnfTDx5Zw8dAljzThRn6AYp
9AhsDO4kqR0MSMhgPyFzpmk4uo7QGDu7s5dbHZmzrl0huB1AJMEEp4D+cuXRO4IW
3tOVSYJujJqiOSDDB20sjnAM46svsCqxEvslEfypwpvVqMI6udnOmgcgtsdtKu9F
Hw6iOBL+vCoRMcX9cIKuUvtvUnK/jshVRYvEQI30EhWJcT4GZVkz8dVqEa7P1YyN
SpxueTIL3Io5Gc+bakMACsS478S9nqc2OYYxZO5e0XxgfotHy1cIJfVjC3F/sNGn
1v9rzSLcHUK7UAb1BJsPuej38AmGGmTwC+uVmvkk8q0NJgfrxNz/aQrKkiazuySs
fCT3dhoFxuYCZV7fv8d4TatOKNWkXSL+VIiTrafxVs6xtti9/N5gjFK/fdbyNs98
PtSefiq4CXbXzOe9uFGvbcB9qzaiHl82bzcNUZ7Qhc0douZTMASAu7GDH4lO1LGe
rbHDEbo8Uii0PnRyUQYHkZeNxtKFOgwAh8/BIDi11NJz/eRJ2WoxBXvQ9Zs30R/W
m2n5hug7ZE9QodPYDW9y93ceVQxWDev4+kMz0PiGJqdVMA3IosJ9EuC/aIfsWTEo
A9jIv5RSaj2Vlcv/pwGpXvKcEv9jijbcaHhTV5wwd5GXDQaFK1gjWQ/uBUfMWYaO
nubcKXAq00d8EJHdNUZzxHyBsVzEVD7sU7/Osbi5gVHVGn1/vUOFxFLKreiqVKh6
m0bBJufRK7tZ9EeurFI10d3nqX0tSyfzsBfLrgr+e426nWwh+T4LzJxpZD6NYUX4
fHNq9zUOC8sVzjpYACrpLMmStPLdMsgPAFN2Os4Ga5sDegRC4iEnXjH2ZeHxAIkV
D22Lbzg45dlVRZ0MB/ewXsxbqBxsZWnwxKs/ixOsmXjTUzrLqHjhUdbL1MZKdPHT
i6aeJR0AeAuZxd4hcAQt+bhgoxjuDqlmohm0Io+Ejo1yPKmaiUpDbSHX0BG2WIa6
D7QFFOVXdnkOhiHV+sDeYgJ5suDoweOOAyZZ+OWU3Tazwul5UfZKRL0oA0btu6KJ
GfFZdBFEIX46/BDOw77QdHjKeWwtcl1KUrCCgvdtLSIpcnkWCpIMu0HMd54g9W9s
tWw5jdnPbfVjJQwB+n5OUL4iaKFR4EllnPzlChLAiboKgvn5Aq2FVMykAUuMIZVd
DQDw6EYd6AilgtbXavc79Fi3qww9C04kvH+0RgcCCmphenLD5nhhfRZGjOtm3LA6
wW83uUFtii6lDahnD3t5T2ImF9oMWUqvHWuOCcKWfRG3s2MWzwhywZeQ/sTF7K7Z
go/+U4Ic+DHL5ZNyUxdOXt17XGZJLvT01zkjKUcyZ3vg+9IEXlCNDbsem4UHBeHj
p5+Xo+n432ogRT71N5Qvce7GCev8pz4WHBmvX7m1CgJiIdCgRLHBIz8G/izY2446
sgmYuGuUhIWjdPGAByKrXPAvXZ7vzSwd5QxeMkPfbbsbBJwhYy3BJ9qfvBP6UQWq
gQUMOHJinL9qI2xYmjfF+L1WWMTS5+CU/2q6ds8Fsc+kvEbpqAQIsSG9d27P0DBx
dT1sZeOT82oPdwxecS13PSN8ZWahkvEads9DVhu2SdO1iJmtBnWuXHmOfi63YFBa
go9Y5enRJ6IB4tn3zWHs8HoKekbK1vrCECi6i51VLWjgilfoYkRQth3JQCIcUiIE
b+LxWxbITnkCgMVMH8A1dO+BrTJMkojEdUp9ylvTMaPS2KrOQ/cNeC2BR1c5TyCO
u6sE4QJX/xwJvfe5IgulLWbXM6H+2uIMzXV0dd1wUk7HXemtrHjOpGCH+RsWQFO7
FGlExnuYEVDtopvBqVa1aoMmEdNxsktyG53uIu/CXOmNRYq6sJ630P/jQ7wQlSJz
hyGmUE2e9iM/fEttcc9TIXUx0ptyt52+VQ6t2w0GrqOvrVrH3YiRaabUPWxnb8WD
bWb9LwLhajN+67Pb6VxK1ol7QpvL8oO5kDitAI55QZRnE5ahpq1gYaTnuTW8zwin
4BuHybHmkH0d1cc2pHKD7wgRERPF6B16hbQyP4J13dmJCU7qGQ5bxXpmy86YbUr5
6g5jjImGGYwaSpOg2hYdvslFqPcBc2B4X3QzpRdRfBF1ofKgaGKhFTnQqNoHSFT0
NP3L/r2iLpNaaC48nZEymA==
`protect end_protected