`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 5952 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/59UwEX+aE7FohaWu0/8IpTj7mav863zUNIsgIH2BWb
Abd9opeuBjbGF/waQMI2vMJTwD1ie1YueHc3nSNpEh4OXp8P5ybZFY89uyGz3ztU
W1EsuUnchJoQgbHZ/sLbgtGRgsrAFn+ZoIeGN1d6RAF2wAESJmYP8zw+p00RvjZ5
pBGEHX7wooDexzkaqKS5Gz133fVRsZViKBvDFt782bl7eRP+EiDUVLXyNZC3KTRR
XOshr4WaR/+Jg0GoRNSj2hpRhE4vrnDPmr6guYt0rxB/xLCYeB37e/lkpbebtSOr
sF7c7T7mjsUxTIlWz6zMDpISsTWo+bAsO23mQgAR/ifwHzLfA8JT8TOANSlAN7py
gPlDYlgWSdWuZUlUvEog9ab0xsiFf+NQWEGlU0snRpGuT5otGo1SpKv6j85v1n6g
mfftnPnvgDzdKFhyJgJd02NAZCWgohY/k+WGisiDRDS0hco9kNdQVolKnRstIviA
HvecgZ41HauxzlL5lj6uf15K8vtotHI1xrhnei1VfXKj5pQgrCD+BjWg5Qmhmsex
253kvRy9G+UDyv7ZgWtkgxf3qaZ6M3fDotf1GdV2nJubXsKsoGZpLOG1Tp4KBOGv
TUiGntD3zAD9E34G1LIMOJQEO/dBWNzk/wM+fYkV8qKUlyUEaGLThCEQCYZOHp3N
B8ThyMm9J8j78LkxBjSgQTXfWVQkoXrDVlIet1KINuDX/NVOamaiih75LUPkqqyn
oi6zE7h7+6zD3GFUvumSy92Kg4uh3F0kLVpSkM4Gs96YiX2BPYSPjgaEVRn+qu/2
Jc8uYZDcu2nV0QZnHYw2Njn1FDZp7+0EYWrhlBktQMwPSa9VW2PHqqf4YT5iQ8zB
UCNLqvb+mspC0L/SMTMBEPD0FJ6rir5SfY5fzqNdaGREFY15wQ7fZtACGskShQ3M
n7qLoc89ziH5RV4ryh/phkU1Xxm90IO3C+psYlBCGYEHqbvp6SY5mszCRVq4knAl
LvqA0Z0uI6PNmcZ5mVyV+FRcO7FcRYN3jCQGYzJmpWtZJMIrpZElH39t0+jlP0mX
wQ0Q5j9FKEe0V7PRaiUePeA1FF4pmSbXO2H5m4Q1f1nONh73JLhpgqqaEYQ9lb15
9XuetYbODDnnvkObDmqbWbmvAysPLfFFCy0dR2c19/He3n/YXIQoHYySDmhx5zyq
LojxdiwGuaYFDIt9XBeMI1MZ6YXseRFzQgqWDuxYnoP8lh193vspX6SU7q4J9kpJ
R9GPYsCztzcheItZ6XBolINNPUYN35FfK6479SyKrvmbJYdnB1q8wB7fXX7L126f
Bu7wPVezvujifYLYOP7ZAv+gs1hNFVVq8yykbv2CHMD3q6oSzopyQcRBKOi8fulo
KGDajGr2uCxZSEVl8cu+DSTBDpU/n4U3GAzM48j05zWO3EYDh9HYx+gHfsFhfkKt
Z8bnHvzHaYH6emxhki+ZLlKv/AHLBALKTLStQliDxTqU8kwKJ56GjVPOIHqLU1pU
9y6BTYssjzliLMGR6d2N5+jxQ4A5PKYuyjMvp3OSL8HcWblCRFpG0ZXXrCWRiiVY
ROkTxqHe7oeDdOtapHChhK9IdQhFcpz0+2DL+wEBXIt7K9XmKX6g8rXpKe6M6GcL
pcm2diAbbLfCrunsi2s3Iz8/DXQ0TFXtWWOM4tRGaI2OhTkumR0h7b5jSTW8zgVl
pX44StUQJLDcSk6lXZ02Atf0xsouUSEdTL2SRJehwBSMTTPRl/aZlnbgpauUs41G
4FiWgn97Sy4ss+wk8qNNefOFSm83BsPZ7sK3F1SgkCJYwGU2a60RAo0QBxbZYmYo
5iSMZriAHRtY2I58PauCFb4uVyP4fAUaZeMTAGR17tYLtDqudgDU8tPtghlHV+Z+
vd19LfINSigaGFuKPkqqYYg8q92XZPpyfbARTiT1wrqVhPybc+QzHMyAreAHD10y
4quKYKxU8iDlP2TLI9iKhUy/KN/ywKrXkRyD0VHCzqpbiR5MJ1cMk5FySW3M2W+g
IrdT9uZcuUUYP48QQCg+2LyT8ROTSIBDSdHyCdfuuV9QNmKjFK+uarGaUknA+4Mn
aM2EhQO7fUSVqbAw4wNl4vV1nt/Bqxp7rlsCEow7BVzbuTTneSmWKFgy9SAkX2Tp
hohGlyTimI+oxB6ZptI9HqUhynGKf58DFsbll20I0N51MwWRyoqdRm7KZ1jskqDv
8Mnz8A3YvhyNimk8KDY4y0cyO1cZ0VxUvXzPh35QKQII2WdejCutKOSRYJkMlsU5
fAPTwhcTydQo2bGzt6in49UQnbLDpFpWxvOBQWk4w9giavp758yt4Oaw+Dga6pzG
hfBRO2dRS30PrhjFWaHGUL2pNLwLaiedZjAqjrc2xHZbYNIUmVPELohKWmRLrkiK
pu7KkvQZPxdirg40wuClHUkzLRTp8SO4Bj/mjNG25ToZEyA6rCuyAYsltVL/Gkjv
JH9gTNTvjSKKol88uXFONh33nRMyI3mTixCsFk5GQ3Wsp0Qm2cvcCKYeEDGlDtZ2
vqQOX8MdwbgGm6HhFaQmjz8flQN7uPSni6wC6TBjEErAEbH7FJPIbmQAr5Hu9fzT
WhnZma+O07W2ZjeZCn9dDGbcHx4iA57raca43jwTxdJk2sCoaSmQoMiQtfUrwiaP
WWzVYpuGmZJukDuvHXJKlxnobelCXSTDTMtUMOZ/JkIEcQRNK0xSA84JU5ZRc1v3
P9E2+PyoXTKedgURfKH9ODVzizLjGeGebmdkuNtXBm1d0e0ATJi5rpb0e/dbLxLH
s4SXKS0hRVRj9pEZqmoghT4ken8ZB3ug65EH54VenWPTsLYY7tDgb5aFo5WcM3YV
NNMvW+hSr++mRJNiwwzGZ5ll3auBs6J2Pbr3d4OjQtKtb/NjpXL1mz6BpOgM46I4
q/SBfq6mUaugqKWQHNd0wMgC+R+DN918yRNUeZTj49TOMugv5Dgo4L7MiQkHLM6Y
jhV/Wt06pPbPnW7AyrFGre3MPeomT8uss4bVgGN8qkkvN9jCrbqJ+GIl+zP4/s71
6ElJtC/QuI77wlwNo9yWmxMUmvE1xTN+T+JQ4tqNp63aZ7bl0ur6g9+4YjliUWZ7
lhkopJrwcC4OBtBe45rbVNuxrIvyz13jG81EASQDYqwidUKNTAJ9eUYiHcGswpVW
DsIZHwBNSuhKyKvg64x1j2Ep/NVMzhR/Oi1ibSZuEiKEjtX8GacRR0AaYAfyn+gj
wvb29TDZ8ALa/SK7gqWRBj5f0yDzAfWvH4gj50PD5Kj4GdeNTRVDGjPgOBicw/+g
DL2OBYbVGp63zPvReTH3Z6ztU6DhjvInh6L4CJdO+VNgAteuX5lqifkQPQPVivbI
aD33NWQP0v26UDdWXTSriX8U//OeL4b07XtqRyu2fVvcypbdiP95UIoO/V/1fSdq
Z02U+yO3ldJ/SRNbixas23sAX3JE791zSzZwpoXZSmCQjnGK+yZVQoegtg4Nwvqi
GaJLa/BYWnRXBEhoPfjtaETnRwmpKC2t++aXv5xqxDL3jQl4FHFxnOmSjl96LQWY
9+bY6iXNtep4kXpykF+qYte9oEaqfIZ63SYtLpfEboO+Vjn0gkOmQ8JS2NEYC6Ss
s/jcCPBjYE2c9j8UESM89oHo7ubStQ6pQuqd6ZdDivU23Ln0j5AHfDGw2AIZawO6
Tzvd061rx53qPYrIO4YxI9eLdTHtZ6Fn8dF5grpxXFtuyfQpvERABEf6qh6D9F8W
I/1JGCvFdU+qnzHhaYcJjRv7TOSTQr41SmS93acAyLGbVsBVRAjPrQRBsFB1MXQH
kg72L9bURLzOZbqAy5Wb/LoNq0Af/p3q2yKQg3AIg6jrzNpAsFVSXaNsbYynReVk
kzc9AtGpLWK85WV0x4uJ/yiyrcW7ak61Jupz1tELhN2oojODI9o0LshDfKqys2AT
/FMKeJSTkPs0heHnzNiAx2lSQcnwKwxV7hec2BFlcgBlI5ZxgSSFSlF54xuFIV7h
JoijR6QZr9zBhZSc2vdP2LH4IHUmb9yF7mxH9Eh1mZa6lQK8FZFFHcNtnx9TCqXW
f5SVmfI9B+gDGtkxj0Zm+fSozOz2eemR5k5pH88C3xjjuIKCeZ9QYvOJhEoZsmGY
MSJ4n9L3leIlzjBqsvGDzDwX4QK4nR4an2vrjYRv16oUP0j3Ipw1hGLgM5SZ7TkC
x0V9HG1TnuIPFuVU98XQjBuhjGt12o4Jz3ahXMxafSQFW80aqLI1Vwvtq9ybBk7N
0gJihniU+7+eHOwe7T895uGC69WpfjH0MSCGLQ5mocuBqOM/VvoVnWW59g6pMO8B
vnz33i4pzFed6i/EiKg9mvUcgI+E94tvrx54w2wDQaJI7L++v6Fefty7abfg24/K
F+GSl8ebmt+ipoEIv9JMGF9xTIexz2JLMAhXA2o9YyMXmKCi5Iotdg6uSkXN4aAP
amQzeT34vET1MMLuJznJJMrVBTy9o7rBkluQWwEs/IpTeYxSAxBipGgb4LE6JLd2
bno85zM/GWNb3GXoEEPc0jaRqVAV9ZLiEebE/2B60XITIO7vb7mtLcVBK+VZQSyH
wYmllblhjYYsIPQE85U2IobkDW/B52PDABzKT/qgsX0XqwiQa6zXWFY2Q+s8Oz82
hmhPzuK4v3y+XNqUc03hdRB3dn41l6GL2zyRvgDUWFvg0GJaGdvWVdDHwwKlVYS2
jCv3NEm86K0L3x+MFw3OOMxtBZVuCw0/PtEU5u7hXAbhflMirgiMjERPLKLGe2Y5
B2nszVSmqVYxUcCgmfdly3Tg/wy8WmTE5dEzi5WY0yN/bOH0NMnDeiulFaOjDzuS
zgUG1iDl6JkLac5Cft4SXf/RaYPNDw5EBF1iWuL5AtXgTiRUYFr9BVA1jv+ZqDhB
7KRzR5QUX/YqaqPbGeSOCPQaAmC8Qjbc1pVYI4lTO0YEGxiW8lIaaYnAMvJiP9b9
9czO/LnHaJmZux1Ndg8waV1Vx7Q5y0XEGzhNMQolCnW7qS1gmmO/AW+Wdqy9WiOr
w2+Ex775jmfNBTrbuNMhdtEYvf9aYzyLgV+qMOuQEqmrcJ02ENQD3BVh+n4/Joje
0x7opCF0EF6W9/sNZBkWbYjyIxkOH5pd3dAL8In+cHMF/lcge6kqV65r2n603gnL
Bh7+bnAL+aKfQjTq9kKSrfJBik4m7LRwZN5S7rlu3XEaKG320R5DDrQUNADIm7/f
y0aX90n2gnJL8HYl+cHjlKKTnm5yzmn1O5Iaunxmz04jngOPi70lJULiX+KXzW4k
7PblVC0XArDO3CRsEL2YndjxXOxiPpt3ZOGbjMMEvqBpdDCxDj8Q2c8QyD92jm5t
rT6IT98+jls0QwzRBYohtwb8yZVOs4dJknleCvo55LEQcLMAea2UDF/QnB/nWLIr
hDsSnefhjaD5pnRtxN6qqYKfq0xFMNd5Y5orxF6lx1C/AcaPJKNKlo7JvjorSVHL
mBm9XiiWfasIobvkEhZfmvMYh0CdL/W7sLRZXoLZvpzAEiFbK8sbIDTLtRP3lHKC
HdBygqN1MUgBAyKDtgSET0eXFvEKD39AzwP1VOJHz4mhOyvFAUJJ3EFgopw1M2rd
gudKg2i7/tsn3+JFHK+Y1ejR/ZXuuJNEH+XnSSEiM9FcE5BdeXynGNbI+AjU/pML
g+mTKA9DkokPyJAFGQdRpF1ztvdAOxUWNPhjYrnjNcj0ozEJrpk1+e1y/7TnPB0e
XMUslG6+/+pEDotqVK99SNJx0AJxynEtcdRREzOxygsLlmqTEIqbOV6FE86yja+I
xUBAdTqABNaQ0pmYf0AAs4mjS2LMCAp3Q02MhnenewtgUcjfVG9w6XXrktZTjr80
SPZ01EPnNnRa8UuknLkl8BKH3GyeIaTF7lR2JtZRoSKFVYgiTbtiz5d+9+0GFmGk
3qaCrF91dN5AkJq7FLLHIdVP1Ch1u+APf5LijNf9kqAmnugDRkmtdOVkCLHkDWfT
IXJ7/fVyPtYqxPLla79bENtvfTZ/yvwjnq/ituzY1lds32IqOelJih5S2vdNrcli
mRIAQ4JVGvhRoAi7pH1eNz2DQUdgii7ngr9Gx3kon7vRNUuNNNgsnYlUoMg2PsQl
DgZrRvpZz+Zd8+D2ktTL6wX6OI5eCc+Pfp0IjHj/kS6eDMEGIg63OOsEdBwmOddV
OqCoZo6/7aMXQMLnz4tUWCv3T8y4n1ve0xGiyca/DzwKo3L1pb5AghoNrAWK+cEz
BbSMq77QvQSIvX4l+ZBKGnnWbjIgLx5evkK8yfHFjykU1BKCUizSf7K7pQRNlnRe
bppk0LVHxeBMzfbgxlGa7LcNWMR5oS4wL5TD+N4xi69lvjLsVMIf6XRUcS7iE7li
bwjBw/EMKCTdmuvTuH3VXp29EtoYONhDWE0X9aJdl9s4mfRH63Wp/FpapmCVUllT
i/YIdMxnU3ITYc6ovxSvnuZxQE/YjTNAo6JAlAOs/xZuAmTzljS5LGZWPHTz8FUt
lt9URNAUK2XIPSmnXyysuYbNdZ0eWkNgPnTlSoSlsMzhSWvvhyOFj0TE0+89YN95
hhDe7wsfS8l5QmyUmYfzqx4GB2nFgjIqCg8HvuRFyUYG25iKiHSXRUdtH0BEyP24
Xjaioce2Zahr8Ap5BE1NzkPVDEUq1y3pl89LXxfa/zfxmkRoDcmJ8dfLmGsDP3vy
nWcriJzUWcMor/lJxBJaA5+TQqjSADlSQ8gPnIkFAwgj5TRISWUqwyoqKR098Mii
HIp8pAByEmQNlsInOM8/9EzVdJhPJ5IDMvhY1JE1ogYUfiOtLwYrtEAu6bagvcIz
QTX/Nyhz2a3+LRXItQbmkPg2Dcc6JVU6/EQCpMlNwhox1SRS/YtK+cbMIWjSwncy
fQOn6+wiqPMzOjOXIGx0qkUJdQBXC7gyBvPpgyFiFSmikDqcYldHoKc4n+RBh6ym
9hebNj/JaFXTxhqIhlhUU1udcR35YFb2wPm76EcfdWOEj7pEubmrv8VV0sw2JyCq
zBT9Ey5rNz+nV9f5PidciIZqu9L9bUaTJ8Qg1dRIdPpYtDJ7b4+fOs1sGscG0nBu
eh94stvUJeOPVW0hsvAgWNXzlk0rbeCrzKvydNE390mReLQKd5nD08u/eqdeuIeu
1TSguUCRoKm+TtIfr6tudfTQJYoFiHbMwe2wO/iAkJHORgoYpeZNqXDSORdFs/RU
TCBpB2xdq6fZ1hDJ+GaXBpTWdcqdId1iH/K0Mxov6hxmk1mh5vslKdbCiZHO03fQ
2rWiqZKEZkbAYiKXM+3fSjM0BH7ANy7mlJnC56Oz5LhhW9/2ETtaHX5e8g2sx8nr
e3hA9TLmbwEnEtvtX8b5WkwDFQBSnlCglZV0eVENnOvNYWtmy40mXn6VaOp4MvRp
m55ZtrdCQEUUxIYO0L5P5hS1NJ/njkLiw4Z7NZ+fFYFLkSTP+w/gB5G4QyzOacmf
HhWe+h3pDiqT1lHxiyRw+LtKO4HLhKKEDi4NUdnuaw6waSfB6csyjkL6R8lHIplb
7YWZtDN+RoI/Vj8YGhnPjp4I70QJQZ9awkPgXgHJaaEDVwOuUtvf+k5FKwOaXo32
17T7jGsTI4fDTcb+QWtfcxYewgPQW0IgCSEY1CxKH25s+yVJHdOXZ/xHbq0U/WTW
zS88Qi/wu23s2QARe3SJpqpXkM1H7bZTZkvgdQbw9cAm3PdwAuLKczpGgnkAp8uS
gxBYzytYasgUUQ1KP7PbHEkAo3V1MgllbGIBwYd5wP7ZDaVArfzc+7NzbRqe/Sgi
frbbeLtXa+rAUv7MMs6t05nhnDiVGDAFc7mlg6tkYLNfYhIrlFVlsK2O7jWJYjSW
BDSbnc7me6BDHlruw42AMR9O1T7NfL7mDSWxNjoBfs0la8EamhcEdifmi5/YpNlk
`protect end_protected