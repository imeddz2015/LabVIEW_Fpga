`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 2928 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/9huKRhRMtvnNqb3Z+UU7TahEoHV+T8U3P3ufru7l1O
3DlgtZzb9QxCbOjthp9+wDkjygH0eUfDrEl1ovhZG63YVlySfK0V2PzXssaUK6EF
sr6EKn5/2v7SoAxx2kUz4sFN3K11piPHvVWsrobtCU5zJYZkuFcWx15XtXY6Bbo3
DpVK3DLHyAYGDoCUtcE8LrxpFk5AWdciD3v8VMP2UFzzWNrCt0Z2Um9k9H9Uw1GN
YB9AOZsO+4txnwxLXiwYBZ8aSDchkJ20jbMYMBJMXT5k1QWy93QooA6JYjwqM++L
b6W/ngJn699x8m6L3+gkcZcdfB8PJIlmiloO90QYEzJq+PlPNiWXvx2Afu+EDKRQ
rPmRu+US0DM+p4q1oFd4UlHRZMC30Wn/Ou7fD5MN0j6i3jV0ZO15Bdle6mJJDrCE
CZ6OvUc63sBLQ+JEE2AdoYX0LPs7lJQs0lE7VLs5eZCi6O02OJeU6SRPQXSuUxOE
+mvTJRE06ZI1/6JiEgMzPfh8G4+qFL5XETbj2UT2/x2ioL+wpd4TDdtCjppLHthX
y1eIGf9bBZlvsXJAQcSJGCAm/RzjsU6MO8QjtFf9uXJ8fi3s9KW9630pQIp4WI0R
EBJT/6mnglOuui7/FnpGYLeDrCKXHYouIdap7pTja+0ypaa1OAlQc0kiX3FzWlfz
qK80lWNw64t9AbNOCjvpyMhXOhC2D+oGxkeJw/fyfV1vg6zLTDHd0s7SX5o05tCe
CW4TXQa7iDgzpM2kp7F9jynfvQ52feXvF+dMq15KMWBIxyMC83qpY1HA6DDozdfs
fU3R8tGuh8fOkc2tq7GY4N4eTgAYqyaeRKP9E033g7iPtOwfLC4j7oTqCs2m2oAI
n4Ewt0GnwPYUhn2KrKtnmdrm0YZRQF4hWJBZrTQm2s2PA9PLuRH6mxvm/78gXati
D9rXdEnTDuLRAWvWuoBaNsb3rqKjVAbGI/i1Ut6SoWpUHRhxPLMFSlD54BWSqUoR
KZyU88qcwLd+5LDJHIKm/ZLrnPewy2L4QnIhyj0W4yrPIAoUd6hGbxOC6se3dsMC
GkJuy8XqyYhgGwvebMjDVc9kVgBzAJKFC+LBiyUB9lxhePOExejb/N/YKZe6K4ye
8kmR1vNuzzMLT94YCsvsGwedwsrEp/cO9z00/yHukisVXiW+FZ24UAFaTg59tML1
7+oQ1+m0exT31RoQ4+zLmFOtmq1TbNtH4smRA4Wpu3c/OixkwpWEGR5UblffRHwR
uleXauz8MAqxVL4EqDlwY4RXQX78wG4jtUcJLwlCwajuIQUYXhzPun3oskDOEFAh
xJYMSa/4HlSZoWnWJRlmwGt1C5Mu7HX8+crkkinXAsDbDperhYWMB3mlocsg5r9k
3O1BE2bdElnraZ8ojwtiANjK86a38o41UjAvNrQ9vuLkhRMIB/vXS8NbEoXSJP23
Y2HrS9HNQVLew7EfPMNKy437NkB+SFh48YWWrLqmRh9k/U6lTzrK2xR34nl0FyMj
4kkH5abMsBL75+YWQCFlMDjnn22Q2h6OpAhDpXsJeLLfFCciAyvNeDKkm+91uhWC
ZK5AF7YBNUpUgQBazNLf+qmpQYuDR31xetT1varGcM88ID+O0qQlN3JMSZSd11Td
Qq4yeUeeLMMk3e14UcLZbcfFnZePGA3I9x/HgkhIpfSpfe68y1AcUI+DR9w17sfz
Yu97H1FrdZIvtP/Jca1E61cpsHNnkm4vJOR92J9KQhbRG0cK+0EhjUNqPJ3sLx3N
2H9phJAIfBXkMtPJBaUNf43/gdw0q/jVG+jYg45+XUEly2PPaTpyO6FCuEO0TAh0
RebUkiAjz/F520QLJB7erQKyz3nPL2DibYUtU2i/VTZ6tCwXyzioUlXQMI4Tb7Hg
yTTMsTT8+eWtB0SeZcDsN4GxM9YMyBzlKoH3uNkJ4s3/OyFJ8Q0VvmzoIWCIQC2l
uj9kOTsZ1qiO5S/uWF/+AyR82Vt/ar4Zy3afi6pJeZInzEUzHn3gGQNmrdhIjmxr
ytESRHT33ys+9b8npC9NR8v66Q3dNVGyW/PPMt/WL3h+od3CJe388n5YV7BwDoZ+
FvPgCLDs93/lw6YOIblNQfBgSEoSSaHc+CJC0juivYkGnLNRrqjEp57ASnOmvtFo
OQWJb+zaWV+EiVZsrb5e1pNYezRKQH6T2PZRI82I0+VElG29tB1F2P8j/j1QdAZp
9bPOBv/sYLFZuEQcgRCARCPaOqSctu+PliMfuVNg4fMhgSiUubSTdJQ2acnvO1dl
FuotL1IMMuC5V7ICSXn5gyAb6Ze8FUlDja1QXjKQZWiT0a56zplPjLF6uKltZXeO
tCjb5xHI+w1GB8XtmGtcaoHJTXsRPURoCgo7T+6YGdp0/qT9ebv9JRu9dp6n2/28
fgxXRPkcIHxRhwDPwWxsrxr5YQOqD9o79jdU1QPddpsEdpNj4Sn5ZpKvX3qTyaVW
RGmrV13gH8DX3kArjV8D8KrxSxEfQ0vBlaObrig6mxO40Fy+g4w7HxO2H3tpXOII
e45QX5zhUf06lc6p1nq2pq7C85ZrjFAttoQayThfUh+DJn3fwb7xeqdkdaVqBWHS
+5LTbqbZ/SWnDPqYSSEsPbFHvrDNVu57OWzgteIGIvBVIF+meWHjg8fK4enL/SeX
NFoKvNJGgPuD7kLa/nlb4ejNnudb9mbtgxAhIA7pgn5aev9Tw48gP/qHijjnm49M
kSKHokfigFFe+X7ScpI4LZn/y1Nr/2STmOt/vKR2aTRjTDgLi6tb5FBhbXbNgTuw
03YDuJh9hacliokrGfsAXeohQnL7lnXYPjC8DoqR6rSAvNU7KuglvpKW54+yu1Jc
JUSxRs3nUNf3lTvqhPJW6CKYAsSTblOC2AJ5FKWhhGL7Ua3YsJwY5aVfmPG+Xn1t
iPkGtL8SdwNVLpcfKvxAGiQtDJHr/rZufANl87lsokqfkziDDE6pLtg41eHC8DNM
/XvoX89fxMzQo2L04Sir3+HyKPEG9mXJKRY3btmp+T0gxUUpe2ofsQOHnmdnWXLB
o0VGP1928YBLYPEDhh6RaceX465QF9+EiluU1UGCYrUwXkuvhBlbDz/2PTaj4cp0
ORBqj08V7DI8eaPn7Yzq/HgdeyCEpI3CnXGm2+gnPV9VUo7i7xEaGEwVOWK0Xv3M
XK5x9SuKpoquQz094CSedOm4FhweJPupXCktYr9td0YswpNup1/ZpsgGeem1BAAi
2mex+XwTYpdnnHxBHZLsbkBbd3aMOt+egqbE+t59d0UrBr/UzDox0Xte/YXFFGFr
pgU88xPXWKwNuX2yZ1Qep5MBlxdwJVwX1HveYIfeRAhKIJ+FpBOHKvrm7nnEipW6
JFO5eyiKawtp8t4XQJ681MlQiY5xbCIBEmvxa7J6h3GRoaflRRlqjaNB1v3LqEen
KbepF4q8L5bFQkPduQGFQA/usFkMaxtG1n4mtrKeNEKnvStiLzumqEBZhumcEUFA
A5KvHUZEV8ZceGSdxw7bh1T8OhhkdbhZiJVfQZxcbhVADqZBm2ubCiFbLCcD7vgD
k4Gyi6mOt46ESo4NlObhYfKZrUSh4SpyAp2ItiV7NkK/ZKIe1Uv8K8spmwB1KHZL
KNjV7SH9nDtrn2ToXh7MWFzgQGhhP5rzT3q6wF3u7XbR8NrSo7n7gZsaBXf/VFm1
sExk+yLLfxHGqqQV5G/K2YOaqWfryT0lKkXIlE83StERgxScQX0/36CHCC2XCyIE
4Yq5tVuS7etBw8m/PPmpYlsLIcQ9cR0Kc5MkDUzzjT3T+HSIgSSQ5e3CXXNQdSAO
DMVpBPsyji6HrnAXrJk8vZLSM1ztatKpTTEYhyZxDkNPH/gBBbJqLB6QO80du+Gn
`protect end_protected