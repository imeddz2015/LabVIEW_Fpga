`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 10096 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/59UwEX+aE7FohaWu0/8IpTj7mav863zUNIsgIH2BWb
Abd9opeuBjbGF/waQMI2vMJTwD1ie1YueHc3nSNpEh4OXp8P5ybZFY89uyGz3ztU
W1EsuUnchJoQgbHZ/sLbgtGRgsrAFn+ZoIeGN1d6RAF2wAESJmYP8zw+p00RvjZ5
pBGEHX7wooDexzkaqKS5G1wYbGesBHbRKJMhACyYQGQxL6V68zlC2Ypa1f9r8MuO
ieXyxTh6baTZBj+Nfj5cuJ22x1cq2jGnTb1irg1pkbworSZUlUc+lsLpn6t7Owme
NDmWIrt9DSbu56RJdBJH1qDFGvtLo9whISuCJv2KIFdBrNuvOh5U16dodQZ+Iw0h
WHV+Umu/fyIpNJlvSX2qnVa7UyocULeIvAOpQS1oGq3y4idF30Bs7sODCYCqCOLB
DKfySuKJlBAOOvbc9KEwS/FPmFmOewXbbzI3uq9duTvHuEI2eD9PRp3Uqi5kFuph
71aTYf9+elkYYAbFyeFPkhTVuQijWqDh+67o6WSzTf7wnSK14VMoNN+az0oZ95ok
PrA8SrnCkFQy6MalLcQKRu0TVK+j2YPkioEPX/B+J0hjofh/5vmwqTSwyeIbOwzC
9C3eOsFvUHFVmReEiN5vrD30QZqtpz3Nz1q108+QJQGaGVbxXdKT+m8vhGxI6Z10
N0ULZ0fJ5dBEwxgtYbEPHWaHNhxYnOKJrkF3wIw5xWLXZRoXTMbBvNRFIPCp7age
x8zsfPuIAqFqdGvQ4corUHl8b70fxKQb/07++AL2P+eAlrZEeb4gy7uV3gPCociG
im9T2YLf4jRqAsu5pJgwh5PqdTieV1r135CtDzkdSjEmqMt3lDskjNOxi6vlODbG
nckUx7ptAPhgrkVMZNx/2kvtPRREa4vBkM6NFRwsJSuqfic9baO/erKTZmweQyf6
b9aE5wSjum0siZOEhASzxm3t6DDnDdbCpxqSDxV+MkeoGoGzJd3dlZiX6WJzRBgW
XQFc9HktfF6Q6mU8/s9x1kTd3XgZsIw/DvEDrpQ2LZwoqI2eohF42ok+TlEHrQnA
yJ2MiyFKDYaagcp9+wPMYWdfcYi6IIxY7Dpwk8BHJC6Vj63ZNG5emB4noZvO1vLR
ED552+Q0PHxrDiasDupI9yDU7KFeOVJeKBblYSnyPN9R8+tKu6bJGti++N/fK21a
XpXcNnuu76MPvwQETLENVKahJW3I6GWXfUtPt1SVbZVdxxIEJGR7JHEOWEhNK+ti
ZUsE5RvyIpvZTAjJuIcKENA/gvFiGuUV1/SMivFpGOXN7TMad1ORyJLOjDsxcVMG
G4lsgJhq5NOPvFxEf6EeGJnod/+EPx7t2FGdWTI85NBKPX0h/BSePc/HJ4pu23zL
htHHndIjuFdcputcMkHgb3J2kvLUDlpCutsDqMm/XpBwMkXo+MSk7gGwx++Yl0vc
qi8aCMkYKuBV5TlQzkyVr6VSouwBFG2gdHMJUm0rQVcc4hzSwMa3G/WRFkKFe19x
gX+6eI2yodws5xdRCJygyo7mwQIZHVe1NgXwMPwlU81g/XhtPaA8/XQ8s/QkPNiC
pNWFlebtoT7GYoyp+mT6LHwfoHE8FOIFF4P269/9cZDgfYOipHnMJ1CmDNjLYSYx
+qNB8YtnDr0Xp+4TGdD2sYI+NfBnpmRKxm11dIjewwyOU2o5Wntnte2QrAp8Ymkt
oKSaTfb5fbRwb4jDrIOGxCXrPpUbLhzhBKIlWXiH+APYAcSYXM8+BnFCJks0DhLZ
8TTT0c420oCXQIP8W2NE24i5EahcDK9185HDCg0x8i379ad4sztZD4+4n4zPbHlJ
YZZRFkx3VwPTNTUARScXCntSPaKORYwVB2goL9QXRCkeFSjGp4aeGgdZZGJd61AD
F12Mz31RtnVS/drOFfNhP96RQDnMcBcJR7q5GUCYPlAvp15BnncS+M3xEuGDabHn
yxLTa1YhvgLyyR1Z/TPsyZ6gZitNW289f8Kzo8BVhSpfZ+RthtWYMPhA6NM+FTQV
3dAx2leUI4nqngf1v+UF5kbXSlfzyVw3IyoV9DQiePgHeB/GZjv06jcYrSOywzsy
sc0n7OJYHnU9B6dKIYOQUy1G5+dpugQIsqT75VZV8SsqTOT8hwfv9SR4MBop91k9
JHIYKMqv1oihInSlI/MZVR37XbQLuEC1ZD6CAcuxhLRxhbFF+sqlwdwMb0pORNvj
C5f5N/JMCfJ5/4lH0NuHAz0nDAPf6e3mk8YkZlR4liXSdX9RKfLCK9JaUrcXiWCK
7cNU9FxG3Eb6OgotmMucD2dlpog9vu6JRKMb/6yKiYOboxLTK752YkTMPA8th+WI
wIM/602cgIVp/hrEJTKrqh05SD+xi3gy05T35Ep/0mVDc0IgIlpRmZUwDKS2YHii
pMrlz6/3/k9QuvjRajfb6uy5BGPMriLhYxgmqFPAjzrdAGS21DmICyUIYcjT9ptW
Yz3exMs3MW54oJ16/FQZzA3vq9KN17KAYi2MncIu65IvUw/bPQl/sRTdLwUOyt0P
O+PYPSXaoovzPdJtlyQK+caa360t5FU3sAxJ3DuchdxfoS8CvrcvnqYwCl2YzKOO
NY0uh3mPGweMKm5knt3c+2pXTFGkDWCxAakw/pVXxNMqvMS+UfmOi8eKUsSPkECK
Dw49yo2hdlpNFE01SWrwH6OvFaWgeUo56Uznns6fsfVTIpJ7o7w1Cs6GQO9/ZMvn
AeEy7SZgm5Nbxt8k55P6LkcwvZTVLLBtdSoYNidZwpyMY5dJHBq0yX0jjWA0oNtH
caxVFvmSV3XX06YpZ78Y7k9mV/YTyp8exdbi30dFhD0Y72LU19Gg9ENzw6fY7TTa
LtZkg+Bj3ehiBsw3t7/XDilTIQgA2D9bciyGiCn7SNFq2fH5h4K+QrC7zXCLDanQ
InklTd/zRQqM4IG5l/CTk/nVL9qi9e/zt/QYJFINM0kATVE9EgPrSQYQHAeS6Sod
LQG+tUpPdCiCBtgNzXm/prtL0HMAJ+wTw5os/muKEpsOKitzAiNFO56fOPPWnVpj
mGYirdG9TLYtwMt9VHKtMGtpKZEPYL8ktNiWw7yYxQsoh823bgmVmUbpwz87WcaD
VmBPUyFDFkUXZ7HmwEMd5FlqeZYxK12fmpoTy6x3ayJnC1llYaSIzcU4UZLHOVAi
sHC5/QKgIVtgtxneq6EvLuqgl0hdybDHbMDjaDd1AMhUb9kYUydkQkRBwjNk3t/c
WSfKZ/z/EY2UXE3J+jeWkNb0b5/3vOTrhYT1Tg1XT+DHupyQvnMyMH3OR3BZLuqt
SO6qm4JwCbWR9BBY6e4jiexcxi/FcZGQMiqFqDRNCxPp/Xa0MiyA8+9CnxEBxt0i
d051PqNgHXdiGbrcIub23BM4VkCzKQ7TaMxZ7OALxRDf400+pWD5bYuvkm5D7XA5
2OKC9+kuFPzuTUo875nvffFTrHMzhg3mSutU0q1WRs4vzUgl5LqraEmdXyfeBDiR
GMePULIZEYgyMz0L4bCcRO8YilDd2QnMawi/Ui/jt8j7nMltP4VD3/w8EVzW6eKq
A1MXla0q29WtnncoPIcFfFW64v3hXRWtdhSXLGU21GKOtD8Xl1wsT/BYYSXFTHN7
0jUBZyIq7XzByOyKhucS/3E3DhsFgA0kDH3ov0iOcizoyU3JdKN6BiG/WNJxbMAD
9JGpqQC64+OaX5iuOqrcDQPZDieJ2VrjeTauG7MNn3lYJWOagbGXqOmiD/GAdfet
1PFmg7IsAoe/JaoFA4x0PdJokA+1RI6KKapwVAlF8CR+VvGASncjv7HjIjgifmpM
eAx9LyriqVuJhkEWA6kr2e3VaKpV3LrTooLd8UT7kX3FVhoTL42jII6fpdcUhTw2
kthwe+ky4VdOuBeH/QQLPPovtGxd34GGnzPj4Yj0nE95znIod0U/NaYB+pY8X62z
l8LqjxH1sCtheWXgXaVvh99UDiI4M2yA7eOvENlUl2hbFxKqu2C3NcSPY7GZHo//
teViP8uXvAI7DORXpghNDKfPypHYcSoYm6KvbLwVBKTfEUw/9wFKwV+syxB8rZSJ
bY1UT3Dt7bamy/cXDHmW/NbA7Syyu8ud3SopQAk8NGQtrDL5XTxWebynNpm4vYWo
z2LYq6730/voqi7vLHNr7evBxOtfVQNjII5Lz0Q4cXrGWPl5gvr/JsWZOTU/sFwz
u4fgbL+ebuY2rSFjsfiUJOOIFZJ5dZ5IpvR6xtlsd9v92ncTSIy1HfqcYStWCSM6
ZhNDh1QTZtk715UJoAhhXauL3NVKop2P1XxKXSCwXZCJ9kg/WIhPJtwAvVZ77jVq
l8AOnZsg/hW3iBv0bbRjpeUSA6cMuKVFTI//4kUiBd6oZIKttKmFVrZSgwqRAuyb
BdZv978F3ZS1DRTIINpbbcX5DgT2vQ5vnh33flcG7pJqFa42qi27gaSWNvhlqHq3
jfSRtwdNwXjD4lhP0tRrEYzrxUPVyXbqzMFDwLUFZD2WcQYHFDo4wr+AL1CYdN1O
d+xXjUSjlMPHR2UXNrCsTvH75anYInzr/P2e707LrH3gofdDEVaZCvKbSoii4fFM
s1qBXJRwYzGZa0dz2TumHZZ9QIjfI4GpFYinAO3hHKmCJn+5Xq/VKlSM6ZbrVYZI
5IlUPtau7Fc+eozcgDMP3c4MqNhvt2+rgCZAGHav0o9PEDLR61b0FOb6iXcowHKH
69eWCAnlI2ocvF2/7a6Eou/9utZlngUZWQMybwJv+1QI2BTXEqFQgNCPndSB6Zav
0WxRSXPoRK6A/gTtC+Xn0v1XRkouON0nZpUW9kS9aR83wnoM+AqPzF0fESjbuSEN
lc9eI1NayU4OxuuGurm1sIADzhnktXDehXahNlNyha4MtrnppJNJz/Wp2agNBMn1
JvgL3F1J2A7dOmzFviJ/4CIYxCFJXWumeslTn51rdidL281/SjFcRRfOr1e1pu8A
620SIbqjiLHzvalYKKxc7b2d64gaEWdsmLnPaBockG3KKyLpG+Ma3Wv52X56ZFpl
HC895pvi5rIdULdMw9l4CTlTvDzH95xvnFUdL6KWK5ZDQEiddckgbtagoc7K7+FT
UXBwnvUEk9BB/MC3V6Wjv544kaPrUZb0rWyD4F7EIFxma6bC591yeVExf+Xq1nr/
MecjRTc3vh0uzmUzlDTCgQ0wIsv8rWsKkm9IoZpNtOUp8SKFuk3GKoVXDEU5PG82
v+fpS7R4uGla0ay0E8l6R/eTmxkkmJjzwonYBe+8gJ22FvY2OUW0E4StISSQX0Xo
tstPfZ2voLk/9mX0MNAesZ+4cthERJ3/GLL+ImYfiPgyKeTRG1xhOCfZ0Qfs4pJ7
6T3r3FPazwhC+4ArQUP0Fdos9/BiEc57CfI0HzW4861EGlSJwpXU2zNZJ6WOP4uj
oZ/Bym8jqJDYmwV8H84XNavEuXuRA3FnIi7RG/nSkS5d2H9jgAyptQxuhXrl1DcF
0ZMyIyrFb5oRPA7BoG6GDc8a04C3k9Y7U4M/WwSMEeyvErO1rMFB77D9oGAefbWD
Ga1scZIWpclXguxa7qHiqPTkjdrbtzAycnihF6+uVOjrIRBUkZvuhcBRUUncw0gv
X0TJjxecHPGdu6jIqCm4RNKw5fARZj1xbYYE6LU0H2mg5SkuWNJQPYhJy1x1IWMG
44WjqgmAUCvK1KgtOQ4JkKluY67vJzpHmjr5jsPER43jOBZAKOZOcjIk40UwzsMJ
AuJJW2z0N1xWKy+lqr8JZUwUZiqIUEZBg9VhXomS7+4mVjGU3Sy/mRFuo2UnAae5
WRuHyW2vDFFUvgYyEH2T+M+q7jM/+Ay6yDLkMwE9i/1yYBJ621frfoUwLirlA6QD
cWjiToplxYjV+Zahuxrj+fP4Q2SuTkWybR+yu+YP8Tiw2muBzMn5B3/3PV7s7eg6
Wjc0dpzuPuRodR/htsn3hJOXxUdqQ0Rw3bt9w/VvW5493dQWA5+LKrdvTdMcFCVM
t1jLG5MaNo9DEY6OBgTWd0uBMARJQe8NuKKIG5eQEDZX3XMFTpUwD72w+dyXPRMW
fOXZ7pxLFt/hCxo/gvLN+1ha+ADGEDezNSvmSk+UP7/Uh7DOjOvS1PzqWpD5dlm0
sTE+i4sP5WhIZ6fT5SptTZEeg7Q1LaUp+BRk6KfVc9rFIIKlQZHSaKe7e8c/zYRr
LEFlLioKpj1+moFRRgS/oWDbPN+bVhU8WtgdQsXwNhDauKKX4Dd3tUNV2wLzU3dK
SQ6XdC3tXoe5EfzzLmQH5Q5hoIchSX4wr2st2UCM+51FLFT+oFU0PkHpRmxrlcwh
4PkcUbCsaC+RnoWwCvWpIsOvh/KZcI3MJvK8voLQtZhxzRVo8dVIgOB4vcU/XWa0
R+d4F6cft+/2A7RWNeGBPelXX5Cc7XKAYMIdWEHd2sT0z0gNlBrZRyXDsAKDXzmV
kiULYMiMX3UZRnjXN0p7bQGDJEK2vrcthbwtkT0LoOqOWUNUpLVKe6ZRhKT9piHX
090p2MLA4j2wGoOA/8rqq9oQUEPAQ+cj/paKmW+EC99sszNl306aU9q3CT6nysXg
6s/tn1WazKANvODa/hbaDLOssuSmRmIWEVh/2peUTpf3iee88r480vWU6oXoZSfw
FLjB2wY8JuDNUfOCs07S2YqEKu50/Ug3yRHESi1Wh6JL4GRktcypROAsvCy664TD
NzrOhtHQT9ppL1pr6opexoON5Ikv9BI4ylb8xI/xNv1aK3ZG6uEraKoc1v+/F4uu
DwKZ1Yg4LaGBeUACGfVgxudhbGbuIoKxM5PDmmw4GS+/P8CGYDbiwByV0XxnaIr/
99TVCA5hO91q1vP3wXRpiuX8VxT+Ug3AvhGuTMBQgV0wMFvyr5ZrFqo73nc7BEmF
ybJvjyMliavlvaKSqn+CrIVrgOxxzNG6GNzzPjmH391oGZJHFaRr6649ZHpG0QZ2
iCzE8Zmrlks5aI+kD/xqkCZxcZ9E5vFBHKKrV2p8t+BfxOT30sQsaekYG3yHJGvI
K3JcA6w8CVs+os9/FW3ss86oaWRbgBsoRY2KBc5iFjenG3EDaaGmWpnYDMp2N193
pOr/ys5zXqstngODsaSQckwP2nRFAJ1CfpYKTXHr1EniLxui6jg5kEPAH3bxu639
I2sMZEKHvwnXLEzo4OBlu02sQNGooJAcKmJJ0Axjhv5ox4hSBnBI9W2OCoiGQhs7
y4FfWW98XXLfr+gvdRvcoIcmqzqjBBnaK116QFSIWKQ2295h2GXUTyfewEsdQphp
HzVmY+1Pc/4soIWFrri/d1Ioby6kQhc/OceSHZKD3LJRaqfHGzxwI33N9mpgpKNw
aQeh1+Y6gR92bFXWK3rfmzUz3JrBJ0RN/ZLL3+5AxPAjZ4TRDRYM3yMR2k5APBMn
2s5s6tDgONL+k7dA0kEZ99C4kEKlO0zOck/z4nllR3dB2CSCz7RQlM9OzCz+vt6d
SvhLGfGrKucDJBCYR/ry94zJRk4+11PMT2CAb6kqmmElvfzz0JNa8qohFw35cpaB
qIKzI4Uhnnx0Jt5HVjkwmkarvzJzlKBOjXElp4qcuVq3ISRJuPus7332Xy9BPoT8
mEnA42kjz5Cu6UtgP7BqsizDSRhP0AfE408KeE2wY0co1xtsNkyXCC5bVpXhB3II
ETrOLURzMd4dzrMmuV2vPPRzJws6QVcbJcjea+57j61RoTDzsqH4jCIqbAxWmKZA
5vJDyneCoApD5ibGSJH3pKKx9169DdHLYENSQfs1OzgzYx7V7h5GBbYaREWdVPxV
OCNIH5ckVADDXSn2GWguDYdnAxfZlpW8NvcC2oDYlzNgUk9GGTc6DG8xeuMefutk
RTdSj4iF/fRTp1VWKuDrv7FqEvI7P5g/QQMhaVdefsx7IV5+2DIk56BMYrmyq9Db
3632HEIQyMrWb4MRMoL7F9pOy62hKIJRNis3u8qtupoOJmBS4SSmycnHnfY6C1kL
+C/TnaEEB0KsgJBRYzuTukN630EvIOMfofbfUZp4ciDIYtHlH4gM0om3tuyznoLj
SBycWEEuFxy5IyHTMwdr89BpprlsaDxO72HBJGAWAW9+Usuto7V6CI0JEbKB1WM7
xcCGuQqYA7jflvMWxJQmLPwT0KzbjpgJ3bnPs9K8VxjXUWq0Hzeqv4RozK0Jye7e
hQtD7+79biWPA8fB8Y9q1KD2fla8uR92/Q1Cv43MPMFR3h6d/kHNdQr5BhDECT07
CwLHDffkzoqTcin80euYuozzhBFVL8IOmvqi8dwwHLmGOq70MjoZOAEJEe+iTqer
GU4xBXSbdSwLYevNdTz615a3R7z6b4gHQXlj7/Bk+bMOOozNAefpy1O3AFp2T1+I
0XTwilqTto7Ura+8Kw07sJ9bXJkaYxnO8z0XGQQhR3r/fogb4Z0iazXsEcE9/ANM
EOeJu8L9riDEkHH7FHFRFO+y7sp2zzwyrwvJs/GgwlxyZL23foT0StJEX5YJJ4Nl
5mGKTqfXORq9JU2fQl5uCvdOrAGYSx4h6XfWKUf+r533uW9Xkw+nfidB54gdjKBq
gOnVAzeaX+6YWRRW/BGRvKuCGyJqfWwqZ+HcPbopqUyEB808EG4x7OZbCWOV60ij
XpdIkZURRAOhmV5Od67utvF5MPCHHaxsdQ/GzDB6bpZH7aWgENCbGYrvlASY1AV5
R+JSBfMcswd/T5hMTXrnqWG2ZdV2Ra2ocHwrbrfA1eaiB1Px3myTCt1GX4lgAbXN
6UX6gcbQGJcLDg7F4t+rdxB1xIGUpA6ZdxikcbnQGkcLAqZHKRVoQbJ6mFVQeKai
jDI+NDgfHE41P4Zz99cwBBVhI2+OOyUE5qcWiP7QW0JtfSJAB4DYDDvnPuhYFoqN
mt081N1la43lXjq56CCA0xx9xJQ/x4ua44q0/xfKRXZnbK6hxRhajOaH/cGQiOFb
OEz0qku2ltqQm83uTRYdmuIfueZhjFnM12+7hP717rsGskIEfXjKPFf0y6aTYS28
rsa8TqKQEcp59oZpkpxdWpaufY70gYjUbLunXJwifbQNvW5JVm0ItWCuO04U7edT
di2S+QlQIumxgorob+rZ/S41OcL+cCsnE36Ydx4f74EPT6iLC4sXK7xFEVnIMsdz
Ex9sHhhyGIUhQ8FdYu6+JyoPR90sITCw04KubhQY0KOr5kjZS0rC266rkfUSZGdt
yvFX5s1NqqgUVjQ64URQp95MtO/whD9U9JxLoS/zdNnxz0fqU3cf8draB1QQcWpt
fPserQBEPSwBL0mY2T+9pBIufeblmbpEP0kuyeVekB+SuokQZ97DGDELT5K5W+i4
0vOJHEwRXBAxkWWPMPnZ4j8vvCOSd7agzyAQDgavp2SEG5h//mh9DqtRy3BE9d8r
4UTr3V8K3SYf60/i2v0WFeaveR/Tq4XYN93eUigXuJuVm7nQr8lICA+uMcwqMMhx
cwOqOP5yGcGHISZQrjQ3HZVglP6WSgQMXmTUocFq+QbjhQz1GCM0tTRJUlm1q9IP
Kaq6KfMJs6scvUWHJx4/2ODxqTb9GJSqn2YUGBfis8JR2zf3/wYFeoW/rfv9Xj5x
eECImna5Ampd/qU22/u1ZAF9+KPf1CBU1U5l/++0fZxqE+LvUsNn1JMm+Mcr8iUe
8IN/p9c5Onl71v9GFheViODVvKGvwMPWP+8edYpgEqzsmD2KYK+wjj7N30N3GE9D
3WPfwBma5+ABvcgKisv3Qsbw978qtsVPXAFFE8f27HajHot83zeBo+gzjEn18InI
ngHMB0rBrYyS45wvVKe898BwALs8R5CD/CeUMY1E1K75+NawqXn95Jj13gg93DBE
3wr+9drvfNfgCT242uodqQo5VP0VQvG/pQjYaTsw7F7z3KnS3MR66YKwlPkS5QDx
o2M7msITCGqXQnyIj0Tisq1InN7GiBmzwfC05DSgqkHmANXyeDQuVUT659CXEARm
7ye0oAOZdjCCrmTYDmdXe7x/IWPmaqbUmG+U0lXvPw3Ji44IBmU0Kv/FZDCRXxSc
qYyVRcwa6+O5+s+08MzSGDgazwBBO6CSZv40xNkGQpkZEr+cnZDpBEds/XsmaVUU
QghmjaMGsWfmzbDwFRM2M+qBa2p1F8O+Vmzfe6+p/cj3AOfD0RN2oLmML8+Y7kwV
BY2KBKY51fjvehWRX/LxTj1Vw82tK0jdXYnbgifygdDeMdCDiNs9KuULLUgqA7BU
mMbnccJpYYa07YLxIHQvAvEERUhjoDO5SZ1EciwWz2NQj5cU/9gN/P80iXebTdlx
szt8EwRKslampN3WyarfPTDaWsGJ2kCANVoSixoQtc0roLxFMJVtZCWvSxHZ5oCG
Y5l5HPJwGlVvKMqd1vLy+OEx8p/wWgburSf9V4oX3skHBurwQBvw4rN49nG44lYh
LlsNCVTqaYr3bsFfoJGKNWEr/C5wm5aCInWauSR5Of3mvGSMpdLlefhLMDC1Eyj5
N2KFQ94Ak8iqLCjElguQAAjL61o3Ez4kfSgLRS2rbI4D5nCKfASBg2HIavtt1Jkr
+8fh1aMxoZlxWR5QN2ImgbUW74W0hMXZ1fOKti0ConlX2O52VfoBAWe9Ym/K+xb9
v3G9sUXTNGKgSE4aJ8m6EG8WXmBhXUtfSAnD9PRI1hYSxkn2N8mIBxDm9kFg15uH
Uf6lN49WLR4ibodY6wio+bJnJuv8/7QWFk3zXEHPX8kU/6I247Mlv4PRKF30CPJb
EHc1bEabfA1LooSWhdRCYhujGP1JzCuGi/6lknVqB/2LIcGMgal5g1hIu/tWdGi4
Z8XmjLPiiMHQjHkGtSutQXt/GoOY1yreYUb2H3uuy09F8RtZyIdSmwZl94IXGCSv
PQB2kU2paLKrlYbCoPt7FxA1UVxwVqMDOgpGewQFWC1JMWteby1M/jX8JQSVdoMm
5SG+00bVZ9wRqXFGDZxpl31pP4/DbdJTGPZ5xbF5xTXlzEEKNKOejpjITAQ5wuaU
9NqMx7gqwOx8qqdW0H4i0OSvdkc3ub15NY1s8e6alx+24reWX0PAZYLKzoEvjz6Y
Svc2dec5J7nTGgiCWqANbKQa/mjF4lOSsb+4x+CcovM6VLvm4aR2LlMtfIecsrVB
KpdciA7pQe+t1XXaQp2Ec8EjWPmDAi1SGZrVvzAHC1OUbDfJPp2SPb01T5X/cP6Q
tu/CahliFvngKBJ0Y8+QakaTFE9Du13GZrpfYP4eeQwr2L1zPaky3nISKm4nR61u
taqqVN0FmCj3NJF0MkbE08c0QPAHH0p1Q9tRTfSgXjpx6AHkLoY3N9opzX0cZ/rU
O63MZ7LDSn1DMunhnk5gxOdBhsbztsl1WJ8M9J6uSJ/ohsx7BYK9R2ncYo9N5Eqg
dmbVDaYoz30QNrXWjWzzaN7gvGjV8WqP24Ltbej/aVHWyXPNE/IsDBuUKrV9YvMq
px1JtZNXK+YbsOEYj5vtYzT7C3AVyUcYLxCATlB7ozzZ9ns3jav28w2+oAAqIsbq
pXtDxbpX6C0cdnOemAyd9IORKqUA1MtY3/C5ckuWYoAvM2OC4ox/kku7TBZW7yzD
DwjWbn53M7m4KyfHglh1WLRU81/4SxC9esTdP1Dz0+0vDIH6UgpjwP/TKAei8fP9
/xTG22AcElJQ//LwSHirEA6nNNGFbY5GstQSxrmkV/RWQ1vFHaFRbz2IQJwxuYQj
NrEzjM0wAVL7eAd3Rc6FjvRPf7zr7gfah+ytkIK2NhaE109olNXeQ5iJbqhKdOyW
FxLrV9XQspwXxNFJG9MwAJMfBSrDD+g6w3pTCV8kWhQqBa1HZ5c+Ljx6vEp1dxXC
5uPJ/uf1Hj7htdog2YUAEgh2FfudtVlk/FCjMhDYiricI/+tXa+HRPZ/puP9zqV5
qJY0tlwaJY4bhsyIMiOdUX56tyPkJUBr9fsjPwKm9U9/wHmpl9kjdv10CGMCQraz
HgFWFcsO9XZMorSpZw4lUsVFeMpix42f+WGLrQan+qE12z7Nk+BZUt7tlT9fLixU
vkij+jB05yYrRelp8rBkIlQGHscwnbdFcz4DixG2sYVynTmGsBGwwU+WUv9/PMDL
H5ocDQv8TE0RVfS+jkTUN1IldMaCRlvsd+DXb56aEIpI+/vz7D+ZF8jY6PsOLg6O
q1AlEi8nLhNAKpQ6RPbyyQCI1fa7jWBVkRpt0dfDDJjIMMZycIS8qp18zJ5T22zG
pudtGD40cxMlT5ty+iF3A8/4ow6inLN5a4ydjadzn2rge3kXNVyPoB2RcubspWLv
HZduuNMl/1VeKpwoLse5ACMO9q9lW50Izm6fsXZBGaz13o9pWm6RPP+xnmLgGKyQ
YVJJ1KEDUw+ThVMu4TtTnfDPrj/5lHaEiePydXpysyVzaS6jQcMdPKKlKu91+XbX
FbDNC2u/Co8S7qLEogRtVC+hw2ueH+MfG1NQz83wjJ7BvsJCYkVwuq6DejDLgwQn
ajvXzvyDVX337E8lVELeYn5zwuBqL4UmYFiYAPO4oxxE91D7PPomz+U7c2Wy+OUz
+HWjeiklH0QX160ljoXQ4VjPWy/4UWEVs9QaHI9q1vcEijprwQe1MtIN0+1h9rlI
5hD/kAvqlZ4LKqsPshvQraMlRF+N0N6gba1C3WYissI5o07dsIDqagjiqrY452FH
a+zAuuFuYS/xoH5A1BvphoBpC3tqtrVPea87ytJsyiduWr/32VwzXna4hiJttX0p
t03/7cdMgklMZ8eBGaaxYkjTp/UfI3NUBkLUC5UtiZn3hdGmHZWP5w15pszsHMXg
icoAE6n/4G2vFcVIrLkRUrP8HZ4GBJKUvdN8x7zYJRrgNBzvXmRp3qtx/W83tsfq
YirmZGKM2GcPPXl8vkc+2UkXH75I+IMMkaqsiqhhc7DLeM5rnDFa8w7v9HJNuhBW
A1DtWSuobR/ikPEpIK0Kh0wiAPE0BUEI0RLmENFn+POeGoU8/tdLnaU8qyDgWm/r
bNfMzEivmndEgSADn0p0mBKgAGnaoMMeI0NYTyor8jv/YiuRUxluD894yOAUrcb+
Me28KtVOJKnTUsi2L6yP4oaMOJ4NYS6xJHXAO4l58anJqyIedtlETwxIKuzezi7K
P9bt+ghBeJR2Pm0RQuKwNNl0DSjitMT4mxWNYj84/AB9TvWKAneqyp6+GREhkRU3
jwNJ2GBUV/GILiiNDG+UXYxyrukWo0AMPZTTFpOg1E64VokmBFnQ91BDkvuGkMg8
btvwFlzQ0GZWTK3AQI8ePxs14y6IFz6OPsaINTB+ts3FwXmuptm9iLj9hh8wqa4I
p+b3kh3FgyiHxYfuXeLN6bDRzWu+rLBd+vrYcsbewio6lFYl82ycEPCr8/zCz4ra
PKoS+JUlECwzxgf7+qIyFcUB1pU+wu3VXjtaKNlGiQvJGgVqjmwQnDh8f9qRfF2m
wgS5jkkmJBvQfRKbEzyu4w==
`protect end_protected