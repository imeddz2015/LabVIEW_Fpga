`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 15616 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/9huKRhRMtvnNqb3Z+UU7TahEoHV+T8U3P3ufru7l1O
3DlgtZzb9QxCbOjthp9+wDkjygH0eUfDrEl1ovhZG61NroaRT2tO16icpzELd/Uk
ooKmi2MzijpAL/xvQdwZNIIyTcJ3EN0tfPctFNQ3RJApyqjs6Wolh8CiVW6KPM/e
5AISYDiqhF51i3l5o/cNK6vtYgXMTcYFzLsyPHYFX0rnx6Z6r0qPI8f46D/5Xh91
51YgK5nYwXOxetshqp7Y//fEt5XRoRjoTnElXT9BOdD7fHYcouIZShmkelf0YXVq
TmMF5pB1d9eDtKp79NEdbM/vker3Myg8gozKV02nUa6eY/3SZ9Vjq5Gmiw54tsuV
aJ9YKInebHRwkXiUVx86MeoESyEeJFgVtLs1D2fE64zoMyqJpEdSBD9pFAvdZOPD
VDvSxmXESNAz5Xl+x8pzzQFstuoKCDj40pJVF6FSGaEpf1/QPWlAvFBH3d1HJjvD
+EjPiO8fPFufMm6Oq2HTZCMosVw/yLdFJ2qaHSMZB2apCRq9zRB+sYHAx9qY1EcG
+dhSIHDL6bsu1TLbKVhGlwHoZ7I4Ydn96L4PhwElA1USCciBRKfvYttEwlvP1IyF
m0mUrqjHWl46NT5KpC8dLJgD6bBhGmFaUewgnmBWrWjo1aod8edvS7WNbOjIbeb9
hY4mRkRHlvA3xNTr4XHb1lLOgt5E8WYZ2x6cJgH/+/wam1GSq5kFdgwf1SIO+ZdM
nVOmFQtq/SCu/RHh+v8qGZtguDBFglUTo25zQ0KFF7+cJebuKTqYu+ekrrSnfFzW
W+EiYAno4Gbg/9deEOf3Wledbkjgo3BsmArKT3OsJcmdhUnTw/CDd3D8H1hjfpZw
jVvuwVGGmP8vZEbRQgwJHaSgXz7GOia9PxioiQ5Q1Nlde2PV2ezbExnUTUQCy+lt
Z9f+74rflk62y6ITtwVAD4VtxDHTbROjNZJ9fUpSoDim2hDD7eHa/ocumGhzx++h
86GoVeBFoj8vrBYPaYob3UkjJZ0Hq2gOUc6hCgJ3/5IbLTedM/JUK1rClJdQWuHy
Nny0rOtYAtg9NUT3n79xoUVJw2k362G757bO5PKUcQo1m7inwW9ZURX1sLi9DNgt
nSM5+3x68GDmlCbt4zXC2+GrYZt6oCuRoHT2ZGczSy95plZ4lFLSTqAgJbs6jwo8
3uUbraOXy51ZnjlcsmnHqGAZB7Ig/66kZnWmvXL0fQaTUasOBwSi3X0yoUDmN6uA
MVBYwawVFt4NFsWYBIGLPureAC+YnS3/QdagyIBJYjhqIw9+f4tIQcGWKIdBPDTM
fASxUhx7usJEtLWLZd2oyKYpcjvDVEKSIAz+d4avNMLEHNU5wYrjK7SmL6gC3yz6
YriIGm9gudUSsxih5Ub7zhjFFxHH4zZrGksPesfCvaU3JopkMZF1OyNaK96yjiNN
Uwtf2+Z7xRP1Hyr7JP+tcppsNXP2bE1sPwM4CLQHUHTaEG42veWRu5tzqZXkq8Ki
eF10VEZg91XI68w4GMeVdY2c/LUDmgHZ4n6IF2yng70BsHewiCgQ36YAAF9/Dy72
mDMNY2/bwb8aBn0J6/fBgYxK4F3vCTMVdkqHbeHZe5qg/x7i8Oxnt/Sn93/BGPe6
JdLcx76tvg/m2VCZH08C6PE99ZTDPJTxmHOkMivGM3vnv1Y+nspgWkrjFcA7IZPM
w144wOyuAeCbWixGEHJVv2AXk20Zkt/0j6lth7beK9D9b1kzNSKzgHiAKju0WM7J
hrLyS9kv0Y05i2q065KoV1OcUk/xXi75WpyZXBZlLhFXRZB3zrGhVWlEgn+lZlEH
N5x33uoST0HyNzK7h/dArZW4hdsBdaXrILHo20YtlXYoFtf9qhiba7hrynge6+S8
LLGrrdcam8mgJ5D029eucg3cfJlO4tz7XVglpWQrNzpTXH3ZOkd38DuZEFXvMjR2
K3AP+9wCUjY8hGf69RaQCPOLiemF6Ueb6il3/ch3TmpLAOAHvBFEZYeWNbC3T6DB
EQFekRrL8IpDJSmZLd+KKDRhTvOnGGkipzZKOGNDOEi0ReFRZBG2/d8O9eCSAGmp
94rt9JYDfFyfDD7vgD97DabymUSKbXyRS/lR55lTaUIAjiph4cUiCjpHwzmDmF68
9yanHT1OjoXrDYN3ScHM95vwth2D++QOuy7r+H+9aWq5kn/uBBrZ6Ak9B3F2eCbe
/P0ePzs2l01MsQCCLZQLAL6N9dMLpEWmxu2tys7ooKHuCp25a264kvtL59we9eR9
gz2fNDUSVXiVY3nxMhSD4YVVgyaAzOnbReIa+HhWzBjJKlsrUhy4/aYkZ1JykLZQ
qAvEYHFj9EgQm0o6S8D4MZPuihvNvqUajSmRu+m7GqSIy2GyYm4EsKBsSv22t2EM
xwIY0j7+lct+X4Bam/b01mkHG7lobR0o6TxzN24AEBmQ+5DGSvnvDT+THPWkstWB
il/B+qeY8nOpHxVhDgBr19wrJ/ZZOfnTj33WWTeDBnhBx1V0EOHEVlhGdgf0igat
igOhazMaDCtZGm0tS5xRWh/HyoY3Q7V4PEkWHznTSava3EIB6Oi7MLOM0Heatp5w
HdNzbp/UGNwPVXCjPPZi1TMGRMitlRXWgIgvnZbA+vEHNq4xcgW0SGYoxRyoujJR
La7plcYgpWzjTPknJTu6bdsNZ/3QWrkjW03QWBO37wA0wP/DVLFO4doVyNmTBoT+
ls93fD9y96gXHjRg4vB3uF535QR2W73ChUh/F4KfyOuAtHoCf9+FWrP2Pb5xjWRC
WaMP3EZumcaGxg7/wRSFBltlac1rpah9471PG4cf/OJNhz0zY3ATJl64QATtoEqP
/uG4K+Jis11XvQa1Bmd2WQgNskVN5GutzRPqb6gq3IZPRGsAlfkM6eCyPb8TM7hZ
HlMIXoHdSxZXseaWjM1up2261wJc15FbxL+PMabmpdxESNJJ4VgBbKZ9VCGbnON2
pmhtme7YpZzhKDr5DGCAEYdwCZFYzu0vUl6FAF6l51VKBuCoZUiLJp4vOuLSsoyE
KAHnNtDrMRxjrjp/nspUTgSsvOpmWN77xQZWhc8rgObDFeJeZT1hFNDnxkvRdr9a
7AhwGYSCwiqN9WfKx+foGrHUP/hWJe4XgK139gLZjZSq7T9116BQ7iY6Gh6cprh7
mDrIsdalsXqOIlHpGxCOkpetWT7MeQ2myZkVGTdvQ6d3J8wBZeJFBMDMTf85YNhv
4jPGWeyJT2jcEeT3MKnNCsnQ7HWg2YBrzy1Ghejw8n4O1nT1u2fx1dkZtRqU7hud
XUjHJS+58V8OcI398AAmLkHWU+2A6fNrm/oRl0gvB603tDcfDk1ynCR/wVWqj2Wq
hiey/1ahEDml4PEng+NMG3LQaWxhHIfEputQPy1wgf2gzCcscf+MpI+PQKwy5Ene
Z2ka9A9EzJX66TJPFz4jqqW/jaYhe810gdXkSLeauPYfVjzhCHpfgLogIbyyL4vX
hr/ZsSMjI9H6RujYfoFb66arhhZPBgsse9TQV6v/FqepxkewSzgi7UjfK3wZGe7O
FPSDzB6GAOeuzoLRS2+2MO6rK5fziN/ENabltv10KeiKJ2Qy50L14i5QjmW+Bp4/
K7DIoIAAoXlA6qxwTaovO7z/bigOoE38fKaMHhIvwZcDSrU58d0LEB3V0u49oonX
4afeXMBn3EWt9CSzj1LNpahJ6vri5q5UeRSAmH5M+I+f8SHTELDccjArVNwGVP/N
MKP85YpA0VFXSLpDjf41ElYb60pbvDTQ1z/3PkqT0bxzotZxbILqWbQUc93H7cAi
rwSaJi3lIUJh6gN8MS6/a8Ozmu1p6/8zwro+NrTW+oo3KKik+8zmuLcxoehA2p9r
Ky/Cu/CfC3WXp+uMOffmR/dLppCgPYBn5YWY/5ckWCnGsW3yYntFHFaCPGhI+KCm
GPk+VODH5936H3yUnz+B7eOFHJfnRnAgn0LDc7GdUcOFMfZ75CfIpHE1ugauafh2
/LwOD6kVpkAzZxg3EmmmZmhO6W9l1Km9MLsMDG/i26+3OguXl+jmQjSSoY+ttPTM
nfCmhOMRvh12V7wziIy/kOmJRDDb8dCg//SACmDGpTDNs6CHwc18JtBCLe5s9UMo
KnRtm9ZLgpH5XwX0/l4BeZNyiPJ6XLDbm9gWb+qv/HM32J4WU8F2+3kC6Fj26+jp
qsDVKHXt2rDzBZORxtPjF/u8ScVc2LTryffxZAB+m5xRj+bSQlDJp4wHKXlPMKQs
2zrWUoHY25LzDlkd3+xk69tJ31DHj3rl49OA8ao2BnUsrPFJNTyDjOXebonr1izK
DSTW93lWkJ3C+Yx3WJAZMkYEEHlD6DkMLfpyInPm5lV+i9hLoFE7PbBZakU9pxwV
Vek1VO/AShAGH1lHdW3SDc7O8U35W3KXajp04mlfMl5u8yFoL0noRHT9cVKm3lRf
3eIO3WCoEWPwVuT1wtPPgftzznzBf6Ev2NM9pqlQY74fvXS4HYMoJudqg1IOoW1Q
0+aL/Z5am09MrgnyANvNObC8RImeGe58vJOon1oe5k5RmOzvtTuFE+3mFTbOoztA
jUGaObPYB78TnKkjvlWZwWph5+tY9dJZaAfktEHirOjyTONNx/tfwkH3mJFXmCA+
rWTAFJFUQEFHUO64f3aC2QTVsdwFHnu1dESSFXTgCGNlSSal7Dj/sUsFSF8aWBz2
dkGSJ8Uq3ViPzLg7QXDpmRsHG+T0lOqr377vfLYkzaJdPPCa/I8zP5Ph0oEsUwl1
R60E4rfza2SoRQPoYtoufUWtCcZzqqi9J5i6l+OnlOmepYugD1zW3LOglIML7KZS
rPpamn40gOZVok981bYps/pnOxyicF9sIdTGXBk1vJRs+MXKPyXhb4gn1W1yJ9Fr
2fu9HBVgmA0go7rMpeJEezUjxd/bKRSEX50lKULQG+m3C3pFbG1VoDHy+19GlN3Z
s+9SOy28mijf16inqNpXL7XbpkVn984gaiDWT8afiATgXVnPgo9u4jydEJWFJGnw
L51p03YwdHscYdsMt3gKneiBFYxw7qeU6kAuN3lRgQrfv9flrmsqD6+slJakKK8V
XWJwkfz2TX55ZRuZBh+J6MmaBmagZxHTOGRLoISflGBoxJjlyH4MKhu4gaQ/8hVZ
wMzuJT/1aSp/g69yZL/5demm/qHZsvVZ8BGi6C4iptBUpJRTXSJrAj9NTpgA8W/1
Df8y0xQmLZEChoJ1AfR+BxSWAvmVoZT9uco9hRkkejtAnW10lzKvKTfJB35ZFvGT
5r2Lv+4h3aVfgerbLUlUQJ1Wu/LeM9uohbLh5RUnBHdQZyfy2kwh0QLo+J02TCbn
pYEHrnE+7o+godinykxU59NnjUOVFDKvQ4AJPstJDY9/385b4mt3QU6pha6zffxN
T1HlxiXPaYI3l+W/5Jl+yfXhxGcIM7MYUTK3Jboz3K8Aps80hOJu/7JrjJDxMXNf
aPdCqSzwWnXRWZsbnZRiHPNPtMbuY4/1DXyp0qnOdynW7nOE3VByGJY6Bw6iHHJN
uIITXUDWfLw9dF5raHhA+D4JujGPS3BixKFVbYivoLon6/JSyC0Gi9w8h4tJAREq
tYemK+6OLQSZM+lRixPf4NLDxzUEUqJQ6fmc+BPRqZdNgbgBrVClaNGT/Cs4M3aO
UCWWfAkAxRnE/Kj9rq6FDbiS4p4NZaT+84DqS5WaTYbb2gLoiAGn2fC+HuHra7LA
q98s1fEaD3xfBv7o4h78VKxF9/FZgXuR2pNN+68sNozMSSdtvhZg5g7eyXd0CX5V
rELe0kzijiXybsIWef+u6UcNoH2McOFvYiA+0tv5TS77w0FSoWuDIteVdvupN1DE
2LRRkZUR79DCnkA2jVsliqfLRfkBighnxgmS0aWsz43d7RHcgHkcwXNB9ZXs8lkP
msh9WDHu5/A66Irq+CLJPzlMRW2DPTewbcpJhJPvASbIQu1MoRRXhivg7IUyN4dN
7MLPBWFItIXXAqAS3NqEUNmeViJIn9TSyBG5mcZ61HJdTRVaxSCx00CmzjxaWlpH
7f8JLZPDGhK+5iUclV9zdT+4kJ2eecwk66P9LD8+y3ts7SddD/zKPXpj5qr7CAqW
Ybmab5havI4S4G4JEEIM3Fu9XA8aQ1Okcg2uHd1syAuRP1vDY69n0TQz+mhVoyo9
CB2NDAGH4X1Vu2XR3eIJk/WndDtmhlEmxcjznYSuU86IshE3Rq65vYLMIfKcGmcQ
KgJEPHcIFs/dtHHruBHK0tFoIBAHuPfI0aYVo2tZpeB8CrdV/e5cjfd/ypsuESwq
XRTEXtisgZbX/L18Omaazwd4eUplHpV8x/wZhxYia9PNo47BrR6LOHeUuiwpRJfc
kvrgpmnEUK/PDQ3vqTILvUQ3SueD1+lPmFTsOJ+Z5Yy62+BjOnw794WvVkqodWgr
AYYK/HVDeF+HUivlGGpFyccokLOcoGPVpzA5dGaKqRBykdmrY/8YZIlvs9t0LrNV
Z37k5SG5eeFnO442zQNH1xO3u0pE4XMqHFvDjHONAgch0mAfKPsYYAWPCBa2Nhxh
083NP+tmBEFKI7DLnuzfYJDN0ENgsEEGUz+/oPngOiXcaT+HMjuDh3MF0Iud2Lw/
Q4qyap2+nuW+IKPwuslqO7NXdQOnKHZalzZBYb5JoE3WOEaPuR0/J8u+MsjsdNeF
WVVTJisGpC4oyK3pQfOQ23hE2P9lpN32Jin8jCX4lB76/5yDhF/KG88xzFK3Kv51
McIMFVYSjG5Nae8FB/yTdXg65Xqn4JDbiQ3K11bQyc6uajiZ4WHdxjrmUKKZcM7P
8JrwP03SXt5byHDggkdCcjDsg55SBBWuL3DJl1E962NCaB7uXgGFPRPOKc0x9lIO
+Qg9AARyt553Fb1GgrgaL098TnhO9AhNeSV3ynSjXFj+N2vcxgb3hzLlpXN14vXi
feqKSH95s29sWDpNNj3uLhi2jp1L72jC3FgCPcLaPu3Uqwnc0B3gkKAb/zFrSCp+
YQe/sXjg3SL0CY4KYk4DPKQdx8rWWP1lkM8jnFdl7fqBgaqEeSos2RDp+te2PUQG
rlhAvgbK1ygA6gHVaghiV/cmq4YC/QJhUD2Srdvjn0UohynC4zqYK7W2iy8ko6GX
Zcgok2A3HC4cMGqkKtZR+Qm2ZYuNnrYKSY8PSRrJnD/XhpMtaQ3XefII4XjimzJU
hV3U9R2bBUP08VeAmzdOu3yRgOZG+sDvf6bpl5FsuaJNYuiDExGfhRT3ehxde0bH
2/qeroebd5Dkrqonb7YKsh9kI37n7FJhovjRyq8cQiWHLEEBYLqLDYlPWcnWVClM
qOGpVnoEO3AF1e+8bPg42ACYte6KGRZ4asW7wdTc7Kqcy0dA4j0sJjQR8DJvjtew
HEq2bP7Oh0tyZpudSX1gWVnAtO9dGPLx23CTYJ6Wpd9cT8Vb1YqbwaZC9vePjC04
5q9Yfzx8UCfjd806RxB1xuT6BtitpsyP14fFGwsgMY85o0lo1oxfUUWzKHleKnoo
Xp59F2KnG+mCoFfk2qggp9ac7RbC4gw+8w8Sc1YpXqVXkaiUOEKD/f2RWwAWi/7k
RwfafPBmu8Tkiqjk1AdaoERzHuXX4NuOAF/j7PuEVeklV2eitAqIvpU8kBWHveDe
nLFwi01oaSTTW3cz8+Xow8XIGz4UwaCrMGB030nb3z23vjms7Dd48w9gatQ9N9fz
3mcGKqlDXoN+1rfwqSBox+nIf8dFeqFrpCAQFF8xnhfEgdGZ4c5OeZRBvilbWZbH
QC260qqoklG3AsH6oTE6vktkZ5Kslyj9cI5VtpMEvdwJ0FD/TRryE6DJvOax8I15
Q8mpUaWBv9y8Uul9sL4Rf6KSI4kVcUlWLJlZ1A+5PgfxwvLhddrkFy39SBKsXF1n
vgm/teJqB/+wZpX1R+neQpMomec/Y2/t2Z7dFz1eIyRMWwl7WmbAjnPf4kQm9NPh
EzxU/FGQ6u5rBRrl37jtxTRMBhtjfAr69Pui2oV9mHKm+Ppp1JDmtPgyxPXXKeyg
xUfJm4DemSK8M9MdKt3f2xG53hm0o/eZ78RpsVjfDDS9DcD1AVFzLjz/93nnSTgS
xwPm8bcs8wAp2HjYPPPi+0W3R1lML4cqQBefF1JHwzQ5X56N06hy4JRd3aS6Cyjh
AKE9mFyjn1T44Y+QiNmvo9emBKz6q8pqxR5wqH2eSl0E6/B9Ag34dOn+zgPnBUS2
3xBrTQc7KLHwrmfSvJlFIzufRuC70SiLa4oFezN94V4LN8j88HYi8ZLTt8+G00ug
T3XexRPXdnHybuDkQVcv6vMmp2vIU61Ss8RbEIAqmEbba3nJliH8Sen+vqieFPvE
tknY1lh0kQtHJMBeZixFoZ/FCLx0maouoeRnUbkOkbd3Mai5ntlPfRkllwmCA5Mc
5ovtqbKLL/Sjlys+4Nlq1oMoDxksvvaRM7Xqmqwn50sN2shf7G5hDATtAgu7ltMZ
GHSRBt/lJDifeprYW7SVrXc88SH8Ok5fwODqyDhHfQ8kQL4Tc2O2/o7xrZN2Zq1l
9tYpAl87pIUY2CI/C2K99hSeIlrEkWEQDOHYFa+BCFWpvxDILqCcYSyZRJcGDodf
t2KSji38tUJP4MFnIl1kpooQYu+43UKm19vXNcfbje4pxRd9wHrDzNTVGQOa9+vU
VDoTckMUQ3jCD3U3NouZV9Cm7XeK85bu0EsnJ2Kb26+PPmE/XJemjIGw92u2gBtV
d+lk+gGskJw3v+4CQMCOGpRGX+Xs+A0TVc2y3GGizbTj9Ga4nSwLmN/rIGsPCfLH
tLAmFgx8/keNuJltT30Ja7vNa5Q9nFIcJvKjQ3ZNAi/Y6xCIombETnjGArX3SPCL
9Oo6cP8e5isjZT06OT8OBlR7dr/tC5OhOlvZvM1yaCT4qcGQVvnOu941cDRPM+e9
B2lCOudLw5G/YdOcOWjvG9D4vKDKwvaNPFcpbvsI/ezI9eftPhs68uuYsScu588U
tk/G3dL4GHx1fHeDNRtGmtA9XhGOeOFmwbdIMpRLGeiolcpEBK/yA50EMrjHYSt4
CRdrBpkfkdtZjx/0Kg+8ndbPmi2/3O8PuoNDpD8WbLGGxEM8uR//qx4TZgUy/lFZ
uABAtK08HwYUnMp47l+BoMD7zsc2OByih5BSnnXviUo+WpgsUiicDZ0Qe0/iJi25
FlIQOq0lfc5Ziv7oERzUNeOlY2VdlQqQ0pcQybdIcctB22yLJKGdRjc4RrX71Zi/
Aof0RVHoElmgDmsTfELoL857fNLqtG1boU7NlCyQuUA7wMi3RLF5LwitIlm4WGWG
QJsIgJ9Nsk1bbxB9mWIiB8R24igQeXGwZDM7TBnRonKqI9vuFvgbeB5TOboYTYhS
Q7xLm0miX1YIyyZSnxOELmfoHhMrUcnU8FSFfZR3AvaiIYkyFoaXMQNdumx2/xRm
i4I/NjeqD78KNUztMyDnlNWVLog57PHW7O1YwnYV5+j0aJDd263OZPCg0i2hcsCi
MnbdhCONx0AbU7s9jvqLsEPF7Bb75CrnPDVP9YXLCWRjfk0HMK0URlwNrlHoL426
KaF22HJVm7gXs/bjKW+VXioUUUjq4NdqlCJwhyBF/Zp4NgLwqvTraThW0/GTPqa9
G9O/A0aUfgZ7yr8e5MWhiv/bM1VppaPn242+UEt2SH1xBzzluZBKo4bMV51NbTWI
3TWQULlPjquI2SKQttKNF2s4mYZhU3ctjVChwpmTWsn6St44E7y0g2VwTN4Setss
n/H4k+zLpPE8dltZkhPaa9k6jtg7BH9m3QGNw3RVX2+K0nk6kFBHGWXWwa1LJ9Fw
H7/J7eE03i9AHiuN4zi0295AGocFpsmwsTsGnD3wkMTfrDGnwqkIBGYeF4N6qxMF
eCgxXifSt7WAQXir/KI5FbxCotsvXlSOdMxkhO6FqFCds6e3b0SHO8hzRAUcGCTT
mSXNGfIcfoEagpoRAfG0mp19gVe18IZkZz8j+AmYFiI003ml+IVYNWqmL+xzBPFF
kMmjiBYSlCDoLkKm+D76ml8ear215wzrd3zzXXv3M2IbbjR0Mkly3TMhXk6SQNzf
CbgpsDomsrnAlJnnKjqwiFH9BDGoglq5WbLUM1QohdIs7cgkfmlXbo3wLojYn4eB
RdaMGej5zCZCNC/enrjhR9wjx/RafFwl8xD+FQVKGUZfxe24HqxE8fqPf/X9QlBB
sqdbBm0+jrsfiHItPLsT0wAuIABdqU6Qn5mAsl8lHpvacwyAiNR3ECOl9KHCt1zP
AhiqpgJruR4Yzi9Hsx7wBs3Hbod3ldkeWa+D3ZYMU7EINMotlGZHOaEJQci2x9N2
/rWJHb0o1km007Y4zrokcWZKCiBbWCo7LVls0M4LQ3FW3lgenv7WwD0phjCSUGTi
8puPQ7UBrhZGyx+78cYJTZR4Zn7S9CWVqTTScbEwxxcyEGKJmhFWVbr0PiOZfS6J
4zNpsQ4Nd53XUuzjRKzSRX6Tpp8DnTt861e1wPqXS7PCxto3518SMpPEG32eKc2M
Rh3Q7cKV0VqPlKLyY2KQ4XDevzjGZGyZZVFgwn9Nks6ek4gNjGC728KhdGKP5rUF
ba7u6FNeiYC6o2W6/PTwyW75YZpSMePkc0nN243vODOob+twPKU0A7+mQPWRgNG8
mdRqXmUlBkT9HmlovdXYUj0+9zNRYg8BoZp/+HyhlcWrgviMGt4sFAJKp3no6l8T
ZiT67FZqwQNa59ogXRa3J2/Tqw8eh0YybpJg+o6+IP/2J35IWrXhps6tUiPKxtyk
4okESpoc8CDwPIaT5+Q+5JThRD+EWpz0OtnM6G3TozkNn9Ni7Z1UFcMQADumRNTu
WC5Xk6CiXqE0LGbbyCLS7aVOSxPxSMotCiHr4jMq1SMmQw3Ve/58ZA47/NcQjjOk
/4cmptp2sg2ejyEpewROBeirPBFBRs5AV3CyORSGwHm5TLWOBlQz5p7eRvhbInmq
RW4Qo8NAFV8xJx0TLdlLG8I63pVDgRdujNie0HUNGzOjKz0kii6ehuk27ugbOZHE
6GpRRlEV+aIJBx0R3bjdnD9TS0419ud78nmah7kZOtYI3awHVHKf7AoXb1CVDbHG
NI2x6n55Nm2dNGPC+CQ3IULmKu5czb49G7ErrsnU9NbwNtk9nZbvA38zkpnJN1s+
d0whHwNJ6BN1UlufM3K8/xxH2WBasFc5o+A+O9fNsEGlnXhF0+P2ZQ1ENmeZM1JV
91hS6JmpqBt87F3WXCqIlkLVzRt9TEI1rYkBxTeTVC7Hfg+E54O3XOxQI+YgDF/0
HVUKW39dgx1fJZftPLfalUVS9qAneuK6tIpz0t3VFA8PmOQxRpR8V/DrLjWIlapG
Y7t/BZhWDIWWT4bY2CL1jgMT0hPf6fXREFmEx/9Bhy/bt1lQoixAQVgwCwL+G4X7
qvTL/9q8hP0Hpl5gnSIWZjrRjJ+Pz6fkwIbSTWwpLCsEnO8ABLii+6GPcogfpyZU
WDi05qXSvOs+sxl8uwbhKOYG87uHkz30ZTUnFtfiBwKJE38yLoWigaexwiFydtea
rZ4FW8OfiZWFxByzCyxzQWi3IYvtYEiqcWIxq40t2Hki8MJ49r3sLjruNGRt40lW
/uCqqX2ODSJK4TLtXUogbqyIRfPiubmlRyhNBPSnE0lElNrXTp/KsX8Ze8mHGvHD
uX8PhDKfPpYHJKzkgTkTHORXOMM1DFr3vAp/6hjTRu4FOqwpGC0R+sc97R3Z8g3T
Mjf9T9T2gjr/ux3Y1YEWhJn1YSanlJzl3vyGxXUuOOXkHPHxHm5jY5Yt019mslpt
NuZXRIw6i+vuiP0fRBzcM/02KawG6Y1wpa9zVClVVwGNMm0cEefOuAbTxdCB4LnV
LoPAlGNR2QNQficF4IgKB4ibod+N5brIQYZWdkG6lDXHbqXURGvbLIgTT6dp/Gl+
P6PfwZkGWDvd+YpQRXIEVF2Pgp764Kdwo8bxwRgmwAscEhAmzxoJrRBgZo5pz7pA
GNfp3sKXBpobedPEr9xMRTTnerhq+xeK4D7SyW7MVb285rNtSKBIRXEgpBC8wc03
CUefNu0zFaAqmkglw6oWmavs/ZyZgerAt4CNxCOuI/UkU0sIhYTKaFgty5zqltzP
2YEC4CTYvruidwUB7YYX47jZQX/sBgbdmh7Tr3PeVAVReQcleDRexpr4NGMWtYx2
ybIimLHiPGOpEypJcZnViliK1+GqcOM4bxAX7ZDoN6n3hTzF0ZEgR6W+9hkkmF8w
c170fEjWeqHyOSSzQqGZCGY/MyUhEfIS3ttn3FW/5Vj/s7hE/pTHtgjBTJCKos/L
Txzo8akZl/Qscz+eP7v4WN5cxahRIVO1qT44dq13Ni/Qirt44pocgAb7QHxsCTzc
c/stKI8vAsLbbPS//7EIjDo8HVuFvHDJHZ7HPN7A84LTVNYbY+Wf7tQ6Waq/hq0I
69NSQIK3sZMpPMfcDC8ghVrIaqxJwsZGrQ2ebR+JsQ+QY53mCCRhzJerIkNlj+IX
AFSs+EQ0PQMDCBnPFdmTOzGxNmfFfit9iolsLe6VTXvrdDDGnzPYaRuEDs5daEfg
d3P0X2g3SZDzLoq8DxiyoUbvqi+5L87JD/gpilMJgkCaMfL1nf+TfO9kyeDrdYB0
HfMggX91OBgxX11oiGO7dnKd/XlgsWFY/fj0zuFDjaMrlhyJh/nFzJfW96c99lha
fmhIqB8SHaNAf2/XMSaZlkK9UvSrkMNIzZ0Q8weUY5BFP/43BeZu3PHciOZcq4PV
tLjqtEScpCIY0LRsqv6GN2FUZ4fRfc5mz2K+RCvtGAzekCJmgMRHt1FZ3Sk7oO2J
WTjR2NwEx/8NnjHuCgclTP5NNlTe+I4bT9P7fxtaQx7Wfg3VcmSJyAXD/mAvIpH5
5lgaU0q180UwUxjlUL5oLi/IbXSp7svGfEDE138JKEVbv53ZDe8s/RboOLMVlbWj
R01+keWD/OdavU06gPK62ct+Jbi8KrIhOW2HpqaU0SefsZkdWSAz3D1ao6rSyTIG
XsvkNYokBvoVJ5xReMcxk/m/Y9owQX5+RvexVpImvQcb669yMhuFhe447i+yHOfH
2vVAVUOvtQ6XU1ADT9Da3CEgd0mkBpDqP4E3R3cs/f94VlNAsH15Sc3OVKOYTzka
nLwBXpWDjuxl1YniYeGxGa2sUoQ0mi+y7LaAUd9wdxLAws18wEPf1CrlUvYqMnDH
e7vATBJqLpOLuQyd5k2FIun2UKJR7y4GXDFUdxJ+iIoR2+jd2rJ66IVi0yeedLvr
q/+tAXKFb8acWMk1ZjqCHpKNXSV1bg90px3KCmkwgs/6beNBhIZpiapdZ9h7SSX0
giFs/Y/mpKXghmB6K+98KWRedQVkuFSSS3VceyvKeHkWnkH0+rYI7h7SBxjIR4+u
D0MU1CkgcNl1+m6TMMZbYn+zFUIbTpG601TyMRX7ropNUumjIvSFucSdjRQ8XYKn
4r9BhCtu8zc0gYfDK6GINB6cOtM2DdO7/ztQxokEw9FJzzvP9tydC0p1E+nrSWzP
pxEMsiDfNQkD6sTrZOYrZScJMSd4oH7UqKSWXC+TL4WuZLg37IrFErtFxH7kHtAy
7KaRVTZlj4ZpKTugYs9CWuDl6FpoPAVXueX/mfByZSWX7Qk2wX9EeZQb4tF4ho5+
HpaoA9sJYxIh5jvZ3Is0XhfA/xDXcuC6LLSydFp6y9NoMduEERZl10RBHxvCIyPe
cvDiupkX9fIta6ZuSI51sCvHeMT2UT2xDITtAo3ZV9T/8beYHLHZE6wOTRV/mK7A
w58aKi4g6m8xlJg1pAX99tcdVhuuKGagp7d90Vmr9j2rlmQE9V/6bJSG25T5O1vz
sitrmSdF2ntEBIqHRPRepzq76FC8ohDw5Idf/AYQL+6nqcppNwJXpsdyhIclrOD6
lq5MHz+Q+4N9KxjwAWarYOiQE+RkabzwqSTpV2/C1uxKSZM/8xdf1JgsB0bD2xZf
spZqonQL8Yb5SlrMtrmHcdFPcejAiacDAPrbWw+/w361mj42KZHsKZzXrax91GuO
hhjK4WkRgVH/cCrg9fivldLIj9Fj6AKHABI+KE203nViLQxkT5oRTLmQf/FJHr1g
UHhWvi8a2QmznuamKwI4bFH6DS9eTjYeGMMO+TykAQy6STcrq4bzSRPJS6gX/Mm6
BiO3gb6zFlBWKR0NlKywxDsi0EZbmJe351udZ6Pdjq+libE6rUMrLupYtYcBvjO7
7NYAjoEiq7XPtte+f1UpIBogA5VWCo0Bpx8P+D7X60WJG3lFuJGm0XrZewjZMxuN
pEVgRVp3DWjh/7VgR8h/gqxvoLXfHRuGKCTSm+goEPZ+Dj7mT+g0qbeUEj7L66QD
PnuMXhUW+Z/wygGfgVgD/5zz+dcuWPdF6xPDVTMnJOb8FfPiIsSjqJ/1qPCPNYAB
mbnU6ZGvr5BScrM+FHoqodqMoZPShfewo7fGl+TQMBaZ08hr4vEpG/7z1U4beWHk
R8dFTCG93koF8fSVndoVFbQ3FMOubHMpd6omV19tw/+xatAXxQyyALM9yzn5dRZq
dliERlCIPKqoEiXVgrPlII6LZGpeivkqAGUrI9IGG2K8BVKSYvYl61yruE1ufWWn
+TiPiWF6jrwhAlzB1HAhfxewUuadvLrWjCNbM4KR2nWNO/MhLnMR/Se4ySff86ZA
1oGRaD2t0fa6aPWIhoE/Zb1DZRzX8dMkMpMSbvApZFXtKu/RVAPqt93ba2/8KmaH
P89e5KBG67PW6wFcHVXOmUJWxSbddCZdU0ZOMpcqM3/AUQOctQLPzZgXLYJwsqX1
bW9HuMBLPZVu1q5LUNi/kZK7mg/TJ3MlbUCKT1B47aZt2WmqBHi8RCdQuLFrvg+b
udmPR839zgQD5+t9hgVa4aXJJ1VfByKmzy7KQedNDPdg5Ggak8nE3dvk4oEvOxve
oGO4VSZMf9MCpjEqRNw0Jy8WDQPzpe8SEEfv4LBB3lFa+dTPOJDt663tENEP/KLw
YSk0UleKI2tmK0X1wyiX87IymNPk8EIycOWAH4aSa05DDS8wY3sosGE8+m4NZ2Mn
GX8gFiLvgzAt4O1bgb4F3e4oLo8RvMVHnQo469oWxs3sL86ux8ijY+ni0vnTCsGq
/H5fWQyu4XVqpkYW5KFKq2RlgX5GTcuo/nMiYgcrn9MatC84fl66LsNaQbpGvdPI
cJMZgsbR2XuJitQYaAI9dCLTJwXnyRvmIVBZx8ZhIA0MHmwUHRqW58dPEKo0y/i/
24L7JFLvggFOpXrpjCePZ7L63UHV8rOsujCsMkvMFrJhMCZ5arRtzvyNkgrKXbt+
cQhp0d/wQWJ9jbQwCOngJRmCgtfeqZ5YtGGYEL6qrWiqQC9nrq+1/xbYWPUgbSr8
XKh4oJILbi4dUwjA1l3GHzJZJgdg7W1U+t9az0oxw+RtUZZ9JznlBdMMQ5i5UPSX
lDbmfV/QEy3EPUKDtav5Ku3xftoj7Rny2DdUB80dIusFwhgeoDOK3HARTQv56Gjx
746n/enRafljVnOJjX6tn9ITxqAZTkJp6vlArog/bjbp3mKUFMdTew6JujgrXGTp
jwV5PsWR+54zKeuJTrfzBSLKnK2juYbSmnH8Xfk7COS0nGsy0E825bu9pO7zG59i
f5jgesiyN/MpxuSYbaniLfn30lDixXv8Rm93sZcFuYVJhttUEzEX0w5yP4CE/N/H
969oHJgclyxT67iAjiJAtps2NesY4/3bX4ub60inkbiFN6tKgsnz+1E/QzHjk5T5
ye7tXLlwk5xZ/L9b5wDoRTysrujP+hzkzuLyHRIKUW1noIEklXR8aRZZwqrnJ0B+
190qwxhPF5pZzkdypyJ1BknHKohU/oe2nlwEGnEMOUAEk1ZkgqSTbAwNOh+4TnCp
MAdfBaGIWdS4w7Eg0E5715Eue0LzDkObQWGkGu+hSsJuBs1F2O/XtWZITQRC+9yS
13sLnXFT3DY8gA+MpBj1Lq8c/jcCamSqOklOJZ//WNpyQXzx6gkdhnXjGQsP/AyS
HdfnaBuXb6019teliqxvj4s4WKRbrcSqj6CskqjtJpw17nQN7pvmUaPIgjDo1Nft
bqAxnNdx1XFpNVOugPoCQiPb6/pd4ekVLBSM9oAXsBymFr5MXTpxz6cxuxSrCrDZ
iIBhIKEQQl2mqPhy6XbPp5SQ+cSIDgHlEZ5U7WW96HQ+lWAKeUFdCuXt5subRj8A
27je7RpiUEkwe/AAhQUBADTTzzCF05jst1tm4T3riqUe0YdGXf6PXEQG9MmRc6zV
rSY/FKZzuErnex7c82f10mBwKEaxa+WpVlggapUsXVUyel7O4r8i0coJzk3UMMhF
8DC9GryGsZoFzgWTV6llrEaXfk4RWBoDA3pNKskr6XfzFiK5kaSuF6T9vBHagmHU
ONxw57QKUUVYNU8qpRK3C0qRAmBLVXORnRh7fjywXZFNH96LXMHXKAYuDmMFkLoW
IYS4CPcqtuL1YneD9Dwkb0L3sJhK9H4cR8/C4Vu0LpdlaRbjYZxmHLt1olfVHHKn
Ls/+xG7+RGmjIOBzp/3VtCaa4/QkAV184R1ejEeqjSrzjA/o1/OJBmi9FY6MSWnW
qdcJOeuUBm/iu3VOdtN78arH4aNuK0DlH+YUkEebXpt8TtwrhiOQcG1oGSJ2fP4H
eq/x5l4IcX6L8gI7xDP8dv/5up520lZQaI+lE5MW/FOR3uC0BaliIdNHBkgAH++E
IBQEWkyOzOaEAQuhOC0mQ8KCc6L8kNr/lICydBeeoZvLIO6QNVrALGAlzVLkd54i
8m6VNBzudBMzkSxvBOxKtowLMDU+SRcGM/ODPWzeJP+9Z/P+oCa9YI7Ix2xiKdSa
7UvTg+RX0MdXPluzqQOVLKTCABMfAp+RsOl4cgtY6sQyvJsshK/T5QJcnugAdwys
tTGQlUvrqhtaoT0E24U1Nd+qPTrLdhx4diu8qww4EvhAHUPQ/OMwH2/HU1TcSurZ
jnji6XiiHWMxCp/JNZevl+of7C/Lffx6WJewaGR6Mbl3pNmi5uvX+jMjuUOvcBNQ
Ph0bfNcj7KJxiF1i2i+SPaoEZUS1NtzzC4qHeobS+qcKOvFbt+I7t7Haum4rnhm8
HZ1KpWFdZpVMYS2W7FyhtooNc5+3/5fkDETEiFQt1KmwSqMrw7lj4AM1lOdAaGqc
8y4RxssgGUALrOYQ5qiH4LRR6JXP88JMPMtF3ZTDquUFnbjzt6qzb4hs3gXyTSIW
IZluaP67UWDSXuUYBDWbvHnm4nL3gSANYednvV8dAqRrc09GzID9q+Py6uR/lBgy
Mz/oY6ptII20fpKNn5BNNKE9yFghDTDuV8U5d/RQPWLVRUoCr+pNwAcz5I9ngpJM
pWy59PGFyxIdo/y0kmwOCvQmTn0H8Cr50s6n0T0cuqo2x5K/hVXHsPnNx/Hi4nSs
yZPTSJ2+Wd2w/yt6fDoEKf1STLDEVhFhSzVmnXOGo7QtVaqRqV1ue0PJblRSPHg8
WFdFRaZA7DN4ACtnrU9RMQHL+8h7PF5pfegTMFl4ztG18Iubf0iONSrS91geFm73
Gp9Tuph2rQqtanfC57aQRHeBlpmoD+bLXOL9f+rx2aK4mKj6df+a9KF8QFs68LsS
0KUTrRJneYZJZ+Cgz4mEo+TXwKvdU8W9tGOx9q/RuGWnT6S4JOK6yjp6dJyirTKs
JIhuFxG+4AVg/8OrNInWiYbYBll/3n1lkypwcEHYUyhkQPgatgQU90XIkAPozfyC
mjWMlcCi3139XBtffqsrEiHmbQTFTRVHvrfWUNwtAWF1gD1ewgi+7SVcm5VlcAPz
QIfhC61xBvagQNS8VMONmYCnwTGW5q+4Cboaq1ua9rvP1SzCoARm5YZhaz5G7VFS
knZ0Ah7REzmcfYwzF4zrO7P6EDOq7f1OImAaxsaAV77Ree5h+/W7LSvoe9YMVjxJ
AnjqfOfu2kS2JHc1WniLQGLdpysTtscfyh+QpwYSZFXIumtRkfBY/0jsq0xBYTpv
3F2q7rssiXYkN+8WY8pUB3XjZHp5g5k0R+0wQuZWjbbNZ9FZbwj0nWdu3fucyqsK
6U3Q4eIQ+f4eYT30Of7OitFS1eJ78epA+YGaHpAlUarw3DrBC2SAARcMHKVhGbXQ
KvNo6TxI42QlWCS0NMEvSm/658hV+0VPoJaMeWTjWyIG9LOtYu+Fq07KmMp4YhTw
yUmZv36UT2ZcGxHytn1dUQcv3O080k/hECjb1J90k31dWqqV+fvusdEa/6Nwtl04
v7kRXp+ROu2OqNMpH/wX5zWs2TV5+TC7lvR51H3lifw5fVJCnKPMxqTWv7ZUvyL6
NUCiXrUobBzVM8VR5K6YyEOBFG1ukURycoOto9x6CqlPKD49SPD2UVEOOZxLh0g7
31mfwDCioH4GY/BPt5sQVrDevpHC0uBtmqIBntS7l7T1y28my3WS6BO59kTL4q69
LKMSjElodbPa6JGfPwLTUlRy/Y6+8CYB7dRCQ84Le68E1Yu1G4mk22UT2qmCHkmJ
JyUpmtHcJ48rPxZy5IbqlS4cfKYPPi00R/cMkoDa+oFk+KbnggpgAUuCgZf1u3GC
VtjNJ6sYqtJrkW9sAE3e5HLsG6ZDlRi/ZPFbV+IqYFdx2/uUOPUs1dCYq6xVqJko
kedCiFMxUcPLgezyx1mPUxTrn9iVoMAYeSFatgVdJgEZrCM1rP+dGwPk2MBAg9o0
j2kNfisJn/odK6GeQHFWVQHIEkLqcJaohbrSdQWjszZXXVV8RtgCV/oOXPBlYghS
MxAf/f+ZafsYfOdDhA2MkqsfnNlvQBS0UvfuqN/uNPCX3poyCr2XDh20veRhS9lh
+4u2K7tPdsEnPPQ3YujtB1XZvwNoRHxFPTWVhNNWjuZKP4wmUpOAdPRcWBDF6hmT
UqwKFjvZNMqKM06aNaxiIsqqN4UF8rIrD8VNbkDrU2FSCu6o3xHcfZYibfeXNeNn
de6JyuJwOIM/WR8TaITF/UylrLnqTFr+CAWHo9F13piMFUYFtg2IfKTDPDOzjlEh
N6/EO+SNhzE9Dhwct4DFIncEv28uMPtj29StnC1i4Kl9DBaRqu9y8HvAEWCmgQZ7
abxF24dKbXThgO84qUwerSBzHH5v81T5P8PpsyuSKgsQ/AYUdD4liH2yqIK9u6RC
7DcR1MK2o+WAA658yhKqS1cjBdOF4MnWq7in5AHqUPqxR0mUNi13RBiw/ChtISBS
T/dT1I6kZ82VGBrntKn8S952Id7cmw2VvKULD3hI+UOcT2B00LQgmFyA9QSpGOyW
3zQ9zLREqr7GITVDGa2/SM3PetKwS8v8RRjuKwhZgs/xxl3BXlI6DeupFPWXL5JC
Uya7usgYKoUqsdDbE2JjQZ5rdr5z+OpDiFMiBbNomwHkMjq43D0KP2ATg1GtUHcj
uffZFWCQcgfsG4cvmXBTcEigNUQDeHMlmfvQWffIEwHgF61sNcLGDsOaNXp9t/tZ
hNeHQbFSMKUu/6YaB9WNSLtRo6Pk4Z1pCBngjWBRcotAFdCzMWs2fthowwmVnf1u
PLy3Y2bjOKGcG6iUzQ99HawIAquVOHG9xzCW0dT0iMBpNbgIjPDtH8jV5D0zWld/
fQBZK/sk8qtBq+L6dBilXCmwcki0xxOiNArswzj4Ui9hFrHzv3zq7qyE+TvnqD44
mub637EBi5+96Xxpf7olDCUTl/JyD5LynZHxDD9y5kphFvCIydeYNg9ktSi2J36w
qfDV5xAtGFcfncLzMilNPPbvpfiHR2WOvNLzGEgXPF5dCnggfCz9LNLzvn3sWtAj
n4yQr1Ndxuf/3GDe8JejJDGYYJESRr7rhdq0rO26sEiv/z5rDn5/2pyrEEjI/2nH
zUfewrOoV2Q4KGv8KidN9TRSUeowObC2WVnrW9dDbF4qZxIZdkBD/3Wb7ptblicl
RZswmLkJAwTln9knkmY6j5p+aWWToivdsIkU+PJZ/GZQgB6ekJeYe3/P2frMPZok
vyTH1K2PbQFyJ2AQUOhiFYWVJej8kQaPe/XQUiFGSDFgsu6BMsd+OhVGWgRLqmkm
L0xAOjxdJOYBU9AyQzRmEjyTCOYllQhQXmTEHJWjGqRZ5X7FIVAplZ46Op5pybxc
qkq2avz1PG93HrwBsvKhVi9GrqGtzK9tzqNYHh3FsXMS7Tj1rp8V6igTIRwxB3Kt
0J/apanPTfi2TIwqJOgFgAtkOE9ZEJPGSbcqhrai2TCzpy4LHeuzvxHXE/oyu1dQ
VJ2NFimpArlZBrNrTAA2TDG3NWx3/OR3EpqRdWnLKsRrv6XB8+Xjabtqqcsq+1mo
fTmZTbtuZkS11Uoi/luMSZ8p58Q6k/XHyA9d9NZKGDmv/1Y/0zUCNpBzihmpUFlf
Bp+DTE6DqKnM3jWF0eZxMgMhC1EYiKQSVW8Nlk8tqA8ic/luVY8EGMxHgMD8Ljjo
HZ1hCn5JtWjKcgHeTue6VO8mnvEHickdck6Ejp0C4hpYW4bpfRdz6JKshrApiQ2c
3iTJ6BlQm8Z9Cr4KTWmpOz6GkJ5F+y/C+MTRro4NJz2ebR/gFD7UBB0Di0xTAOVy
htBoImkzdrlRMX70eZkHNVGxoUuGJmYMyht1EDcKsbIIChULP8/QMGwN7GclhPiz
zfLOoYUlH1HPkTTXqzbinLmmTfcVU/88/nUL5blEmHokKuA7bAUjbKvvTA7EJ7Nc
c52ADfsZACua/vf3dr68l+ZJ2bm8A5hpw/MHcPmvEgIOLOWNPZCH1pAqzGPIN/fj
nAdefzRUGG95vlzCB/9E9Q==
`protect end_protected