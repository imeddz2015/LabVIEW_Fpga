`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 23152 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/9huKRhRMtvnNqb3Z+UU7TahEoHV+T8U3P3ufru7l1O
3DlgtZzb9QxCbOjthp9+wDkjygH0eUfDrEl1ovhZG63L76IY9a2P7WcriX4qPg5m
eRzGHCHEbecROZhZ2b1EXNkHSjSIFwESopBR3Mb5KUBJ7sLsxB7M0IYTPsjw7+U0
qlmnlWK+85CYmsJgpA8fDP3CEUK9Dat362nFCC3CQchA5UwidGUmn9Vom0WEwy2Q
iFrvrPujJo2Xh/2Pg7EhYU5p7Y88ALUnyhziFMJF+O70DGD7a3YMuUObA4ZaI7Dc
aQCLlsAMC9tqRLbX5C6jX/57gHcq4tiHdxwzGVhAAkEezQEFOKUskWFdptvifM5V
Db0LKxXLs+chuChBwCPeIe37BPOpAm69X8k3wZgXSIWur3RpRSvNfjeV9ilLf4ug
ux38g6h+SBQip2bm23lNozC9KgRVjSCyS1bk04fRPj7/u0AI1eU73cfIYkdKpicT
a6+n7CCLucek8WrBNh2Ma6FleNpXA0iJWud7VBD7b491K+p5LmEJpyCanTfrEK/Q
5FFZ5e3moTxaMbZf7b0S4I4Qdo3dUFWNTmx/LZdOArQ47RJYVwKPO58exfUqfwcA
xWvT3h2THNKfUgQ1wV+LRW7/ebdZyxvb0t3j9NuZ1cXrkiWkK8sMkk6RAHQ9GQhu
3hiXtIt3/5gD3GXrrEofBd7qx92lUXY1E/IucWhtm83E+edKelCMrAS+bG9XlBmO
YmkRB9IfQV5PtBs6Sa8CmhCQ36V1OpM7BAz440YkylGq7H/nFlaECQ781UNq9zAy
P6Y1trEwUyzPAz1GPTgjiAX1cvEfOkuMphAHamAFTYRkBHaceMOdXzYDgblgbPf6
Hj1oZNu4SPmSimbipb860ejA3oD0Qc4xzWQAQpHREtS5+XP4zz6eNZ1WKGIgVC59
VuI5z23dLR4h+TlIBPSqNtxQfVRrfYI75kysr8KPzIj8mdBSfFuJEI6S2RSO5Fl2
50HwUtCPiNsujx/v4klNV/yiUVeuB9c/xwIbydd1fXnZgx5O7aZ69vpomsayO7I7
IqXfZA7a+kao9T7ZWuQE9DfKzGsWHQY1mdJyMerpmayE+F19dMsHsFPjtBMcwi8Y
0HfWAl+K2klfmv+o75DGviSkcuLW0GtUeDbZKX+bz8nPoT6qJlExr3O0CvZvcKw+
wSDpQldVkieLLgzYlsEcvsTx5n7smpiewYI/+1Vh9FuHCXwfjAJYUX22WFut2zIp
DLNyNTUuwVEZPFy0lsTx/uEeoRkfhe8HxThER5FPJbsHhPIE9pwBXnrQk1uQjIMv
/xcnEobdt5gLtDWO5SrCw+Y+/z2stv0WvDw1N5BLpRis2iTgHTWLC9AeGA0aYH1u
eetACy8byjdvIeeNhRHUbVcJZzPCmoYw/rAsuxiQ3nVElU2eM7DWVL0vwc0btb4J
qIuzoDi4bQP/mYqtnN5bK1CJzAaX3O5Pghw6//0h+IexSaD1Z/AFBZMzwwg2HVIc
jBQK9Lj5j+xHDt+9NY3pdQncYmRi2bngAD8TSzmfDNPm/fDdXagm9t9U+AqQPHtV
t7nOpItYwOkmvW+WxUqzPHuzVGMksbOPrVTGUk5P+I59ZeOR4zxjEQPnXQQOdaMe
VbAEAsJhK4MvotRIshETY0j7qS8GI1XuVjdpmC+W25P44vEQR1f6VCeaLzKbAhlt
HfnBJVKZ6bSrAtPv814UVkfzd9acUqi0T1T9w1x35u2dnMRBFwfLg77ofi8XtJbr
vWx8ZJkMeOHE8H0VpzJvO6qLykNn9PNudTel2BhTugL06zQopOCG2P2zp5QXHzvR
B4hpLqvP+kHX/IHW8W1UxN0pl1x9lS5QFbb3Hm0F7uycGKMYrFiPY+qdz6dFrW3l
8y/zHLAQWigVlq+ipgj9YH/HOKObROygnO6lOu0TzuTOh8PfyAzNMWNTAN6zmk+R
nmviDxRYbIQY92NxJvmuvuYkJdW2LUY04M2y8x2WmA0/j00DQDl8vIvXmCzq3xq9
cQq5bAt6e8tmQ7SkLF1mzX+dsJe3SSPnwaMidpBElQ+cCyks1gALfvfo9gOZACPv
uCYTOVCj6o34zUO3X/DtukslwKrhJrtBl4fXIT514a36U2whk/4eVX0MOd/8aHpo
CzaWPqa1WIGtrSdmBZUH32Ob0bJFKNpmrQsrBueHfz/HyBIneFgygnVP8nE0Md44
9YvFv86R9Ko9hYvfE6gzJhuoqpXuocun0KYWg+w1f2y+op50NVEp6vYMcBXCFElm
Ec0fmK2oDVKY2iUauuP+wcmjZogFiabZF4fpIdBxPytqERZFkBIsFLAomolqP2QD
mHbLREokI23b4FFrXz/X4GXj8/PM4WtEogFccGYC7hi8Pa/LS3CZA1KVLRPVDrDn
2vKRwv8bfCoHDv+UVxbXjFLgbP1ibKWtNey5QGTpseZtolBmdRj5/1R5FS2Vwfxs
U/0mL1AFpc0jPtxT4aWZuFIUeAH2QiNN3/DvWySHlcgviSxoiU66zPNhP9yqikBY
Wf5IseHdDcFDPBCXkW60BVX3fxUAC7blgV6BAC9z/AxMfz2TNfK0g6+g77tS4FOh
YdW5rZPmfEz/QkE4GTs9juFnctiDbj1anZHdpVD8LNlJV0uVF/fQmR9QJY620jmp
XbmOeLXKthi10GZETyV+I+p5JNeen1VRIx3eawHf5u7xh/XZNCKxnNBMsszYI48e
bAyD349Vw0eOFGWAa9VMn/U8mQVNoZix12Oj9JQRp9u314q3Ojsq2NgT24ngOdKs
uktnNVi03NQhTJ2eVhtgPc3JZ0FcOMb6MyGho1mVoZf7u59n/Eg/EnG9kK9HDq1J
/Esvia+LPsujYpBQ1GPvbDVNgXyBlgJt8MbHrBBWBBHlsvrw57uEKmGdIef/9KZ3
sTnfJwAYzZX7aDT7dm7f+knWxoegO49WpHov2cYmEYEaI0+k8bdghhgyaxxSL76A
cWZ7y2eM4uEJxeeeBdVbQ/BIsL1l0P6eeczpm5SPvPrVv697CcE6/zldUud4eWqu
A5daaGuOGRU4i1tRkLyxeqhP2VXHURoi84IDV6wp251RCRxVuulZCjGsbc6vf58x
BGWHOOiAkZb6f14VCOEE+N1vgYt6QTaa6oVUMc/Pg/39Lcl/IARbopT4jMKPlZ+K
QGc4Y6pyIbpxQNI+i5pCHyLrzXjuMe0/efJbq1O3wuDTO3q0vWFtiSONQq09C/oH
dCZJQ8+UF0acJlytupglR9eXdwg8pI2XTZk/sPaK2kXN8GvxvtuOvcNsvyFIIMfI
/VPCd61jCYNd91REfrhWcyp0xuD8NZa9pWVT3Xn4fgsfc0GD99rXIPm+QhOKr5HH
Aux8m2mFUmHb7sKOcl5hQc08feHRNW0sx5nbd1lDTS44c66BPkMGXQkF7hSe4Ftu
lzxub8+/1hfS93w8gbLOIfJ/C+al7S1JMuxtukz7LNdIqvitILTsC2cIe6Ze5cre
sJ+NJfO5Lz+qsvxj2mcmKAZf/ez7MwFlnrIR/YBpfkAjoDq2sZ5WwjpFPLT1tu86
BAQCym7VDRge74rP7V/Ct9iYkqdntCkvkXMpbMLpnRBXjGz+UmMTAAlb4FSnx2NU
hdpVkziQ7qth5xXMLO8nDMO4N5QPl8ycwpa1iJxe7qsdV68iqoTj1FGfymW4X+M4
8s1LZypr1rYFY0LdnE2UCKQhy/7wGmsx1ESirxmH3UuGj4UJLAInS1Djq6hNb1mo
4bb4/tNyyyQYoPD9dGaY1o1l5E+Y3/s8ymnaXCZN8BYNZQ/XDR8eQV33QGa5nlT/
ZmtDXoa+/d+4Cus7BYmVuIhkrM9moGEvqelwEd3tgeHLVbB/RV9S4ZIOK/Hk6ev6
WQyKBEBmz8DO43WaJe3uoDur23SkLU5aiUnvb9BuN9AmQlr83jowUHtEqldSoFlT
gnY9FbwabcTCRJxCp2ktZ6jaMlO9SOgjs8d+OqkGJDxMcU5WNUmfGospr+r2LMmy
PBAYgDeXZdSpAba8QC5cL71e827ozpqwXrKGWxyPWX5SVhfAs0rYy/GyRRQAF2ph
gAeBPJkudMMMnwrx3vWTUFlAqh6nW0c0rz+qrpM38xH651fB9n3Nqm6wEUktbOXq
OKydgCQl8rykfbEeVVUspTLQsYLJtDEpHe8QOhTpS949rHz6o1O8FA1O6oEkv2OB
BMlLaOBSoVhgfxC21pZhCjbLiLiMBHdNWNWQzepeZpgRNnmJrlqX9//qY/oH/Yki
W7TOSy+REqF9nMNfHnYPyC6j+MqJfRDHy+mXB2l3qeUIm92cawgndIozNX0w5cNJ
78jqHQ6237OFSTKgFyY5W3BYUHwGhHtbG+7bQxp27cf2d5M+VtcfZ6JXxQ140xyC
hgOVsad245YtoGB9RTc38aD4Xqpy7cim2qkRH8UDGjog92uylEskQq+dtxLgJAR4
IU8b8hf/T388Qsa8XiiZC9DQov5jMCrZZacxT/noQiBk2SAeLwnkmfvu3HjXhnf7
s+SlOulZwIpeXCwT5yWzg3/pgiYM2OnMRDCG1MbWklDad3P299VxZTsTJvExcAOI
PuujJVO10re2wEsin6bC0BD7LRIikw6hIwmT9PLmLgw7VHh9w4bYD+XhkLppwAEU
xK9AF1JWppM3R6houNE5J7/aiF/pp16sZ4jk30TEL6wUCnv1Vq7Kh/U2XxVc5837
tGZnb3el4KNPQebbCYzMvPhvXAgZ4Kgv0hjjamIhyZGO3WmvGt+GOMDNUVAPa8nD
a8zZeFrDGfPiRAcfV4kKQ7g3d9JYG+oP6A4z6UUtxHfIUcbGReK3+/1qLi6HzwOf
93Lf+c/78nWl2UYPbx8Z11tnKTWTa7diuG5dI1TmtTS+3c/YhN/c6X3TWYPM3XOx
S2qq+eQq+bR3w10auL2n4gV5FXWh3v9IYkPZI4biwzpsWVaFzilKbR/tZzehOteo
mao5Q2RBoT4B2lJRJTwli5juPJPxIm9ghjcGe6kbzLCmEdCFOVV9G4Q7sRHEZTXr
YrqpylSOdwZZM1AJH4+0Dz8qxtU7Qlz32fXIZelO02U0RR2Pgr2FxM5f9iNr98Uo
m8CAHESM6U+lQCu1+Whmq7dLLtIKAn4kYHA3TQJ0zDsNJX8YcmhCzNlscTrQtbUF
3QVI1/gLw0UctyNh/3Z+AcULhAmouY4UyLxENZnWgMfIhM+J8giuk8bfO/d2HIaC
LwNIWrQetcAh8Fr/hnqxDRQRzZCZmBrW+LsrJ2DlYdfDqkPstfqHmkxEasQFUJBz
QYY8kav43KcB1llVz31gQHUR5E+n+cBr+sbU2L8F8ca0ZO6K2cWzMmlpvRqQ5x3/
K9Q1mV8W642aqY+Lrb0HImHpyZ43UAA7xVXP48Y0+K0sB7tQsfQGkzVb7QWtz2ya
chA4ULdFInXfpnGnbWGVJaZ2ESf2raRM9rEns6TfZt5qZkU6GGudTn7MDpHnu+s8
9sCPtVtfBf6iWqE39Xrl9MNcu5p2Z6YO/o9SQefFd85DcrmCeQxetj8NWhxck7/t
IpaqvoQ/fHaLc4m4yMlbAiZ38MAStUbN5eFDt20Mx9+WuayWqThlphhiY45Pzht6
hj1MIZCn32CoW7K8CT1EWQU8ff1gydblp5CwES5eetU97lvZlCWjym7vEfAUKSbM
TXZ+VOzl0f3OCoIDnnb/6SqntAj1TgtYWwI50J+OrLPEysqT7Lpj0Yrp71HT39wO
F6ylkmSVoqyCLSbs1IcAHsvCtkrXlbh4F5Z5XfW1aAkFeYaIV4q+Tejj1N/uaaIy
CWgpwlJj02JLrllZr2xjyA0kB+w2KtEa0+911oQpv5679+84PqZjf5LbrrBDsu+d
anAm0y/W5Hi4MeaWACR7qrNeyeRGyBG+yBpIr9+9tXn3E99PsKIUfCtb4igr0eAs
z1fZsiPTizIydG5zYxmTasn8CDBVvIdaNAFQPkpJzXLcno338iEoh1IQAMJ7aysJ
Z80pLYDuU2wpqkLb72seeO0rd8CLC+yBBJn3FDk4U19q+hLGNr3c0yRYggbOGaap
tJiOwmzbt/OnubTAk3les7XDxNet1vbNQSXaojavlILo0OGCobi79/nfo8IMWsZF
SC6G0TfUENH5TEZ9t8hRGfM93TbFxkspseISLxhLqkhrdCbz6CP45WwakT0tkyjW
Bb6B27c/J6Nbf+uIy6fnQyRXDGRwmR4p0F8f+gzCRh/2Pyu8wLvfd5MlZcOHPMFQ
KorQjxXzFti/pRiRSws7wIizCF8fsi1mIxxxbXurTPt2ynDmCEfnAdijW0sUMbXd
A+MjcfJcJtwA3KbtA2wfcos68fljxTJvPExoDaQAOFwJdrv0cjnI7Xze8hFu0m2e
BHlG7Xr5OrZeHBoVDFElYW5J2XbZujO9xsDs1Op936NFHDtRHI0vGtaPbkAJktOZ
onyOhbmm8UV/fl72gZSP2fDEKxlOdFbcp0Xu6/3sNe3XPRlwkg3wrtMrfB4wbHZq
lyByrZAB82QmotSrpm/abVS7LU6Q7WYuh4logdEYu9yvykXnSnMu32YhCBjfp/kL
BmxfXwiLDAm+sAaZ/NVdrUXzXfVJGO1bVTjwWWcD+DO5y0nWVpxd7PYoTSwwtbw+
lKLUj1PzOJzTGb6zpxZR/qsFQBzBbHvJvLD3ALXt4iPPOB/6LwD3GwS9VE2EA2fs
WDOLWAcpqS5dX8DYumbDY7/QKryR0kJX/TzvQ7GWnNjBPkqUylBe/0oMU7BcFMKZ
gGBjeR1dmFEaASrl8yw5I4i85IffneVXxpgzkLRslV/aZ0u0+shK58WndczSWADu
/3gtPMD0usAQfHzvJbyoKRXFo3NI308ykmuFFxWm7JrEuKqEZbxZNFoQyZxdeMtz
D6JzDy90HRQcDB2q+ZFEawhqddOX+IOvdX5ytLoi6YXvk4+cdzFUtOgOPPGILGUn
V+ELqoJPK0iKQK6iU+T6r1po65vbL/3+V1Z/9XWzENWqDWct/TvMCvBCtq2Klef2
sLynHaeLAZgw5yBJxMcOWfwOpMl6aVXQv8D0fovy/zATI+t3FiYkvFCnJad6cZvc
heOfBPxcAfIPkhlaqZtVpbVZLAsjiXPejL5E8fqbGX+rLe2xjvJCxNwZDvvrlU1g
qNCEooqlcTOO/1YK1N6Xf1m4AUM5ST0IoNMh89xwx9tI+rRMH3xNRVRO8cgk/mEA
E7HugEBhmohjqU2QapTzPyiaMwUOT7Guv3r9zjWro8BXOh3gEpkVZYQxDA/N8TcV
/D+uxKDURo/iCewJu/pgEEdWyXsw8mwEXV0MJSMeUzavquolsiNDwiR8i+9MgAuN
4wNTBjaI05z0xEesIywz+jtNoHmg0LNE/ysEqsc1qCU+zybhEu2ZWFINZycTyg99
TEastkpo+Zz+mINWieUQSui/y9NWwrKvY7lMko2VdXDza5M+emuVfn4t4FdO+WZJ
+WoasC9OZCC9WEc89WajLCQMqFZVV+/52R+gPPy4tvXHRMtHaVNVrp7Q4bvraXGy
FK/hrKwiTxptD5hf3Q2HD4lskxXzEsXlkKhSHtvJzkFsyd5wQ36JEaDYEqMwkBrG
siIq3n5DgjXEZown6Iy82+mtc0fnpox3qiC8XnkTxklikfjaCeTMZqtis5rY6ut3
zU8fTzj+jtX5gjojoYvDf5XIdGPXr0ykZ2ZxGKFH5Cz/X9PApCIDNVgSqrblQ2Sv
gSxJgXK44dGfv8FMlaNrAXUtKqYiryr4p15M8QLQzYsnbH1HqLmVwPcWR2D79Q2u
3grA8kZJsmh7KqPBWd4UAHLEFgUu5Bj2c80foCPVz3Ey8kKuxORVpFO7x5o0b9up
jKdgNSP4QKe5orVpMdb9KMlxcDfoOTvFyYnHB1gkXzD33egmuhOKeb+CdKrRRrs1
HCiT5XPDalTJv5XDE4JY6y5kZ0qIRo0WrB29xubZdykfUOP4od0XGyoMBDKBvkPB
/Xa2JSFxRkDGNrLJiv40/gFCLtwrUs8aWZeHFTS7fXm4GkYKwmz4mSfN/UU2IZIT
uaIfYusgoA1vc43ukyY7yeIbHhVvFhPymD0U3lML2uGw3fm1ZaWPME9asz6CKYJS
z7PJon2tqN/AUD/evOQheLDmO/2C+896wIjRzjm7bg0FOJVdnWQTDfCJv+YpSygb
OFyG0qKWLIeXhCvQe88En/hoZIblM/WADejPCiSf6cSOQ187ntUJFjzajWkqomwN
G8pgTXmO+SAGCRM/VpKsOH0XwC/G05ay61DlR6ME5SbXn5NCaq9UwsoKQISNkCfj
+2TA8Bou7DBJCUPz+ZOA0HvPB8k330gZ5PJkB3iLAzLr61vU4ySgUHPmH+3C4MS/
lyYRcQHBl1ggc91iqG/oJwC6UHnCWeSIUBWXkmhVtSj2o8vB8a0cOWuTi0lzB1Jw
MF8HsuQZZJskaWndfK09WLFEs+GZAFdeWOKcfJvD6CQKNwAK33bTvAbARsfipyan
LzcSmO3T5dx92pQRMXGqCcdqgZ/rUAiML9oTsgBItZU6oAHaohVpRH8vIX5nWi6y
ZaBSTjUe4j2hlR+KIpddVCq7xLMIiGt81fcTVwn/35guzCWJtlzU9T1fcPGtG1wg
pcA4pJ/P0fSNgjiEfPPDUdnfSzhQ3urmXRKAaY9J6QGLLr75HcsabmmVwcO4mZL+
uomci7XoYPmORcfa22uOa0M/xGHgvQ3RTwBr7lg/E+npld1eEgG0ZAQeDvbI5hJv
2JSeMtIELjHaMPA1qIm8AZkd/JyDMF72J8M6G+nt1/YD9BSb2YqHW762Vaex609a
/l34PU5Sg4/1rcC/h/PQlkwSpumrdQEu0e9gQVZ8EWLanbae3XB8wsAbbAgISp7d
Z2yVAyCCtCxYNAroxx4SK8e/kbKqak1VR+YkbFnYvN5Q5x2uh53E1EVgV9cTPUmQ
L3Cfch7jhTZT+oLk/G63ZhtupAGyXikhO3CFmnngFGqyUepy+EP+0/2jDRKCWICd
vxok92aqDwQ5c5atyCKU2Kvf4zk8PqcP5uND2vYTnUUVZQrCcP8rz7nTHY8RL6oU
jcpRTU+DOOFXSHFZxXr1QyORCPEHRUEJl6jnP06m39s8YolLS4otPUn68iN48iS9
8VNsMMywmNDVDhLS6KdOKQ/YvDvIFP0zgNmd7410weX0XUguTU/L/9oDfUgs/s8o
+03OkIlnRPSVXLjV6SYupenJyy00l2uPvXCL/YyUQ3oVSLQyDFJB984Y3Bx/pOMj
8/H5VNghbE2l5KHclu7TyQPZJL0PdxDyVk+a6k6DgjpnJIdhX5O+YCx0BOmWd4IH
O3J1ciiaph2Nqw5g3gNDQtWKXA4DCszxGnjD+SISP0HGnC4UAAmu6ff6oFSmfpDI
xNJxqZIakddVQKiNcgCGb4Jqqlolqq3+2jmyjKzsNnVs1bgkZSHjsXiiG2g0Ki5N
h9gPDxH0WoEeuwpqPbKkHMcxr7bcuYvfTZbZEFKDdH/wrtGL2iZYEHlu0XqICWHJ
4NlF2tR0/T3fOIbBHM5q4ifUYV4tWrkS1Va7kZYveJMVxGVVV5ChKei+k/2nypAy
RDCE+bOwRjwxPyWztLb5sl1ELzSEOjMf+8SnsIsxEijlmX/rqXdZ/bwiNTqKgxiK
st45TcfXCNA3v2itd5xC/gTOarmb7iCsaGTwd6Sqq5Gk/rIUHZVssgHma2tvtOat
RtvqRqagq4xUxpACbvw91hPy2TvB751j5QOgwhUOoGIOi89vieQ5S+SDK3iqCaB/
nUIeuRiG7gZqCdD775L3DOJ7iWtHNuOKuC5e8zPv2LVhc4yoa/I56TSyX76+QwSx
m/VrNIZlW3FRprlSXyiZFXqE/8ZLHYHDBKSYrD/z8ac+bT59975HJton2cDY5ji9
V+Pfc3cai8z+syiULqCjZXYR8z/UA4DXqBcpbSc5RDuV4uiY4LNfYhedZbjKFAtO
CYBGNzXQXQtEcNtaGz2Xjdq2qaotqojFnMrhFsEHTJLjJWoV/1Gl+1HyKg79Qky1
MmMQTukVzHPK59eFPLunAjAjbIGwr35EjzIWS7uFBtQ4KjZdFDuj9bZeljDiJzbs
RvtaVm+Ms1k/K+izblDlu+twiRvyo1OuXz6G5200eAqwyll/L9sHHzd0zR9z2M/9
GT0u0hm7U9/aVo1ASCmtDf4HbQbqJBalf/rK399E8IixJOe1C0B8tat6C/DGfqRn
IMvLZG1T/orrrMYnthM7oLOf8yYgroeQwA5OI9CkiC1+2HnzsfjxdjjChroBL5d4
W2Derct7qKMbHx2ed5/UkDb+fQzrEmWwgD8bIiLpqx2wQE5L6ptHNLYDUSxWlPdw
ktg6jJpjpCyh6+cEKWGHJum/ijnk9HtkF7jJEDf8cEoxijEik6QBBRIc4+VCQO2N
/2XFa6uOr+Jj3trONLHyskh14MPD1ivxE/UiZUY7GPeYh02LOMwE80HuNtaS9uUB
airkH8d4fiaITLQVZJXbgTiG1hEe4usQ9/r8ekjAX8YNcAAMBvYbxuTHFTC5ss3z
tfvRL8B13l96Etpd8nOUwcmoWNHVibhA0mvbhtt8SYFp8DpAybTppshd8L5pg+ym
F1l5lYsqUsoRVm8mMSibZWUpYvucDWAEGZ0G6gpwKFWo130S6hiLSgREVNVsdi1N
nK5V1mLZg7nReSrKRg3E49gwMLV4s1wzdT6NEMyxf0nG5pPO7BhUMyrS+0+ftzTm
S18svh6j9zDNLmHILOXFb6ZRMa9GBWMLVsYET90g75RaZJBmnAPLt+Lj+MwyarF1
S3XeNAd4We0J95hxXbrdiLQbnyVnf5+n6OiN1MTl56bpyGkUaMBxwppXBpQAh2+f
tsCl8hIz+A/GqCnJb+G8+fF2M3w8a84OiDcfpEU9SKrtm5SejQG+n1fYuEiP3NaF
p1j6LWgDPMyPf+8qjyxFYYPu5EWxlUAwNJsKwowcN95KSpymL477w+4idg3dih14
apScdOpuumqYJnWOxOgypyZK9shsntwF0qpHAxDK92zS1FCHaaz+Q+wPyVz00gsJ
7UPjQ6vOoccl7+WOscnr9V8TSZLFzh6tCol9CkRuUuXo0v7o7gboLPyfFdFN+xXH
8Dh7o6TTkLXOd7oDsFTmpy/4//+ns74OD/we6XbaSrvmuM2c/Cu+TR0v2PW9MEAV
hY8PSjb6s5lR3DH+gda2TWFKSFF2atFGcSkywmiMAWqcyTFmI9KKKUZrDoOS/HaD
hFP0kHJ/BrcxP5h69q90/tYgJBnJHFoqCyybHTtJme383QgF5jDTsfV40mPttCoh
MuLHM1jMGwpy/BSX5EVBcI3Hxd9beeuorocPyIvpVjdoUE1/mgm3QuDbeK9wveX3
v4W7HOrIMbo4MgsmnX2aeDv1sDCBXU+c/QrcWILJNGktxNYAbllxChzAzx98DL9C
D/S4RZH/RSTN+onoXXrh2yKzZwm/IRTngAfU1TmsUqN73S2uIhudUB//09l56ReQ
Z+sJUb6MBeaL1mVfZuaedmOeWMyrVBBHE8aMVP7OeFad+6WlvcDotcsipNr40VMc
GxDUub3EpQqKT+cx+Jbv/dAC8z/IhGdLR8zQWlOfisz59jlLWsHPSOqhHb1Hs9/E
4Z8+SwD6AmEayxQUZ9lvF7n+PpA9iMA0eXxaP1y8wx6HbYuypwbz41gNik0pPG0I
bg/7CUh5APd/H3gFWHiaNcpvyPO5J3hwTCR12aRL95Ds2vln+WpEMvJZGoHrZ+vn
lemx4GZ7Y7w0RiOuihxyZCUKogUhG6qmnCBrHN+r4dnc6AM/VNBMqpZHT8iuC4Tg
aFcoU+2FoltkcOCnzGfczA7t4+QE0nzcDOQZSuVGqn8ki3UB3z8hnNW5s2Fpepz2
dBAJxqyLo/zWDm1y24SeXDUEgpQLqC8KK1vBtRKdKrvgdPU/+AEU8I8Xt4gQKTzT
/PgvHOIYGl047pKOKYSomgHXrCk/W/4bdqv7dqF8I5W8k0NfUlBT6j0hQzNWPkBI
EhWE9auy2np/p3af9OQRbV+TFzr0kKSooS21sd4l/XuJeJqA1I7uC3Jg9qzViRiN
/O+Vjumpe5BJW6TjBt+8Eujxc8UuvoVn2VzSc6G/T7XASbP8RPQRHKbvwD28LAQW
wqt823oIXrISW/fZ2F6TPDIyh6jBEFvVZK/2/Rgyhn97AFNI+uVUtHB+d8TUQoFO
aH9w/agdtZWJWNzXOpVIjo/wwcXng4klnWXDmj9co8GhbNZTva6+3889IxQ9IUCP
spmJ4tJkVzZdZlR/BkjiHG6YNNfsmjxndyOqJ3XW4t1QkJtfgZsP41PMvhXOf7kD
IEQJcpHaS5QgGWcwBRtZAeHG9spi1y1PPt8y3AFqQtxZlEDSuQ8N0s2w9hF3uw55
Hqqm9jM1HWjeCp4fxsmVWiJ4/RRMTWxOgUjFaGnlUV3O5E4IvlVAygbT0A9sTYaC
NgJw329C1kfeeivIWfKcdW11/gP78bMaBZGdMnDCBFLEPcAibeodrIYUSYeF6O1C
NP3HTinuLwzegSrURRry7T1FURGjEkuIrE2l3bT82CDFJQ4n9fntlqgb8T4paLCw
UUaj+wKQwgx5+U+3Q2L/EKZN2BSILvlwGq923P9R9q1Hvg84RmWfOE2wwEZc2ZC4
NCNefV7f+O0LnsPXVjsspVj1VbCFxWuH4zVIP/kIlEgCz+WZ7OvMCR5FWxqzlztz
bt0lofGokkKw9Br4ub/d0vZLg3EJor16BtHj8esadhamBDGbRiKNdVCq5sHuyYGZ
mF2dfZsNuQd14wLBWNBY6F0CfP4HvptRKpwJdletGN37fGrPIBSzirS9alUjKMm2
Axb5BE6VH8JJmh6C/RH0Y2uPEdAZ6UOeKH1cYsl5TUxhRWRBvO2BHc1ysUXV+Orb
Sel2xwycIChluQrrYI+RfENFRqD7d3xfdBdYloVWyd/f4M3QVV643jodTA1xSewK
zYcdDSK4XRkxIJiQFFgi3RBgnR+E8ZiILoEHzkCNLWpEIf6+vQ+7XNjrd9JI4D3Q
2TU/bNuo044r+FMCPnhTPUjeunPsScre42wvdqxhPJIB+Ob9wlyOzz8muzhMqoMD
4WuH7PNYmEEqyhxXPaX8iBArkiibzaJhnwvmmh5uMHo+9gz6+uBHt/HrAIV2jhDX
kgs3dmjNCPawWcJY+tkQLYTFqFuEsJgcyQB+1GL46AmEjnQIpNyRIDCGQUJhzziV
krlIoYZWzlgyvFRPhEmfrPuoxLM6caItiSR3suMuBw8qimGQARmYUvx8Mrm5ZSQF
PdJxUeZ/Lx8l4gIvLtkiWg7ZCA4xXW6OP0Tb5/keI2PQ+Rjea/3txnjDHoTZd7TL
DkJ7K3ht7u9g8GJJ6FMKuqMAVKNoEkUhqLlFtEv+Og62n8ky4+ohZFD+BQ3ZHPHd
cZYTB5ixdHCSP+Bxofgf8MX4r2NzEsmyLEqpg9qeVMn+qewbEud7QuzXu3IrDxX2
rK8j0t9RIzk3Mt3G1wqrqQhRPJ4jfpyKD7ylCsCTjByzMllCitjYrJn9UuyBCZIs
RF7oShruyISqMdf2//Sl7bQiqNB1EtIAqYO+8P0xnZqaKBKhtZX2UgbdZ6fbmslW
/n4dkO0+e+AGG5G6D5+L+pdS1jmXo2BehV5M5P5k3SLcIB2w0x2MTpIClLuTCIVD
C2+/7eEbj2UjWrmlfjJihkah31AEgQU3qqQKWe/bXh3qKQhkbMdMY9z22ga7txVj
Sgw1k6yfRAI/eWu0YYHZKLppQQjq7x0HsAzCPbGcgL8WDt6omEE8TZZV+am+A8A9
D1tHeKv1ZMC1nM247e6v/COG0n0cPji+U3YMEYO9bIOCmkiENa3DkUL/w8KQ2PeX
8KHV2YLhYazPF4AjktI8D8euvPkXnpUdhVCrRGiesjwaXriTX02gkoTDln/Tzxhb
ZcWHnkuWdyW6DoVXCmMiwnSUg267pOyUBYUPsiT0B68CZ+aI2uKDJF8KduQf8j11
w4P1FKGZVqwtNXM5a7IEU7GXNH0wPr1Cd4yuttF48aKvGS8o/HJZeMhql96cloiu
v7U674PXmJ+1c+MKFpNjUJj6B7kbgMbfhA3hvdOgHsvSeju4goQU2ZpkDeI2RxbY
meKWg5Mtk/wOmzg5UOzxQu1X53EwBHUTvOH99bTMAuxjLZdetD5TIw9heVzApvql
Lp+urptbHHbeQHv5cRhG0HEyNtGF0j790uu3a/Qh6laFzPjSZ+lGePQ2lvy8jqnM
whXm0bDwIsSb1fCOxIrnyxclH7HLDVznJU8TAD078UX4KsnbPVhZ+Y/+Va821MtC
aT/PrYTgpVuRYRFKhLLkY0/ZU8NAHcUSMKPJdf7p3kGYHtFAygXeEO2KlQtuj0Bf
/ixLHz5WDI2oEyqIcler7IzbU588IUSIdu6wAuwBUrm3EtpuGXqKW4z7YE575eQe
UQpFJNJiOazK8Kfyhg/hpdz8qwE8Mp8MdZviBsHPX9tABSk9Lizmlztf3UGVIpuJ
rHlCcyc82wgxEDNpYQ+kaVEyFc4Xvn3nq1wjsrYc1LP9HgA22FsQmUU8tByibQfN
0JwKo7UTiuDcUWwm2Wh8n1qsk3mcxMYtWfUQuzny5pMgJLibQeJQIt0C8tHKtymw
OS3dvGj5TeYRakj925vpyMZmK/eMfXqNYww1Qkx8L67vh6u9N3XJeDLacS3jASLO
z88taDlGUnrD2xJ5861gGD+Tfx2h/nx0PJl6gN8iAZqvoWRMNAcIc68utIyOwpIe
oa6HYCrdv+Iecbwv4lV1TMLA69qDwJPCs8jP2BtMw69oOdjhJpWPBfCKJj9saMZd
cqYcTW9gblmRjg5Zz1drnep8NgBn1siiSE31FEgme3yt2Zv2/ADyL45lw/+G1p7J
EwtwJyNAjEkMG+ESHRUBMGNlbSnoiCvuieqhP6wT7ZT6JTl5ZOnvqYDEfpKqazMQ
J9wwJvDvitvihwWv1Tlc1D0cMfsry/xUXaZ+0fPhij8IzGjkgfdZIP1j07jha3X7
/4x3OMoDD+28LtN6nw8NRBlHzdZiNoUQ9jDf3XF4miY3RluVRlOQjmZiyuxT7Odu
dfVMWBelnoLCB8tOlvs/+ufYXT4sXrIZCi9HmL8XoeL/8rd9uGml2vWBb3JEet7A
qOEjQTQLISG5zQ8eE6WCZi/iUjno/7gj+Fqeb3uLYobWMJXkSKeOBLtoPbTRTX+8
sAE0NBUZ9Po1QySng4SahXTEMj3trE9LjIqaU9e5MEtMe+7jeQzuaydaYOrcjYEC
mCwFL5AGsfFmQKOcjAaXr+lbulytY8Kkx94awy4PTM6Olt+zBzqnXREyiAWuHRps
5J2ooJPB+XD9LUNFMdAq3pzEVsZp9daD1mZYSdkcJW7xpyHeB6bR9X2zxOb1fs2W
2l9WhgOYHhaToNWHlitnS/X6wuniXtb44NpGN+nmqWfynrY7rZNX1bjbs7WwCrjq
1RWJ0+HA7qEtOVyxDA48UXqyf1BTfU+992/7ntAwicdAqvhRnv0XD9tkVRbesfv6
wDLaaDNAemmL9UrEAi4n7SBGBgO0QoXPxqFDFIAVrKryFcvbKBrqLIKsI+qaz8rJ
QGDvNLqu9ohKc39cotyd4c1B4pF/iE03rF9Ms2Bhqa7wFjhck96AV/mqjoMZHzoV
lT5lwZtUFYMC9bu1oz18FCBhfxO559zjzE8lBN7MeNav8ZjHxp1y0LcgyiLXCt48
Eh7BYPyRrWaLj9jwSRQ7DNoLNeS1vEwI4xdrvh5VbPpsxShmeoVx0EARX+hLBFms
47ZQHIFAFyH6Wv/XO6F8lp6prJI4s8rDeeaBSXlAW8pT5y0crYaFQJiBf4n929Rx
SRVKUpTBLRjHrtBVvhWomQhv8DiHZ32roMIYSf0uCWY+X/6Iv2KQ929wgO3z1C2u
APHU6pG69xNspATZtOO1/gm3RwnViFnRpRyJhwvuP24dr9hmcreLwriMf2KFR/li
D/n/YF2p51l7yF7zv4zGvtLMn9AN8OU11ajwF5phnekTzUIo5+Lkwi3hM2HU3rrF
FziEIfbjUGjNrA5PbGMjPNDUmfM06KSe1arQQkvNUNnpA14VDg142j2EcU6wpNRf
4UB3k7JSx8Ng6Opg6p8WJsnDSZRW/AJ90ne73337iCl8STfTmJt5Qbw07qyzpxc2
vMizvfI9F4LC3nEsF7FPtnueHDlaqo+pA2l9LdUDfSYm0icUE1uFlRcWknVotOpW
vwrVarSJad8SuZE17ebHojNW7kmqpaO6XyDRkKUJ7k3fG/kcRto2sZO0DrImxgBo
fIpNJKo7e+50WSLsyuA2z5yWqMDm1+8pk3KmyVitl/kTenPiIsW1e5RoJ8wF6rx/
YABGAlVSGHERUYgM+p+NKxwCGpJaXf7B+ab6H1ird/X4vMkcL7dsdP9D1q34rMSy
BnIDQdEuElkyJiuTeeUKIOXncwtYHGMNcJwx6/gZ2GaeyxRdcxDiN0iJU/DKH5fv
HjzrBCiBcY+t5HWR2VkRkLG2WVpzdNotYNo4vWHclw+2ZAAuIty5OpwPUkqVZ80J
Xd57KO1EhSc3ml1hkas6pXz86gOJATXOgs+umAWJ7ayEH6QjdivQ87c1DRThUMvS
eHrBLxY9qdYSYSBsYn/2tF1JxD3l4wUw2LzxKzS40Bxa7IWIOAjoNZ8wFqVvDCGu
CLYg0wM633ZFVNIDoDwmVt/Zc9gypMFdx1nnrw/cizzxB/yLElsnLDS4Ri7R28TH
ZsR60WN0rWC6duxRXrE2jvqxfitZjCnxrqVGq+gHARqJ0AIpuvzL4TkkSZSqNPYN
y029kQ6xmNrKQA91A6REkaYROIuDI/KIJfL4PeVI57UKDsGS81ZYH0AienHXD97M
kVUyZkPmiTnrzUQXUhBpEu4gXguKcamFbgjswg5j61utJegoK+0npuL7KTmYE7Gl
fsYkhieT05yaA2kCmlcX/Y6/R7+BbBcUcedM99p65LFO0ixPHKJQtvk+xgeeNILZ
7xWeVmsCPTXE7oa/SKJX7vZxl86seeMk6kVGcoLSKK9smRmQdcPsuIRpkFn+Vuzt
6f1DYtguhcqHwLGbo4rncBh1lXqLEtJznP2k/6hsdNP0HIcQYc05y/1Lq5a7rs7D
C2i1DhWKOrLhjePdIdaO+X8KorpjVRcvCBPo+zncKypMBndRwDh0XzErDDGOUV2d
6wypeOElFJDdonXgxhxYMwJYy2Q8DfGTQyLUyDGMwuNTjvIuWy+sdR65fk2WO+4C
yoYcpZSg/E4gbVHatiJyo/UEhFfuUgwd+EYqLcy930iaiVCOxdaVR9Q8fdx6TpFb
VWQFGJ/rwSVnwZk3Vh91prsnrXDoFAQLr0DEHvesS+yoPqBQh8Hcm5soJ7xLJGDg
vLLTHvETddC5IfKqQuFrImlM1OnvjchFXIeCydORh5+LZ0T6ydumY0vkqY147rXe
PjE7Wwdjr+J/SadgQikuiGCrPdGHgjcbwMIqNBaVzk/QG3J8Kx5x6s0EG/C9BqH3
N/1TTsTc1lSTKhhDvPV8LlQ0t0gbvkh8CWWupU7xChRndQoOcBqZy+Frg/MiwTpI
MCdblEaIhmdpNj3Uiqrc98nUtC3KVEBZbXpEiyjVSXh6PAR62ZsyPdytsMITKQXN
w7TwSce9Xkzq7pgqqGTxgFYfPoSwOqfAb5za0VE3VamrVaimECzKdOKxSrMYpkHc
kUURd0t+cAGYSScs/KnjWvMiBCoFc1neA7AHdCy2N4KsEjHDjTUBqghmjVtWiYKi
KdLTlziBJUhRKg9QKZnvLJL0zF9JWneIrUjRe4ODWLm9uVUkRMoEvF+YalAKcmr3
C6kWRa7bX7UBmdw3ltsxBgnfSpHUvadri+2pzezSyJEIdNRmj0BX/sn7z8YfagrY
uEO1j9W4FjZ8UdzL4hV73+ZB/whyrwXTMkphw5cWrI9/aufL53uquE8vih0QjTB3
I1L5j+1YXUXjD1qyf++nZy5PkrLWeXOk8JYSjihctRt5nglljcz4fxtEG7M+0zjW
QzbuO0AXvyiio/g4B424T6MSQtYOLrPstO8ZwIa0cxxW9b12Er54lHAbfIA4D68x
sVoknLz4OLtZgF1HsPt+rluJxZNKFcdRqU04bu518q9Mdhjd6RTYrGAe7vnWMPJh
C/SDQBOsHixoNHT0UWpOrWGiSu7QYR0NNoYbuDlGaQLSKl7aXEC0KkujXkTBfYA0
fShuYdPvkkftt2aDHssnaNQGmxtYYwZP+aSTfAA+32SbHzN5GgxVCA9YNylKSkMW
73YSYG+ii140I4miADALUKUF1nT7J28A24iBYYX6/T9oSEtNrIYX1LNwASg7YKtb
KYKfMwKRTOzEpn+JEjvFI5C1AjDBLZf1muTap+bU1fmxhsr5w8fKMQYRPNuQcqqk
hOr616GDyCzHyPAHV12rTjSHswnn6jmg9t5Z2BLadROiQB9HjaeLjWeoYWqZgJAv
FhM4ZS1PiX39X5qeusD6gmq0/I16/0Ep9zA/SYvAM9NIk0yN1V19V5zK9zvIe6V8
TGmaO2LM6u6S8o7y7BF1lJd3oquv7wpH31DaZu/NDnyCfhDd1N3yBnSLZzIADfmT
C1I3ckYIaznNLQuza8czXSSvh9aStvERfPezbaBznVoqdVB+CteMWEdx6Pwp+qoG
+ane095Us6c0Swu9/n+ao/YfnNATdBQ1Tx6C7r6QF3Z3a7pu/wpYCMGnYF2Bse2/
fcTeKqvL9iRWceLAOLB4+n2xtMBT0ulFRqJMOYeJax+tMejxdjczTZJd5D2NXOyI
nWDrbGKO7HyWP3lQzF2pgzToBYXzUyOSaWwUtoC9Ccs5LH0IlQa27ZbxZPx+zsaR
ph286WGiAgsndJRQ2+t+q3bNG8bshNxoAh5z8MXqpBE0MQJZRQoVBnESWsdORV6G
e5lsO3cv5mMzWWcLWmnZ9YBdvd6SmJ2g8s0qG1+mclQ86ZHPUtu2sDa+lBcb8FbO
GgQaxmo6NH1By6W67Iybo+M4YVjfKoG6s9WSOMbF9X8/Z4WMYRXhRGTllGTl9qSO
PLx4u+QJ9JWCnGKzcvtPlZCS2gnTfyWxD9FaV/fzkQljsS9qwjPDJBhH+TXzQxUz
0DRbWY4wFrmOUiLtpZt1FbVdJDEWfaRmlNDxKrZyAZr+bXttjAlwpDcW+GpEsUMH
U/lDeJALvj+strWyze4mfbiUG786ByZV7M1pQ5RLE80q6EkjmUPB9nZRdqDCJbL7
XXt4lfqpkpr5Eo0LSQIg4cWYxfdqH+y7uSY0gdFa4trKJgnHOIyjMqADtYbdbwio
CKre4LhT7/BmUYGnk/uYiUn+kM+12S3Zb03aScGUX+QZGKJVHP/8hIj+xRGYgPXK
VJb7cd+HHFs13HlGi6dkKinCreIqOkhWQU0opTQ6N4G4S7UboPVIlmLZz3k4wrNU
WSMo8mOpz6PU7klv0Ajv2NdiABkFP7dFFK5LKb+4FUcfQ3knDtYIghCF7yRM6K65
LZ4GSn6iam8y5DXXCVHYe6moUMucR3dFX6zRJirzyP/3IFOkaN235zLqyfDamO6w
XxULHBLeiv+Hp3WpanKO1c4I8noQkdhkVgVEO2RX0nXzkTz7stUWZ5PV/EP87liQ
SPEO6QdG37LfFgCXjHZ6eKClkghgv3Fbxg5oDUMKjfzqLLpHMh/rizYABIrS85/m
Ldfnsv2+cQWcQzlJ7JGw5/BxKQTebG8ffZQ39FWg11KmxMMqI5x1bg590Vn5LGA7
aKxqvgBCbNHsheoGIX9zj02zsuNIUDNmyDUL3Wee83EXLTuiQnGdIugmzEvdSf9C
VlWLJyDFlI9c7d9EEinFF/xm61WyKg30Y+LsovaFUxVr7mXbXJ8trvXcWXfAnMzZ
dIYob/3AI1/cjbXIsBj/z/53rKt6UpP0SLbNfVWrOM6cDePKJiL7mMXyifuuS45w
Nu2XVs0T5ceVeGHwsFDUtwpNE06gpYc3cnP004dgGX5XDw0MkwzIiqQKXJkB/DqA
AORajyPm+oS6i46hNRIjOgoT1rSc37qugvdOZRdcDlELbTcbyhIzAV2XMbDDjRC+
6HvdHDjNt1PL8yVT7PHN1be4DGSeME30y/yuSSFsAhScdNobKU4YEiBLMzrhPpPS
5nN2LS9d8LefhceN/sbS5AjPKTa8xWofykJN//t7t7dg5XzOVxX4WwrmHv4NtnP7
KuFHtKPegAEXC+G0PU2hoUEa4MXJa1V4YctXiDO8TpgaVc13Gr70rYvVsfKRycBE
5GWHjRs3iaX8F7fZa10IgEaDWaSrMFGOdbmGZsLOCGaE6xRK341LqvU+xUrEZ7kj
sH9iD5QCvxw0cftPUR0ISWp5PnY83a8FTTIKKIIAvP8x6SwUibGWjlqXVj1yyx2Z
XiwBX779apOi4FuiSWtUlULr6Jfk1aEqV2plmFvvDv+FDq+rB9VnJIhBrkTVfham
D/JYPCvGjt6iBk1aOWR9tEfR1IcOftv6n52fwe+uCOuvUH7qSkMgB93frc+ev0hp
2J2SuYLCn3X4RxREOBIaHwqu85wvf9o7SSm1yBztU6fpapkyMWRXB3wcOWCjkwoL
VhRs/07V7BNeua1xDC+uHmGBSryU6NvyTRz3RbaVoJzk2iDf3L+I7DjeizIsQjPL
0JXEdQ+0TpwHByMZSW2MxxNM0PAMUkOn38vfgN/kb61TVrXNGtO0vRTxkcMH4R+Z
zTcDezlP/eAFRyt3OyWmze0IEfDpoUrhE27YORdNbihRjPPV5B0xPpP978SRXsB2
WwFy6AyZC4QxjRsGINPyJd/2z9o/UUIOAevmxQjx1SyI9KAKaEwUOd4/K1SlJccS
TLsvDEIFeNVY1+aysYtGNRb17FKSXS2rnFdYdwO6XCqnWToLkYUFQhI7CdANhz4N
OiApaY7TjOue0ocDpoifJ1vYBrwpTDTSls4xWp0/U60q9KJargaDyljVbH7FnmvM
39Dlwx5/XWh6yh3YYhhqkhVO1E3XJp0Z54fSPIHsxa8mAndPA47rAhS1Dg4bRn0B
lKLNidpJtf+j4M6DQGnJj4wS70sbVJXNoFT+WuPXpOAZiYcHE+/oAfCFzJ5LpQwX
i5AKCB4RNBQINDK4OLD2e0/Sw83KzKNkWNbvjpQnFT2pxujrBs4rIq1B97ptJ+ZG
seBZoHqViCs5QBBJCyTAfB8J2LFkLmkbfUwxqxI2Z3q6WOIO+Ymf9s8GWUMAdR0J
nDiXtXCcFOIRLFVm56VMORLYpVHS9/HRAWp9odAruJhXEB9pO2UL7Cx12DJEGruz
j30kFiOtrbefxKdEoQsUuWGueA6m7+yzd6J8Bdfz2qp8ln3togs3aVJRsyO66cId
FYlaQWwueevSx4ssvcYotiYXWDm0e7bgoEqCQuEUlJZ2FAHtF6NpLuhFnYnBQlrQ
AZONsbo5RnWg5Q1Ak+lVLe0vydmPnAflSvG3iZsle3y7TWETcJkW/IesMHUy8uiO
U7kIt1EfJNBZ9D5eBW12+WkvJIVHNgx06yzkeHLAgoWcGHz8cAU2ahpio4VkcM81
1/GlAtLPiEWEJ2zvURk2IVtbWkLXmg7x2meN9jBQVul7tu5mmVQfYpoUfofpMFlb
XK7OD2LNb5hI0F5OXXedgUT1/CIIbfGSO9svRza930e5FZbECyh5A0EXIYF1/NJG
EXP+YZiqCrQGhZoFuKqdoGOyC2cn4rewyhaMuILPxmsvjIg0t2EuY4Qd/FZC4VzW
2jvoAGPjJ7HbxjuEmOATg5qpuRk3wkyM5FDtvRKM0o2cu3CXV6RGdXoCD5dlynwW
/7fJiQVOuTz3lDk4R/TqCXGHTexs8YC7XaGcFBA7br64uCvj6KYq6vvG3JA2J/AH
oM8Vj61Ro6wf4B1+K53uBD+c37K+rF/dcCTOYbOpavKSWe7mESBZLKxHVzOTIbfU
xH69HZpMVkzjpxph0FSlqSu3NM2JndwBM8WMvw3cZScdrgd/JuvGyAfa1QpHwCIO
3d4muwiNGwiSU3wbVh2MRbPvHM7iuEt2vbMZuiBmFnC+PikAGL2goccinG5W2i+B
7ItC8Cspktls4YyBEbWxRntgYlrTH8t+8faPjqFbsBGkeSVCBIKZTWaH6aDTSX0H
FWiJNxWFo4px/9A1qwrvzFW4hjgEtJVlKYzNvi5KroNjqTbjx7M6OE47Ni1jgnZR
3pUmLI0GpEQxJLLJUw7iMq8UTLsgF+dLP27q+qGRBeeNYMiLqpoYDK7/QzrGtPdk
qTBebeHgs1OhA9tpW1qGmxaXIUwpanw2TwxSrkUF2Cvo5ctaeY70Xs4VUmvf6PAB
HU8rQnROq+PXPUL2SruPnnMhwgeGkYOXEnaim+h8BRoF0vktOGj737ndnw+tI3iy
xWhcqiZiZV9tEHycTlHbR28mjsMkXvuExM3s+aaOUNVfcr9R1YHDAQ/2tvf6TFnc
6kR4pPYYZpyQ5RE/FMvxDi83ocmGoQh53wgxZCLxF6ZlNEHwiCwznZcQGdrlf+IK
7atAn2qjSaiQBbE6HckGw9rp+Rvd5Fp88VGpnXn/OfsRLvrHJt0v33Z4PXAwQx1t
YrSzsXDsp4HO2R1BOw+KgjhCUubOK7wC0l3aecGyAQ45N0uMJz/ATRqzR+4B08tf
8nBEc7riUs1GdfFuChWmU/AJaFBzly4a3PxTB2C+H/X4ZggMkp5RwDgEKva1/VCF
LHu3w/LC53+Ymm4IJFC67Sx5zNBTXW5NCuyeqHyAjVwA/42sPTTB7nMX0RKUYfgx
EgxU+LX8WYlaLLqhfXdkOAHwQ5UeCIIDZAgQLiUdW+qhOg6LX10m491/LxoOdRvT
6LPWX3wSHBo8AnhNi+wG2qfJ1PNfI3p4kwwXXdLQG2oM75PJ+SJ0AJxFcgmL3ry3
bs0qI2GSO9qBrSibEs+Q/b7XzBR1awZpRLt/q7GEZcMcNu9rUDeTPlpziwq+wN4X
Gs6dneBPt6VX5mZWFpz8tT3sPM60kW1/nqNdTyPukhvG2YtoYoHj0Zo8nSXaQEX+
qlYuEz+0/OPFXAW81cK8V0Gm6Nu6ni8RWtwBVo8nHPrYl2arrRHR2jOaw6Zc1CVm
/3cTv+oodrb1/i9lZXbvw0NUBlVzB7Hfihp39Hq4/m0BLSvUmp+egkj6SZCw3ssS
os0ZKc6COdiUhSlhrwcx3oKv7mxz1LloQG7hGzVWWzmiLtgaET2yyPBcFUSE4+5F
fu96J/r+CTRjRbUtEkMNUDo4gQNh/iHANCqQh6yhl0VrgxYqALmde37S9Tce7yH9
+4+y4F2k8xCxrZCcg62A2zvVdVmBJemA9G+aqAYqywNp8jJCvtcw9Je86v3BTLg3
eLTm87s7CK7TfS6riP4k0I+1iDIAafw3cepEHP96dG/QguZuFU1UIODLVd50qkwn
TNesiOA362Hq19O0dA+FKcLhxOeNBrBB8k8qWArx5y3nhRxqDGvqY9BkcXmFoEgv
MCTd6oGYMwC8D4MululRE+TzRqmUjFXqCplEbkWYBZOe7QgkRQAHXEh+qcJY0gG4
x9P2s86Z2FFK1olq+l9Wp0JdmfF+yUQsJw4hSIQqRd+uowfMgeMegHbj23nKGuI2
DY4dmrMLG6zE6/P5ilVThFJNbhC8oaMoTeFncmcQhE5Bp5iS7qhFbw9go9sV9Z9r
YIMK+OfBE27YmYUaFPM93P7QB42H7E/ucInT068XRT1MJG/a2hT/bH4LTR6DK5Z0
C8G1dn114y+f5DpN6SGYlHV+oMeaZfj03d580qOqLriaCNBOO2wcsJVnU/7iB7iZ
cwGugIjnMpGyJlQydvjYfG+mP1dLcMPL2seQj5I4Si4T5ffaRMPsLRYvVeVPEzlA
LGoD+Biiv/bZzknH4OzPYy9qdiz8M6VIsrMvupe7xSSJOMZkv/vxk0Acc30QDGOc
yqvAyZdBJHuX6wcHy47Y2PxygJ7JGW987jaDpnuPiZFFGIKeCcftnA4de/1A4+Yl
F8oR2ngcwk8YfzapbUxxbpEjX2rgXO+6mYmDZjzCDJCshXv1F5C+cwyHRqyrnNoR
G54+cw80jhA2UBmGoiPe4jl6l2udDXxxqRKQ7IZJ6bYgN80sqPo1+JvjgR3mHpgY
SUlaXUnt1Qqgj2lQAfm0H9LjIXFuhuAGsh0jFVAmXNkPlh4eGVBgDf3qlVaWuio/
aN4h4jJw7OYirAg8YpxtiNHJvju7WY61fIBnAEaW+8ts2unbmya85Er4z4niegFp
5HrvKUhL6xKcKOrb2bxxRXFgr/+ZMC1qYnlTku0i0as6PjtKL7hQQf1OOdWn84VS
W4LRHzOLFHjH/YrVKHXMKAqURQsdg4HYgh8/FvQ/nA70009dO80dWSInNPiopIVg
3bhelaBLb/tuAeZQFtEafAxIXb/Jo6DO1zUiFz8ztUGUf8MjHMMLyxS6nPc5N/sl
zJfL2Xc5GhIUTwGMIooptDltxOmw3jnfzaIvCGrf9fdkeQMuHYiBRAd9udqegFWE
iQzNPBMinzXLgao0z1Ji/TTh8jrlLtChv6OANjBTtniaMnuNJZziOSqB9+Cl2GtN
s23YZf3qsCfp+2Sx0Y4HrkH0nHIwNdJ7YPbF8SUlyBtz6/83lpSevd6POvV2Du/F
uOmy9/TqG7YTMzEOki0FgfyJTpclhCQ3vImkC1D7KUT7xxArK5t7A5UCnkIMpK9x
r9ElMszNwVMEY3lfHZp28+lyD+Ws2lK/QW2BSwpM5Z4f3Wm+SFArXNF/8zEcodV7
2L4Td4sHVMhbE2kxHonVNcA+2rr4+xSglokyK7vcA7I/ahkkiuBMHriPfySXeUrh
VlWqClm/Wh49Andfx6WfkIXn1UpQRgQXk9U2YdX7eVnmXsJ9g3goDoLqNnEpgPsz
aQQKT/Ik4A6CriiYWVfH+B9MQkyXeJh0Qzlcru77AvJihZXnzslZCpCv3R0uJk6W
2HsRMab2gIR1vdsyMqgdzCGFHh9W1IainxMKamQCne+3ZDnKMOdQOb1dsuJMdji8
ZmFzB2oBU+OdaMqRg6aRPdRGDMbAMIMnOTHkht+m3g8u8Bo7AbOnR3zbD623fQHL
LJFfH3rCOyENnFJRnBNoV1vr1zvRqZYofwKabafe9U/dvbhek8PiuSaZdSOf1TFF
uFVaz1w7jAiFALGm18p0BkbxbEQSfvvmQSTFhA6VQRcyyEN5zTmOGTdDr/qI2w4w
HbcHrLmFqmcq6Q4HRFsSOVXGNiIFJ3iSwRuWvwGK0zw9PP4rUve2hud6FsuriZOS
/U+8KniQUPTK+ZDVMFjZKfyA/6XZ85XTLp2z616Yzra/l5oHD4IGDzWt0DAvOqJg
duP//w5WgZ7EeC4+PVjvbve7+SIyniXrJ/QIa9kgOGnitbg33mV8x2R6Z+gR5W/Z
A4bFvdi9z2u6lctvddq5ZQCL+rk9cZ2i3dxONBlvX5MW32BbqboC9q3WqXsusA8y
KQ08I+3YwredUAn4OQ3cVrx2MW2R8qGCg8TsqcDtoNJyrpjS3olXUSX2O2NMgtLJ
Y/btKo8VpsukSLV6EXAPzvok3FPzUNF6pi8APXR0+JZ+vy8XkRlAeoQgF6fdDU3P
NZenvqlpj9UMuY042b4KFZK9zUqQBd+6xzGlSAjsBSb7OAHt8hcMdNwpThGKlQ1S
sM6nN67N/OfKaHi6YsZbu0cl2TCxaUt1x4tOMF5riMCOBTp7Ymd4nyF2qdIbjIlk
5eUVqHlSTA1llnGizKl89vXflJyaWXdXa+cHkzYkH2vWONxURySEKqrUzMU8DXNR
21d7pNCK30QC0BipYG2rfC0E5x7Kuwmc9kXapHOSXu0K/S3DcXwh/V/WtxzGDaYO
zlUmKdnjqs+g3LOaK0zlD6lT1wDko4CEepxKwfeTKxV68uoBZ1x10VoxOjzakNLB
M6WaLOBQKpAsPvOyn4D61YYnPRZNrmICh2zbEh30Lfeoa9Tq0a1OyRa8uJvwcZ1p
v+q8GORTXZTI/fy/VoHMp4o0FfVnV28+vQJt4QSCtANRZynJJz8bBxj0A/4wOCLl
oo6UkG6ih0DFufW1bkxYIgDj3qW2E1bl9fwp8pvIHK7Q+WbsPva2ERJSuqqYbJsN
tMqYUmubmKgZa6zgeUjkni3S8AE14zSuUShs9YlCeLFuacE6ZK5aylJlo2QHc5lJ
gFQFEOpaele4BToB2XeZ3T/XVV5nbKAZmLsIcInx4icJLHPIh7uoXCedkmbnA+Oo
eqz3xb+r14yqU90+yk8IYKl7DE91H2+pKcq8KnEKhTW7yNKqJYy6VVssNNSURwo3
te0MaZIIqV4uMrRXOsNtUMGe4P/HKcDYvqG0ClDzgY/U5/KyPcCoNjIab1hqhQvJ
7vzsIzJyFF193huaoEKi7dqWLE2XADJbetBrNG9AS8RHvm+jGbGMHgm4/Tv9+0r2
GbyKHxhqRiDRpqxY4WnKjKyOIa6+ihIKL4awZ23dkn6ejlEIR+XspbJkzGO0L/xo
0iV7RukRUgDaZxuegcFZTJO4KENO2HVwYvxBawictRYfm5T/4mhujjRuWAco75El
2039gOxNjYYr4mfqCGrzM6DzfiMhY8l5piWDUSt1P6KIHmTfOsz3dC3Pu6vv3kVg
Xmme56bOa7KpqTab/mY7M33XpstBytsGKCswXMF8G02+OO1iq8tdarvaG3m4US98
WR1lHDQVpOFdkgKfHJLr0ORoIkSdrcGaup8v0rB8ja1crYr9X1tWk3DOwtOgkNDA
/c/VvK50hPqErWbvHLErn9mR4nO732dXXqWw2ReXf+gT5KhCF0BH0raXhUrtT2R2
8+u+A8gz99PMtmR26gcPRZMXBNWkjRazI809XkbrnYY/vhGkTshRYubYfQCRjptS
Rcb8ZR3lBEM+6sVhqT2lSCILb/nG3zPcDFOj8/Z+NB7raD59Swbaf1NJTKuUj8w/
LwAtC1GbqcDwJ265UsnpaXCeRhQBoMRfAWfqdJVPmtqYogxVLFkXFBadn/2NujZ1
gcXbHFvOUfxI3jwnG0HtsXvY2U9fvHuSGBAlzQYpvvckLmS56PwhzKl4RVoBM55t
C5gjMX+C9ujVxMHVrQVvztOgn09jclN9XT0It809WoiZqo5kJ9BUJjY3PVgaprtD
Q43WrhZGGz5QqAJKTOT2EOR9NOnSLQueRUVZ4iU9OE0vMWHoZ2kopwwTVD5D0t/i
QLCXkWZJJkIdNg3wa6EL+octloN5CmWN528arlMjfbYhHDUVcSOZF8rGjGycDEjP
7dI0p3P8UDoUavVO6xYb4QFBrguD+4L/gZPUi6WVKOIr3HwNuHFIAoUR5xve2h9s
dellacUyMBG5OB6GK4ew9seFzPjFYJA1PieLnM1RkXyzLeWMqvCKjjZh6RwpmkFx
Za+l8AVp9xDnvn+SibNRoSA5feXrrLKRGoQZcD/11dRB1hy51Tg8Meblae4B+VfV
/cfvoAqc2JowDwvc7ZfB8PCv+sCP8oWX6ZT+RoWoVXJ/gGAXCMWM4EN2T5edWzaG
UGZAfHBCH8DcCJjWwtapIB7TsaUJClOsC8jT85EQBSyXOhXHlFiecQErOfEGShtN
5GmxMVmQYgGgY0Z4UwE0MuTUQUUQMH1nM2gjgkjBDRioet8mzbVIFGgV4N+Na+kv
tvMNsNoTs6St1aIL9b8gFBAv93z/4F+rwCRn8unduTA/9U9BcGUcd5Ba4p0oquKR
Xd35d0HyE0Li7gxbCDA14IbgE/4Q4Zo+HoQh5UkuCad5zNUMW5GdCJR4Q+0pXiP7
r7ZVKze1ENKkeDATADgBnfYA0NoMkAJvOgdGyxC2uvKZlboGWPowdgPiuZsRM+f3
rocP+qKZBipmEAPk+NfA0RC04kl3cXJZP9Vrr6Nl+wq9U0g50WKKI2W/Dot6LYE5
Ug36vpetf78Y4Zz8xXRtmWLoMWG1KEujR3q3go6MvXNrglDqgprX+z5NepIvLlwF
8SxRmgTov0ffgddzSGADYmftSlqU9bUfVf30NvOJ0KRCv9WyuW/imTiS2lMQ4I5+
y6ejD/8cMMD0OsLsE9zo9z17hPpRU7KF5u5TSSnkPoEbo2LYumW1WAEvv4mVmvxi
KvRzH0UPYQI95iCctUwIKZToN71s5x1yjV4UMXGpP3DP/Jm75ikBIx5/fUzW7nrW
qrRiy/PXmCBXqIe+Ni8OvR+noliTvsI8C1v6VVb8MrqCgLxTb1H93TW/bjgID/bt
c2O01GG1yN8LSM6rMx7kpVaWRFxqZ7DLAQAJG6V/r8NwA8aSM2lWv/IRQB3g82q3
0+CHLTmxjZG+pODIdrb6jdcec6VYLkbZLwAsUbtds7nLcqJgkmvkHu4sFdNiqoqL
ZZlSOhNfpX4dBTThnwOh/d8hDbcJxtRezmZWKuuMtz5Ii8l+Gs9y8p0FwZNnAHhs
ApNivrX80uuLWyhKlHXWG7+ORF8iObxc62NFsbSOZ0kj+FUEKvbGCKTM1dRmV9Zx
tVC6VVTh6GOXJXTaHBzFIjnol+CUVl0IoV/q66i2SuySgq/9Vwx/E3JYD7OAIOHT
1Hg5rk7QRcwjsfX7CoFHKGIiQaRgTGn5l9lZ283XLnTpSY09jHsaP5kmcPLnsIuL
P76y49AciM+L8YKTxFDURD0ZWiWP+SiWmJAAAEra/nTg1juQOBw5AyO2DrncU4Vh
Kk9Pw4J6Qg9zyE+6F4TW96Nj5WvlA7lbLuVkogAS6RlO6yETkOQ/eAJQyNYdk3+r
VFrT6mDzYuzMR5Db52GUiA1pVebsXXt4EWZYLXUXhMEf7ig6UVKj7V+bgJYDu3Vh
NXrgkwqjkRCE538IPC2VtQwuREp2zK6oRsFgo0v58B5iRQ3XF2BgmIR//kESGVeA
rAiT/Vj2GeYjgAMf2Z7tWSjvOB06+e3dx9YuRo7m/TN1+v+7ZGot3vNyIOP2rkyl
yb+ThHQawCrJD6zxuHlR3fQSzEsi+6pwq5Z2YAfbcv7FI9PDo4o7amuYAaqgtEAA
RTUPH+dI63v06qgkn894lYbdghCP09zJE0wuTuFEno3U1H33X4tnDL3Jwyleuuly
adSn2lrlVNUlvyyIME8Ey5fEbxCZ0I9jATIYF3svUyYKQoopswbRYk1djzO48vfr
OvddSGP1veXFkjEsAhTPijRQxlLZTP0TN4KCAGkLhM01NJNlWo+O2JCuNTRzRa2f
WjxisMg1BX1xZnpYE0sW/Et/bfI9r+wiqqw1x38NtzySCw5Z4DRPrQaD/hHSv33T
H/l13VkXNviNgI7Hb0YJZr3P07TMGSyoBatxakXdMLTxgor6y6VxWxs4vgsh57Yn
UyfvPLaFnQKnadEyabBxo6Zgo0BdwacbSf7cP3OCg5BeB8WvJn9yozWc+kh+bI3p
ofuBtuuz6JilOvtyT19WjAyf5qFi5PqeJjmGKI7tiNDsUFzIy2XtzRt1SdUWhqD+
fLvARKU4/FXAp1jr1P8FpCBZskQyhDhilJ8SBblTaccR3Vly/O8tnYED8qAa9e0f
KBSOPUPX3e+vfhW9Dz4s2l/tTO/KvjqmmocCsGXKxMXbIzRqRqgcpYHulEHxq/U3
lYBg52XJvdEsSoaonFC2+3jSI0LRsB0H6MzIP87SrIrPoQheCR0bRV1WXgg9EArL
ulnzuJtrmL0/FvwfIyalLKJmIqLKrbv2HJ/xjdPD8omsl86DEhhZxO/mn2ffJY30
lVckO9+Mz4W0RT4kNRK7fjLvhrs10oAZGpOUu/vShN9HAsJ4Vw2e31rSDq+gB4aN
WeDnjnrHxqX7U8FwLQYlzWf34WrTTo1Io73hDEY39VVN+PPWdudSW3YDVTe7TTWl
TwMefAM1kwYx44V2VOSfVsilM9WHx0TnOFp209mm7b3aQ3IE/IZkWDGdO0wj02OU
LDDo8OZ9q8cTmZs/j7iCFL+sx/QGgv1pusc6BJmYBKZ6zi6AgYL1j8FbbutFsW5p
ZEsREnH0Gu8CBMvd3ZuVrJjw73LPZVH4rg24BrDFLjjTVWqgXr2yAggTSXPtVcuT
Z77bI71+JY0Pozw5tf37EiPwtnSl4l0KxYVpJxF0phyMU1/NEf/Xv22FFsZz3OKE
sAANbxjinPqwUFCmA1nmF51nbz6KRgBKPSvILe20NrCgLfiz/9b7g9hsrDtE9TfJ
p8YB215bCgV3UxkP8GiE0lKVz5wU1W2SWxaCbnTUbBSEOOIja9+Qchoqb0IoG4Iq
ftK+Z81wdsQ7TKR0YDcKAAWiMCUofD+wzurMaFeX/y9eXJUHVANFzsZN1WfRPzqe
imRDge2b5RBhcMQQP53u6IA0XWly1ryVbuYy4ko2tlyQV7FttBC+qVVsntjPNLK1
ScMc7Cp7gd6yi15xoeQDo4oP/pka02QVu3QQXd4hDtf/sYQJGumjAuxxSsnWyCxI
5Mns6BsbCOvUjGmsDKzM32TZCnO7fth6l9TUGPtDgfQoJHGZOxLnFAKY/5yt+UWt
Hs/pBRaKiNV1dc/MdYjiOQ9qweCIWew9u5LTdDdmFXJdDJqwBMVg1RzycXFZ/jMt
55A1JlZGoXH/RKm3ysZQMGEvAiO7glSZi2F+ZT+YRZy/Y5bqYSeeukMWYI+wLnqx
YgibOQzRbGQ6bd0346K/dIqrnyHn1Yj4QF2x9MJv3PU0y5ET83ZSrZWcC1NxK+3i
uiSzPUJQinmLse6VsssLcUrmYliX+oBFqI7ApZge0ETSYSHy1LJnSaj9FfUJRcAG
mtVDc95RVF8w4yD8dxKNLO6jnhlpfPEK3hzrqjZ2nOJHEc/gsch2z4ocVU6tVkZD
vjKJU2qshIxtuKBbN29FdhVuPDG1BbmNL2OuojzN8Iq7u/iyTAseAS5qonPRp0qU
nxN+7qoiF+uyLOlke4tayw==
`protect end_protected