`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 2576 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/9huKRhRMtvnNqb3Z+UU7TahEoHV+T8U3P3ufru7l1O
3DlgtZzb9QxCbOjthp9+wDkjygH0eUfDrEl1ovhZG63TmYA4cML/ohB6II7ZpUq+
u79oPSJLNTzGJbphhq14nQUVUb3sWLTJslCZ5yTjIjysn5A/MCaEp57bQKda/dt6
X5LJJjX8gVdl1sxTYdGy202Z8Lw5EX4pqjlAb5wiETn4k9SA9G+7mvOCeRyBNkO+
fGNey/kr+uAZBlfvC+4RZd1ipHoZcTDwEjAzM8MGLMy7TbyiJTvn8h2u4JwCGbW9
90rYRxukIO/0DEvTQ5XbJ4PdZZvLC9nUarSaB7Qlf0/XZ8PKh3lpgUc5TZIq2yPl
KF2QfU3bAurw9Qe0LvGxO19yofOgLFHYglwGUNqGTLzfb6HsDJddDMNYmpr0lHXN
hVgblSZtsDNEbH+BxQSQThv52BXXpcUef3ueiGuk6gEaN2ixdFIzHU7RWUzwVbMB
BNgAoqOED41/Pk3UPrkrPeIQxhrUm7LJgYwlnEi6c3YMp9MNEacL80n/v7QeRA+C
/akDubW9zyF0tTwTWB4HXpKQPx1a2+vv5FBGnjvi8i02CkBsD2CyVRX+i4inDXer
UvANXuhYaVr0cn+V9hGoJB6DC70ffmGxZjhhwW1M+g8hYbrXcN3AN+bjU+rK4qBT
seewOCfiWfA+L7e04B1C53ozy7N/ljtgDMqwcTMHHy97/tSbIzOWQB6otcLbt50N
lMkJGpV7DFXY33fOT1RZH0ax13rYpHRXKxZfgMtzE+auoLDIkRobKfZwZemK0yGe
q5YZ5k26Rk60bKZcnjLtYkB3JLeJpKZCWRC4tbn2OBW0gsdwdRI/G+NEQ/pwp8f0
ZkezT/pLfzAeZPkQXYabXcXo1dlokxQeVW18lLMxhabG4/xwbetS1vSrKrWx59tn
pdJdVeHmEINq92Nzi0yY+RBMwALSWt8tUSYDGOIEtU5Nwbuv7N7m+lh3I+ofzQqP
MaduIcQaYTvut5tFKu5lyt1T0Jt+dfMp2QMTH4ZYvvQ8RF7gAAINS4xx+jV3kcjT
wM8weeUmtAwzioVrMMZisf0cZkdAgmoFKvtmyIqon6I0wLcpiyCiBbYl9Xna9eY2
arcMKyx1+vbEHkr+MWcM5aRBTcankKYb7Odu6Grw45vVUCvp2Ig+ekumSfV6ZqHv
JRQQhWRTReGDL8wcmC4TpyH8NrUlXaQ3fpFwMdkcVmpA+bwJGzhI86vcfQHzRH1K
k7Z9tRxgXk4nMZwQ6V1kBBYVcnqf6In/xyTQ/SOG11OjGtEG8uEq/5Qy47rYAKs4
tvpaGrQRhOGaaOofdFOmUdrBNHVbwTwoTGwJdxsr6+aaZ2lZlnBpODFBb2kWjTIv
ES2Wx0Qu1ouaOEBgKrCpR8zPMYSHLloocZPoOO612zykRZ+Ku9S8zgV5ZTI3WRfH
bVTq5NGgsT5gURtsCx33CYfSPcOHbu1lKBePeTDjuZsn/xov+NAdgDtyK401o1PG
iDxGXFMquJKckIXB/jjqI/HdjWAR/5NkDptQOPSJBXP1f9Y3nTSHgf3I5mxiW/xU
P/A3CUWHOANFZxPBgsU+X5mlVxN66S1wRUX3wkjdcYpsmsfe4N/0KaVqihzyT815
xrGmBdfsWKHV3toIhuB9ODOa1HSOn1O9FxZ9el9F+eqXcEw6cBdmy0Q7EdQf7lFr
saIwpuOtHpnvKpcN5W9qPPTHQVu+Kfe3XADeb+HcfQ6TFgOrFBkeLgCeb+RNdjzi
EebpvVC0NlzFwMi74Z5xr0kI8OYIfaGeK0EFmPjgYjYv8aKBQ8wOb1s/cSuIgaS+
WG/JnItNXnHL0DTkYh9J88h6rnNeyJotZrwchbmzosQAxtylyxaTqJWh8+ANWvQ7
csuBkExfrhcB/Mt5Dk4XTyPeWt7OhATQrptHbah0SZLl1ZV35ipC4fSCACj/TEhd
8nC0B3C0951QWwOpX1Sf/pu0zijv+xcBxDxdB7JTKUH0EVeMSDyN4OR8U8LNR/Pm
qQOmwDekeyIzwlIHY4zlJj4BC9a62HMcUx9GBzHwsitbknRWrNguJWX9ORefC/TX
5xcH29Ecq/sA3i/7m0D2edIpiBF8ZrKZ2iWfvZ+7WgwFtmF82xPxkrCuac/+J7Ih
E1DqQhXP85VvUFIrz7PIPqSvkOSL/S3BZfiHTnANLhwgqfYPkGEIu1OPQWf2Z/ie
2TzFRaAa6y9n5dlOV5YeIXXBPFMJpZty3MJywYUyp3ERRknCi1Wy5SXOfcmWOBU6
p9lzKwFFVqhzkNr/5vXogekc4jHmlkiXNlH3lpvU9EJwftqzJ2xsPtaPUIGB/Dmo
kkPrssOmAQjJKdDxPP8DOzgum2NL6rPMREQERVGrDj00tpevuklBbitAE16ByKYb
QH5LXigyKfH+4JTG9kTIy2pQPI/bZBbycMm3lYV4ZzrorEwGo9gY4/7OPsZS0hFR
PysaAgS2DeJr/QM54+Uyo+o5n+nNpyGrd/VJPIX6BI04MIQLO+t/frkXvJsF+vl+
55n3FOttlPBabA+hfe6PRTysoH+WZvN/5EPTeu6Y3RuhTaBz8+45FZoJbU1IdGLe
APPq76EKCKv7ahzO6I9fB0zr6ZYiP83dgBv9hlu5Ngks9xN7DuVQ+NKiw6brf9fj
+gNiTl3TXpZXvmU1aP88Syxp6BmeF6WbH9pDRe1zpAJUI3lQd9QGcDbxObaW4ZMz
tUXhBFYU64H7csX8qoKFUP/6bl5HtxRlePIfuIF7rsZBf5Y8cNGJGc9RHQhyL18E
h479ffy4Ktc3jWnZy3RE9CQ4s+u9J+nPjxKddyCdcs2pjkvu8LcwsPYDHrXgfsbQ
MzFEos4+gqZor+BlJe5xhRUZIFmj2U0GicPBjRUD4/9Fo/BQ8wFfJnEAp5WNC3dG
bJ75ruy7ietiZaSFQ+HDzrQrso4TwHb0BcSk6Bc2bpGAp9RIY9XdlvMkc0VdXHRR
Nvg6fvqVL0zlFr2oP0Ac+54fDAOM7WzvqgIEu4NPWSay1Hpdf5fnyWZPpHamlyjA
FwStQ0rvVkcIaLqEdq8Jbr+xCVaWA5fP7gJFnca3fn3XZCZrQyGwPGKExIuBo6lY
ztoweoZ1TYLCEwjzELh1uAWfTYyzcksup3s6ydXfPcdATp/MoVbGRKLf++usVql9
ZP0PLZy9JTR+x139ns9tzBiwj3iY6MKbE8vszayekXQY2LDsosfpzr9MrMr57ehL
1jIO9bFCoEQVo2mxFOFAnC4hqGDUyedGeVyreONr/ySPx1xxhtBTVVNdnZEko/Ag
YDki43SBqttT9uZ7tg2x6Q8CYBsJnDvgThktM+yhgQ/obmegZy+8F93TM1n0TRYt
/3GhYllF3qDL3L8/zYFgSCCrI0zUMKX6GnJ8/1ZjKog=
`protect end_protected