`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
C322AjKOEq+k94hkAB74AtR+hRiX5ltWnE558kk+r2+AeJwVSXNa1+pFYfFasfHb+KckKbhZdLwS
fW8S02TnYQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ofzbFY7L06zQH12UEp8T9MQk32MkmgyM1pxnYEaMMkxVZT7qmkPcrHlezwtxvz50P7J+krNjLBvl
9WnXn7/AVK2e1kkdihNcD/4z+pWtcGzBZGGpjSR4cYoy264j4wSVdvBpkGSKWThPWbv7c/mnbW9A
FtDAWg+dMdA9gA8q5xU=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
IXMd9uE8RWu+CeYY914H5fGrv6wBgSGy7PE72qSrhvha977IgXL47aVz8iDNHhB7cPWaysiOfWe1
z44Ah2oDxeU9N/ACt4VELUAKFR66gxVBnP821bIV6lnEuGuDJl3Jt6TLksKBst+9iGTzA1Xbu8uw
awvd+dRvRdNaa6kB2gp1KE1bAYqbNMgDqNruZkGtFniASJW3xoeV1/4MY6Ke/rzlIV7+JMoBT0tI
DVQ7gnZUfCWyhBVbusKBJ6+UH1IGvBq18CzC6sx2IxEAvVuGRv5jTaSOssqFhs+hQyG9sUprjXLd
hxcLv3YYPrGUu2v60tYT+2heSMtU2rW3e31SzQ==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
gI5rNyG5c3drysVsOVroSrr4ZtWR1lsLBTZK0baFAq41KkpdWktaXW1nX/+2PBYQd2WuwEzYgR5A
3R9IbnThHfZMUVpTqmm3QCjUOIk8nTQkx6iS7xUYHB6IvuSSVzwXQYY/LqkXQLggQMmEXSMTtRg7
Ork1pXzde9DisVtwZ4c=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
bnYreZri/8cxBtUYrMOxeBRiusm7ZutmnARaEPgJr+swerZuyUOJZp6ItrV3CgROOAJPmjtZ5xM6
8p22vOpGw0kyktH6b/I7eW+xyPhz1bhIfjHoQkmjWC3hZnK7QT175CxgyM0a8/ioZcEqkVaKhUbE
nSPalwFiTDeR+NMIeZCpkb1Dre5ForqsAJpX8FI3X50m3/VkpVarXzYDZwRV0rJ2y1K/44VnyXVj
mQsPxaPSEaNs3ANT/XC25M5+aakN0smvIpd4uv/LSz31BvQiZAUA4Sadb8OP3AXdb7KKmDrq49oL
v0kfRFYGECoXJBlDZldG95v21lyt8fj5NUetxg==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
isiZwfumseLxHBLiIld+QGY4tmJ5ngxpWNiK8ApOc/PKzcdGQqiUXP+VgYMyH5NFXIvrL8Slv/Al
srKlPMKwyAl8QV612cY7tc3fHQsbKD5ebSpDKOBmvNA9WNpA5PTQRl5hXDd3GpUhPpxPVx+dfsVv
YxjZACjWp6636QxL1ZtwQk7em+pvgGpS0osL2Cxkq/x/Nu9nXN4mo9pBi0mWfdIbZsWy6Mdjzgx3
jW9wsPoJ1Ne/n2S2xFex9EgaCrfvH3v7tuVNaKtsd87nvF9atFT6vcr8VVLPnWW0lVCmY7U49TtM
KcqhgUB2Skt1rkmdS0rn2etqleC8vdiEnTMhsw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4768)
`protect data_block
54C0tOwBZ3FVAkNcRAZEHJaG016DWwH4zq1NOqcRsdcdrxhNyF5qc4pDTb1JiBkseoxDjSJ/p/Ca
K2bXO35ShW8tJOy+hThZlkdYqCZGJY0ihZdkhdnFKL5r8ygjDC0n4HqBBhq+H26EyA2s3zGqaw+N
TBoXVlfe3u1AWcgUnRkKJ79BF7Aqkcj57i9A2ROxdWwdPHiMnfAmUQPzYkIcjRMdcSzUhV5OR4lZ
riH9ki0vs85JZ/4tcq/U3EMf8HHz0PrXg+R7rUS8B6Gdp+YLoxvTxmIM0YWMYPNDJH8L05L1gSnQ
wODfrrjnmCP56d2DGS+qXKgSY+kuk6s/KfOkNj7jXdIHgLlL7JGe6ZFGY9qYPYypb2/zd0ZIXM3s
Nd3wp1Jgk7sda9MWnxdRN5iYZdxJKDaP+Hx3eJuGOAPem03mTbS+EZ8LWzP5mDVRjKryt+eaIx7L
nh5dvb4pTOjNGP9FPlYK+JcQzSj9qHZQwCbITr1TEc88tGsDTXOecTOU50fvApKBctcE4Cyt5gl9
q8zZc94TA8B5GegOqt+ughyN/sY7NXs0C5t3U835h6pxfdmgDqP75sQHBLGX56edbzJqrCJ3ncFg
s0wFhBLje3gVuW+ZZo3RuAtWDBS5jWsDD6V1KM46pZBvvhQ+WgdcOtudSSS1t12tnOFAVTHEZjgy
hHahUauo9FxY7Zc56gzQN1csPUmSqxsZNAn0lNAyVFBvq0whOR6egNwm0/WVWKKlpv1UQsqs0uuT
KFRCIiTJREDOqTP//6S4DgTUWd5ZtdN7mCTZ24HhYe5jreLOyXSljANZSoMrQINNlwdwMbpkSKnC
yrA9ZLOSGMBQTJLiYviru+S6M5dn9CdNGNyyytRg8jsGbOfjve+oIym7oI8EIN/fp4PKZVd78rTG
QBQbqKEJzDAOezG+ulqwyZcA3JgiXcn7d2iHNAQqldUEZXpVMqv6g8uLUUufD+E4JUfVztqFfVS8
fO1m8TYPfPYlObpS6QvUfjBmdVEIFTamruOjrUE33IN59qI2nBWsW0rRb7E1BTOOTJQN4dm8WwR5
Gs6dKJnF4VWa4kZqhtN+ypINUstdz6bVHGF6xBSVvBwD9u1pMtQJAE7a4zHFFBz07lRCbwUGTAZw
2l2OURGvMMr8+YqnpQQxIQxv/NFw+AA9koOd8PEgDBpYEu5r/bdsFpLQwlOa7I1eL9ffk+9XMvTS
cRIli9HuhqWWj75Wpp1SeDUI8T/J0OhYAGbWJQsDIlLy4FPN9Lw7lowtI0FWoOUC2B4bmXqIfEXg
vHgaUuxpdWHxAkfrrohxX4s7eHMv4k7/cqOgD4cJQaQVlh+wXGUyMXsduheC3NUTLPuxIaffQLlE
C9kO5RjOyn7g6kRyYdqwhRwNAnDLoGV9q9fWB83rxZ6KrmuxEoveWeBXrPVFQoeZhennyuAys4E1
IJ6govnQf/2FxVH8TyxoKzrUDCWZTSNtEJWvSDj6pGEWpacdq1KFT+ubDZ/W5v6e6qt3hSD2EOAq
Sx92mATGEbSqGJpw21QzONv3ZgQ9heIM0X/U6kvKiMhXQrdIjlWxOlKeDWs6en3LYxvp7nHtRvVT
pN+b5P8YDR3p7/Lifsr1Bp/rAdGaDn9M31Y8hOvnUv/qd7agD3PMA7mLG+VsnbG1z2OVJWiszaZB
Otl+E1JBUxAsIEHU2WxOV7pKzLJzeKiIJancS1fZdvcg7krkTNx+yE2h/JIq2kGCeydpT877VGhx
chrqOGXUTSR+bz+wIDZLxOs6vhxVDpRNjEP6YMTtA44VZlQ2C1KjsuPAm2INfhMJqFzE/m2r2i8e
puR6ypKxUXIDHZiYWX3g2rrnq/O4pYTzAI3xpKGsv3jzXDvtuB+VGPIxr73ih5BzfdmuCKHiGivD
3gldnWTMso9YBznLKLoyfQdq1s6+beVrg3Bvi9k59Ftzk+ZsTv/dgifGyg1X00SYjRt1eBJD1zud
3Buryzp2Hy+ybBm4P4qzEYYh6OmCy6Olta+7pB+LoIBMFbOg/ymBNJwTshXdJ+AU7m/Lphgu49GM
F3LzTvBfyZuUwhpvkcBVEisN8qe6JJMbRGs00RihS3kFlaGt8vBVhbsONdSjsUmY1MjWRMMj2/6r
fIFptvnD2QIiKg6PWnILeTROZo0kSD1+LZ2+qW7yM0eg0BDWnmZfuuCj9cN7fseomP/fINs7+gQo
A/bZgJBTA5AhjDfM9kYjEvW0XUL34oLuN5Whf2Xg6eHE3wQtYrT9tBcT7IAneIObE9ZG5Muvz75D
n2a8Ppxv/ZE7Abr6infSkXb0A+D/FfCwdHJeQnS+OlzWiJsehtFJF5FdxOG4wR7t66XYBtiQp/HX
on4yUYL8FffOeA5yyIr6NDe8qQZEtgrmY/M/45eiuC35i7+2gHgQWj3v+uktjVaxtLC8Ao2yh8Qb
yXo0KV2wW9/LYILFgTBDsV/a1ypRPmDP/TW6PRrwCSHjZl9ml9wLSNSlFWeMdD7VGm2fjxeHIDK2
n9S5OaTy51yLCWwYTZBkyAifjkByPe9T7k2cNaQ48vCm4M9+zAvYRmSyZMkmGpzCxbfR03u1CCoy
0X1GKApWC/QMEFk2RZPSwiZgzxHMuMl3T/p78WR6ap3w2+X+xwEhulESiz3X5gAzZw4tduz1Ujny
O4WqwTZic0W/BWi4XmWiLdjUDPdV2rWX+MtkA9F8cZXRf7lqMGYb2QLQ6MuW0fzJlyhiyL986CMR
j61zVaD6KKJGgjB4SrzG/d15SeyD36ntUbutyVS8fs1tdw0dVuRMqe7MYI7WwR1JRrsTmZaThLx5
DHp+2aIRttF+xvZsCjSwNJHQdB32e/lA/O2L7u0k4WJOO68XH8FaTUI8beDfNUNVtvjQCD1Ufelk
wXBkguCyOtla10reRuX4otjA+gevax4wWC1+3GqkFSb6Daiw4wrTX7AftDeUcQ1i/y+cppW7nWll
mj7yYut4fCzARh+n/C87SIhNhKLCYLhzLkBHFUFIWUk+EM8AirFZfH+aYhsvTOnBP7h/z6ElfLOk
U6iRWfg604smQ9E6jwoSDWMXFR3kT26eZnGuh252E12DOHmJF+RoTkyO6Et8hhSGCKbB8NImR228
ukYwHPG7AJmLj/vEK+ewWQXjKMksdYmQIucma2MH0eDY46bmhAqR+cKSqV3GUsz86iVEIlVNP44j
uXLcYPH6P3YOT2XY7wlyD5HlwqqLq5BPaovvcz77fmZI9U5d9iI2oWAIstlKB6CFFgqWqYML6rFE
IFw7z1h8mAwE83ntqkb6MWPZCKmUoFAGfvFHQPFhKEntwEAGnvt1N1i0arOkdOkaWWAUafSq56KW
/iqgaQuGNQnweVFh8EtngA638BE5i50Yd2jGNa3LVkUY1yS+W9B7C1PwMg8in/nRP1ItQbfBuN3O
FrGW3EgLixJg9pekzF/UsrTrQJtT9ZmZGPA+s8It/Ira8Weug5jgbjTEOINcLnrVSxX2A1yq2mo/
khlBs34WFc+HslqtepmpGZgqmmTtiirUtpKRJag4V49Iq/raguDSgFjJgxZ+MzTGXifHLrmied0S
qFQ4fUzwrcX9nOjjJuAW45dHY/dY9Ya9GeHv6VCZYkpwxEmjRz8qBE6n/0Rd8bXtWmZA2ny4qSJl
ygqQI+Qhd87AErOKyOAInf3ZRhoiTN5wbKlGD3o8FSRCebKpAa0VNMxlcmhTF/CiH8TqDUXYFXkN
FjEBOPg0TLgD1eXKYtkOpV/IHwdMBmy+bRjKzIFjqO9pzxA9YULB+yx0++LC796qVdNN/6XDCeGd
Fj7gpPX2pvoylMoQcJtYgpkf+fgAaCSVMTa51Vwd/k0WAazinmHFuYGiZ4eMZRmF+N89DbyfnRA9
Pq6x6Nq+b9x7x8UC1BGPW0BPVfuOrz0tqi3Pbpn6GRvCzGHHkchy4GWgxFASoIYSxbniFY5BwWRD
dSmkC3jZAsd22mkkdaNy/eJklv5qVZ9udR3rOV2L1LCMF2B/ccGyiVTLieg2z/UilRN9fSXpdXJf
3FdRCxjkCbIDL7Xg6x7U96f5lNBVsZYJgV5DuiZ1c4Xw4THDa9F5gShaXqDl+ZHF2UEGrf5VAtLK
VexebLITPj+avAZ4J0XNYeNBSoQPJ5QqYNXdMm/LDfgkPCByAh7KSf6d5LQiDzT0xWWL1JtzaXAG
6AjNbGORH3wfJqNGxx2wButaLiOWUZkzMpKdqwbWeX8iV0leD9Gb1z87eO4x5pyQxLJarYMhpZq1
uTx1PguPTvEw6IcCWWRo3Jth/Qql2PJn8Lh0v8vgoJzwTaIcybLNBV87zVdJsPRCLfj0vMXF+3gU
36n6ZXD09fBamqdcJpSSdPcsmRkwYBNiSMlvh3btjBGtTi5v42MmZZxebr10FrW218KNtsnxltpM
VUAu5m/ygEqp+kQT2aFLpAMpErkEsLPnqjoJ97uF2+GU2wpxrvMbg1XVvm+xd0vtx1PQaTGI08ke
qHl/PFiJN5L1aQObta8C73S4MBSQYN8Zmqxfn6r07KLgC5NJuITJmSMcX1jK6WHnXtUvJ+reDvyv
wRYncW9RF8QNeoe1GKbztYavTOhm5zN01XkA/6rX3SvtICb4f9YKKlMvjFbtR5UlCEKNLYS7gh9u
AN4IKRTYCpKixmr6e960j89H4fRSqmPtCgCZe+U9gejR3V8BBrKhAKZwdfLvxaGDAALLsCGL5AWA
dGtxAro/DQ3KFGRK1JVbosOlmTLIhKYaGpH6jOgiv4iqbdqJovkHvOlKOObz/SpsYD/E6H1vW/Kh
3uKrpOkT0ig2SYZXnJP4Aa1x8IJgIEBCji2sGFfTc68OfZgcMWOvjgMCWVUlFpaXZRCHrRmJEywX
fi0bzdfI39eawGIpNZkqd8aIysCQCG3l8UilyAFz7XDM/Nx+DdR/Moq0Dqxmu02ZaNzwuxPWhJdI
MAUDHQOGvvF3j0FHoRxSM2UUnxhdZ8v50XG9ZWO+SKUXLcwdHby8onC0bC7tAHrZVeIeOJVSgHtP
gLu2RYekvbm0SfGDWLPO+YZRNgIWzBaay8xEpM6PwXeIRCZvi4StgNBZnfjfkwya0OaaS7tdIrP+
sLgbZ7wdu1dfWsRlnEDFrzamPb50LNIxOX1yWSwKHZXmMNVhKTOaUgo914VbWI6diuXnCVRsd/Br
ThMV0hSOrxplK+/S3YJmSDcGot0hOvQhZ4aW2ZA79PbWbB/sYNfsBe+UpFVPED+mLSRGKIW9kEeN
1Hl2udxh9YcL3h96AQa8KVaw6HR/tgMEDmHryBceZxvKLvNj9cxSzGUdBtryzCXLu6tsYx67dauT
QzN4JxKeuZYgpLS3ewvAPoE16irmaLI9mVmWqBtp3vMiwBg/dDbjHt/iiLZUrxWYMnXkLY/HuYEI
3ylIncQyoRLzqy3CP3iqFWzwdnoMa7eLZhALttvh+nmamswhZg3a0vu1Y5dGn8Gy/ak/FtZo7Saq
SFa4ORq3FkFKEeSXfo1V1V+08Q/5WnDUnrC7zro5bv2s2L1+60fbVTJVFLcHYY1F1hKn71PWj8yY
suKnxflczKTdbp3KqYWqhMOReR2Bwv10SWRI0Jh62uIeSE1CHaneJYQx7nFTysQI3ZyrQVZOeIeH
BJH3eknwZ5br5NUDxHXq+RIbI/7K6J1vaqZz3R/oZJ1/Q47OCrmIbhgTR2kiDqFBYoIEXb89A8HM
/q7/SyUvc112OxilsIyWCr3+JyczmMeXqiyMTSFdrevBLUul10aaZnC/H22kOX2Q83FYb+ycSEby
bh3dcxIDpgikwRN+Qb7Q45YMHSsIs8r33lNMm7c4sulWjvsUKS9cex6HQxgt31U6plwusvBSEAfA
DneKUWmkqkynCR2JpSii/sQSJlxCYFns7NeXwYICXJtQZ17vvLFMYbStccqHTldxV8d627XDamPp
fQXLL5Mtug1bFS3xIGk4yZ4fsxLHnv3cQxldDEUAp0zJMU7Q7YEd0BZS6zp+v0yn1QIyxTJAvUD/
qZUi8eIgISDwusVm7jMesq5xyX65ifyGC1mKJdcTl3pGh7oZ+ZcVOBh8TDBWw1ggrCG2eYCH3n7V
E07u7//EKO5LpYe94xkSptIQgX2ciiLwa6bTNqu0eLngSWZE5gAa46aXE9nMgQpPUEORI/Ar5xBj
KBZ7buN7ZnP6SPJKuLQg1XD8rRgbSMHOgdzVbgm2mECjUDMy+sSrgJUS72OD6IXhe8igtRZm8Fo8
DiG5o8K6raWNjmPIjIYM7L2qqv86PTEee/WgQjOUyldribTsyI9qYec99OUouqtyYKjpu+0iLWon
tFKqVszjNk+BjVBLlg5lmgZE2kPY7QauAYtYV9W3DYr1b0WmJg==
`protect end_protected
