`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 3152 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/9huKRhRMtvnNqb3Z+UU7TahEoHV+T8U3P3ufru7l1O
3DlgtZzb9QxCbOjthp9+wDkjygH0eUfDrEl1ovhZG610Kje4HgTZzfo2Yk8ZYLRo
Rs1Lv0tKTgaXUjVWrUx8LjbxDDiDQDh8ev9A+gbc1V9AUz5XnsXm+FMlhopSDDPs
aEHJBh2AIMxNK4ilMPUBxB25sJVLlGojZvbNARlkDdDlnRZAvwDq+1NjqofgRE4Q
kvTosk7ZBpfdK7D0RL2zIWkOV5XuhcW0GU1nBr1n97iizy9AfEgO/ydDmFTMcMXA
zqGJLBmziZgZQXwsTrG9/kiDwCtQ+J6r5odxszPd/LgztU6aXOOW6PpGWBBHUAQO
jxm+G5OAHhX5yeh6LpCWqHA/gj3n5kxr0sNma3ea3ZT2NN3uAm9lt0VQQ3fJzkfR
njbdnUU/ZD7y4/IjgMmKPOT2PEaZcmDYwaliSGwgJoVvgTKgE+wuRayxIfO+qOhK
JwPb0nZyPeohQDOkAbgGL9P5IO67/YpwaFbJ1CeTtQzfBnnK5pGuqA+A0PVcc6s0
t4gteOVcFEC7YL90zOSG2VeM+9Nujikc8z1OKuvEthcqSYAMG2XlpS8voPYHmLiv
YckTuO9RMJDgrj6e8J/ObOmx3NFhviiZQsKp+K744YxK/WHwQ3GQk1QOMUsfv82G
VRO8xi8m79HIBNu35uo74cj0R7Zx7M77dc8CUkXfXGQWuSj69NGhJPjGlbRuIm1b
kHDXoUQr+J3LjhR8mztOMQrL726LHq2mMSzDUYyGkelihafb/32OQ0kdMDPwvblJ
p0z+f4u3LC14YKuDe/u+qWq9SggbWDj1ZLs3yfAUQhxAJE0U8r3woabMVVLFnVd3
MN3SLQ69nuqAOFS/3qPjenxVyymUrxo9bUuwZ08B0BnHSW4okgoVym2vSJhowKhF
ygF40yFs69wEWpSKcE2pZyQ6GDyv+3xERUBDAMX8qtTEYMzgHsKPH8uTS9LTjaW6
twDQ1kkO+8YeVrPTjHUDLZNU5NdaJvQw09ayfPc4Uho884ZyV4ri2RT+FUqVjEZw
5BNvRQXkrVNeEDM+paHStEwiNi++2rY9aLP6fF5XPAsalFT3hnpkhOn8wE71nasA
rrZCkhzpnS3DlQt3n2/Ry/ZX/1PTftDNriWwHEGCHAlkCsCkn6MiHSu1IJQeihwg
u0NewWZBnz4xaYhoquC1P6tfElwsf8aErYokUGXSyX2wbxoAkXi/DC8p52zztdHm
hr0vL9zHtHZg/uAXmp+xqi4GkQuC2T/H283aBYK2DFSdZQMnO5CttASo842uvFfY
XqWPsyzWTlNM0FuvlXJTzuvCCxoDmcN/9pGioy2ZLSL26y09+uMBwHZdNSOLX0eA
M5SScFYZZtpBy8jZ2P5LUZMGzjF/ZWlv2hXADULDH1YozYBZ0I40jOxbMQU3gLoZ
1Tieh4tahfXP2NWsfQ7Vq2k25v6jsvAYzc3UGmV6Mlqvw0AxQK/LzlzTVtA80axX
r/qikdu/eTx0vvmY5XetANBT59xvrsR6hwdZSQr6nVLRTsnx4mMz1pvepwhVt27w
UpSXFJaaI/SU+1dmlqel9inyQ99Mk+XiX22hNw07/v9q9NcepcnHLNdqoy8n+CF9
h/vqtn2N0h33x7dzntz2Yhxxi+kwNCFLQQQ5dkOI95gI8HJhblP5f9J0AjAq029j
+7KKL0UJ55jcHhZ9Z7PNYN/2p92BNOLT7fIYsSY3dDaUdN+YTh+7VGl2Kor1iakj
FNayYLiMvySzd96fRth+OCiiwoMbj2cXg8JkpEiSGNP9S4pi7PGEGjOwPgQuuJmG
h4ats3+0j3tbBeLAmW9FEqiTyMizOgG3FB1GWzgsM11Q1TxZ/vRjA5ck7zhmbpwn
jzps/eFc0CO7Gevi97NeSzAWCOlyO0nCHgVV8pcZ5z/97rMIyIJ9yOPmH4UcKHjg
x638TCDCQMx9KscZaHcw07FlR61UKNxpeByDHYhZK5TSE7Vmx1GnAb7w+d4XM5by
O8cuuFrcGYVam8X6UG4TtbecUHNodNyfwVndUnuZAQCQKJDSUML+qegezJQ70ZEH
HR0wmaYIh9eGdgDR8+cmkRIUVXHPsNcOtpf91vbDBYra3Kw812CL4hk7BbObPEB9
V6wbNqtau5g4mpiwQrnWHzHv5TUaiRlDFdmcj9L5PkVu0sYZk7vYC8k5/jPAKqx+
zLoiudygDi9KlSuxxf25jBu0Bl9HwHZz6a7WhhIYet47sVAuLhp8Z/Vnj6wjR9zr
OhJiy4PbYXGmryVL8mva8HfzpdabfQJDs1HvEN+XKHEjkAZOweacL2eBkNagmiM+
AlEz2HMmZeqSsRVkP6V08mMWdVrmKKrJVxPv1g2jWroY7qLxeX8Geb8GhNk02dAn
qY8yJYDPHpuixJAWKiobowA7wb9JOcQwbMlB/GsE2eKpKNbWHXpuNiPUahUkTfEv
xjwMugkaHlm3N6uoNLwfd+iVBtkoTt8yE9qIAb1CO05mRn5NytHxDiA/sQ0xbSCa
Vons5hxysRTnXosR4p0pBJuRb58H+Yor+Plx/CGjtdElOvAppD+tlFMfoDHKwvZS
UbwOAIOQRcoT6FwMvH00bnBmbp7/1RT1cLOl32ipy3ZLoUzWTRF1gl4HPTJiuZOf
jlZ7/dF7eR6bKVJJ4YSExcE96eoaa0qW2JU8y62gGYJQbRZD+Gvs/0Qrdx2bdCcy
COe+UhI90/SAU/GdL/l52RG3bcW9e9MdOoskzDXjOkzgx8C9oEUiuxCcNv2mkm/J
tk7U/fRDhR5jQQh1I5DTRB4QzXCGLB5cgcYSArrg3sHDDeCc1i8LUBJoFt7M2gff
wEcIijOit3PGzPi1L4/pG/f8QMXIsxrsnpVJU1GT8aLDf5QdLXRj32GamWRhyhdr
hZZXJDUUAZ44iQzfEOUQGf8gsxDbTJiiDgX62+q0shtYfA6KCh+4yN+/cXoIi1RD
CVRiopS2iAtbBELvit5wAo8vsG9rDf0ViI08azKp1j4apo1dXk8mRmOtYD2F5Xze
ruFt1ag14rbvmXaQoVUgyA0W/rV2Pgb37xaQ0ay6rKVsq4RzJaSGsb4uXmiozySY
hQYMWPTz5ZDJzQYmRf531SFnI3qXUK2UR8dttcagzwk3xsPQ7lrlMOQyz+MF6MML
1V+hulOEPazBQw0lQvRu9BKlNyfY1wOF+B1iEk3rMvGQST3CIHqYhF682mMN2OkS
PimsYYodkgPNOCxcAKF2SbVpMLzPDwu8BY6RyH353W+azsYQkebfjTg4P9A0VOCN
ch6NISWJE5Oo3W5DpAskPnBod+thLMT2Fvf88wVSLwcSW0TkN4jRsWWkTl4ApFus
dvw3GoHTzyauqVtF9wNmtHgiAE03R1GMFuSzq9Z9gzRpGYgs9B3+Dege+OFN9Ot6
unsxw6QEqqzzqvKte5cOmlXs4KSY5kHMNoQYJyipR4LqrneuvceU/8EWquUXNcty
zGrt8JuxnIH21exy7Kjy8mGTBmpHNsCiqC7u3LZgt2oEk/nPyf3U4AdhK6mI2reX
hTzbkKd3Y+UuBJmhI+Wq7JaQltu5OEQpAyrzoX97y0qSWUdKhvM051WOPneQ8CW4
OiPlFuh7uTAXGzXQSI6Xs/B29hHbp/XmM1I98oIvBRqlXAFDrXmvJfYxOqFdEpDL
x2N+dw8T1/qbH7UAGMnHMNCxb3xqjrcoAe5LzwbO1CQSIEdRKhO0vqRvWT6OcYiM
givBxcQ5k41rS8Y/aRHciGVlhag0l0zT7VJZDFyOq0grKi9foZGoAJBImBZWWG+G
68Q2SCAV4EfPLCXYRO3I9oYLs2Vogr17FaMIf1Y5HP/yqc/n0dSSVmKUKRd6q7fG
+P4g/eITgBRKnLOQmwqdAESHaemjXscuKhn6mqyQrokbWNrEG5IKK4G+uawebcde
ZOy9xIzPTNwZ6KNrQj+HPC3yk8DoCzphET2GT6S4sWU8QXtp+vGu8/KSB8kPKFsb
l/FRNyGu4/SLy7sDH5YR8OLQnZwSaNw43ys0ezn0/6KgzmrfvRWIIXCFYWpzlItZ
yRQdtdHIaoXCePB/iODTw7zeUUHjhSuir0tG907FieJ+MBM5/Cr/zjcUROWC6cRZ
5R0tW640EpYgxw4Z/5okLPZfnam3hwnV2lm2q5wj0EQ=
`protect end_protected