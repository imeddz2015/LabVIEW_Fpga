`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 2544 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/9huKRhRMtvnNqb3Z+UU7TahEoHV+T8U3P3ufru7l1O
3DlgtZzb9QxCbOjthp9+wDkjygH0eUfDrEl1ovhZG601IZoIoFqmTwGFM0Ymq9rE
Y6DZ0TjgV9RKqugNVFlRXPhJZqCgNVaJjhoEyf9FncGfAJsgCijXLVIIyGIXUWIk
Fvu7JixabkHq44DwOtbcXj4IKdWF4s9V28rQVzofBDPX5yrSi+wofMoKyX9k9D1p
tCX9jBKL9T9O4GxUalvq004jo7XTOsK7WAIPFEDlndmmgHStb3NTb95RMAjPiO7N
2cdQ7UcHP/dACFOoW/mfjW0905k2dvNnw0PjDXhLf0UZ1ko1VOD1Rh+1SsOyHhf0
iVUTF9TA+mNBXpQIsiHZzq+JoOtfsOb+FKflXkp7N+whp97AXY20B4ko71BPDYtw
WA76ibhJmZrOXkjd34rKKq/MSaHHpwJIiFDCw/uYTB4hN5AuHiEGpiMnKkiQNMD4
LMLn3Rn+wNP6Uc5LzyeyX61YXgOvOw2waKsWFkOqWwFnZbunJAjxWHyc0WY56Ny1
cY2HsOlWjUAFj9mhdfnfNi5nh0C5w2zEnCLU/qsnNSgH70UE/OH5Yyxp5PMYmp+/
OojR079rDlhR5UMsgxfeSg2arn+e0qoVD7QI9r3ZYS5ayH5w1Km3N70Gl4xVeQec
q1F4ir9euvjYvXtk9DIxKC0wEAeXGPQeUTb6L8g7IGMo6BYvA18+W3Bs4dAtqoGK
yFlVfesKbs0zw/Jm1Nr9Nt9ZnIK4a728iAnUh7XR0WeYs9WflNSUBp5Zq7NJOwXq
TZg/o2ucY9TUQHTPfPUosaOmp79XjKYGnTBYnJQVyb9ENKOLmjxUcuuK7MyHg95x
f0xSzGndCq/iQwbcwZWbx9N8LgByUFsWZwVQZHpDyHFyCziaHsKcpPcWZ2P8K3S1
Bw1TBmpzz+oa69Ect+Fw1WJ60bvpO3NbVWn9QzplzzUI4rtmIfyE6GbfOvzGmTrE
up2VwrDGV5lCSIFxj2AjLxF8HrzGKTeXBdeJfdAPQE0Q4kZ9skXp6XN8Q4pIFr6Z
sh8H3p8YUJ0KxFeWRFVfBCvTizyZZN2JZKLf3LX98luLMuN1VP0BWqZiyCf2u61E
DwG4TvCpkzhAan1Yt8mjCeaEuqHguBHbvO5bwCK/DvUzR01QnyRM2+Y04KZyAuBP
tDtORuB1BBa1ZFCxJICWR2EY4/ZI0E2/LIoOVYl6DAbIGV5LQZy4h6W8vK2Kf1kL
FuK8Bbbz2qrSPBjhbdEh/uhdvdzWFd80lu1mQSo28HuyG/pt6COg3tBUbey8RZTq
dRP8phvKghc9JkdUwA/jbARmH4q10U8UwHjaAf39kxdKTScqI829olHMHk1LPVxh
M+LdnK0m1vuUzBca8bsQjMs7JvXrvJZyDBRPd4Bns1KYRApARtEUlhQm4tIiPCbF
Cg6ewwt85WIxHvuRotOSZ7CzhvcTgRPuAdwA/Q65lLLTdpKP713PTCqaiHtq/WKI
B6dP+TZwLdx61CMoidCw2sihRiNxQuFeTvnikldENkHSAwyhZsYKCmksnG/AbTdB
lOgInJ48Ho5VKt5r5zXSRrbvAZNArIVpBBk/SOSBUfkRktzzXB6nOYqAXUPzTK8i
QwWGH8T6Y5Zdfyj9JX+cyxpOCZhDEZ6Edh/HbuvtnhBFglxS6hvwP/Kpxl5G9Dh7
Z2Ja4DVdOEligRGjNA6vIIhggyiQtDqFncm6x9I6WulsLTmAKVYQP3JBE3GngVaG
4BQd03P0nfaD0KubMaCLEfjuhT58F5egXkTKP+SjGJGNFcD5KUtJO89zV3Hu82jn
yorSYTO1XMURy47rgyvdpQaBuYm6/xrF6YFrWX+rPaqj54eHMhRp/fohbdy7jq1k
w+EU9/ON04uyEVjUD1zDFccVXuVozVHWO3oCbL1AWQQSWOs1edkfzJNeUBKDLshJ
cPX93wl2p6xf1uhoa7KcmSUDDuYyGPJdPCMQLxu3V1wHJCv0jdiMJ01Kg2BKrB+o
aMmLwoGWBXXF1zL88IfXxu3VOQ63KJfPFJ9rzdzcswJUeaPzZ4J7yAowBwssTptR
IpO2MieFWYGRhorZ6gHIMY5LLclwLq2Ad/3p85Frz8zh5g0NVvO9+oCMgOKU12kC
cGN7g+5q52JMHrATKSAxTsf+ivEYuytBsRsknyXOEj+p6dR7+qKuO0d5PwCpTmWk
+4QNtxQA4UuT81bAj6nUTy5S9ei5hyO/gFof8XaCkP3l7xIhc4wgLLQv1W5Qnmzv
ReGA8SV2nOHUzwwtL04W2Y3cjqMeArWSAw7tKuQ3qhFsgtm00htM7XL78arCC77B
pSe2DvfokROsOLKcd68xzQPhTwhAewt+iFUsluKs/Fm6NZ9ieKkgEkF1FdyO+YKO
9JJSydRmk1Miv1CGV3q43iYqPTHYtje17HyGH2fdYO0ENiOLiAlg13xtVXMwN66L
lood1l6qU8dzdkptcuUeDIheVhmgsFAYYriP0D+6jlNHGiotMH3Xj8ehYPKnmLxD
Ntn5cd3Ey7sfNDc9KwtLyYobeXx096i9j/+V8SIOp+GpUlRH+eKLdKSBGkEitj8W
Jjsq66pk94i/AIqQyF5lMyk7ZxrtC3GhABsQvpy/HjUFHGJ8VhSY8UoQXIhDaoC0
tei0rq0gLZxDAY8NB/ofmfK/Wb76cWKXNKzqcmyDfl/FXc2m0zZPe7CcHZPtQQMF
6dimiR8A8a++W1Pv1U5MOT9CbSk4MzVR543a2q8Ond30vUu/dx+6vp913ZAFrayA
010sg86N4umr1/KaTnsfMwOJ954SDQzCChgducxpS/hOCtpBZq/Wpb5XgQcj7QBl
eb/Oj35OC40BKuKJb1KEOyxLKNBij1liTKJV7+FiUo5c9gEtCOVb39mnzKadQ3wu
8QS6zUdD27B0A7WEvgbrTOEAHpuobcfOupiNnc3zYHVQf9XK0PjXD+lP+TLTmm9U
vSWuBYfZdPmDPfmgiroK6RV13SOQh12NegEjfFDKdavZqieXtr4PHnBq6S1QKqOM
Jkl7YcpevaoaIOJnbtYAlehuqSKH3Ogy3e8XE+fm0ooDbMehyVIAi394z+bKpfIY
UDWDx2YVA9hUynzICcXc7HC8U8eidyNC7iAdAgqOPpHPvvKsgHRwY43FLM3KoYlm
w9mIe4mfXp13Z9XBy1hv2Q0o0X8/Q0YK3tzaEr36wZmQwnPNghQxWyOg8bEZwV6I
LRjldvkXGaa1Mdkwigbjwj5YcD/6Vp0sHN344CtNm0+Fv+7HwmegfNE34fDqieLQ
nFHrH69RwpGucQuH/EMdklGE2ogmjnQ8XTF94Lu5gTdw0LAFiJnY5W1YhKi4tYEa
`protect end_protected