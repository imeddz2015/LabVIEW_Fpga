`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 3808 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/9huKRhRMtvnNqb3Z+UU7TahEoHV+T8U3P3ufru7l1O
3DlgtZzb9QxCbOjthp9+wDkjygH0eUfDrEl1ovhZG625RRVF4+6Kk2oUkF/bqPbg
dvwvLGeBWS1PgFMOvguG+4ZAYH8WOgFf/ZTf6C7grtfrgkYpPsaTjiU3Z1bdTwIa
jYDS7pqeSXAHW5TRpZuKYxeB6RuqnUxDGPdhuR6bInf9wjj+tntYQVp5xcgUOnI2
D+InfR5jGL/XYDigvSpF3Wl+pDChgcutkVTNqJPIWdsOQ3JLG0Z/K4WNV2yaLiAO
eIrc72R10Cho4ga6CAVaa+oCNuX4D1mGiRzD0ZgNiwZVuMzLRfGZfW7l5Qnx6X8j
gwPoMG9aHlVXaUTwhdUbJNPLQ/Azvg5NGk0v+E6Gf+bvVOjsCAyUc9fN0AW2PNEa
PuFme4v+KubX0vya8JhrOhA65Kmo4X7jHlT/jPz5IksqMecwtl4757gv6Q5V52ks
qJ5xtYV3AQ2DTDj/U94I2hEjKlPpGTo9QTOKF+2Eom4fso+GNcr45um/9dguD8e3
itwx2U8c9I98DyxUdKR8JnfDgEAVdzZ1ZtAPft0Ex6VjPKgSxs8SC0+4LmmxQhf7
mz4PfBQhK5g1xeN2g+G/3u0MlK8uVSeBI79m50m5VpWTaAz4kP7Y2LPQEV602KjK
W5clKwXwTyauZVH86e9Y2tBdEClq2eA6eHjN6jYVNIc0JZyLi+toistUXbh3CW7T
puwUvOpEMbZ4v932iPCw5A0VENv7qkqvDAW2e/muECs8kCcK1qROz4mLeTeP1NaR
9EvTE3ybLZabHcUmp7V8q7EqQyK3CEEOvGr303E6nvg8QhCxDnsCFWPAO8okvLUy
x0Iu7F0ezGNWjzh/TzhwM1WkE5D6d90iZGRkup2NHi0mDOtGKYz49UfFJoUFixMC
a/8+S8ZKyUmcwqeyxM8+8Vjf7+kfqGwrDwrljYEEzugRS2OulW7TWv3DafDflZY1
HNzlFLN1x/AUaSFCFf82JTyR9RogZAOQIqj5bfFrlqaYgMwb7QEbenU6FTH6vmff
RFXFt5SNLUv3MD6/yaktgxnRfTqpALI70r2o4xdY4AGh71ENQIdm+ZB/+iYV62vo
0W6jK2Maf5VSD8xJieLLRa4p9AruMQNzMt1gLwLcR4ZdAy4tzfOMjxUBvaKRkWWy
qXH6i1XNNG9wVkM4DkwnniHog44RlvxkAiBomaObUZsM4CwAmiImrtdES7Ca4NHQ
oP0aNUKqq1AGgBL7UzrJHBVml0oMJpX9Wz0djgcuYYJOR/2uR2JPOE01uXLgNiCT
V3lxmfdzY0vvk5WiWVudaY9kHUmayhmbM5t0e55tgNVPx4BSC1PcfXbPjHN8RXM0
DxSnD08b7S5+VATY8v+3Fl/KcRMhiN5Et5mQXCt2pjAF710XFP2j6gJxb4T6z8RT
Wjts30svNvcGJ4roNwATJh0HozNcKcDe5objA29AVlvJi/5PvjosiIrB4NnkUY3f
m3yRbD4m/XrMS6XeNo6W+VHStipLmod1kxBvxj+dXkG+I9Hx3p6rmmkbtDCp6xEZ
xAwEbbUTv8cx0LUCLWw/awJJE2/Ycpq5kwtJkY40F5VGab0SdIh8PxLkMORiqgat
E16baebFK6BvItAVjKTTk1isTUMdEQcQlU/bbcqbQ/BMo4kJpmAd7X5QkSR7gaEh
C3SOBrA4Fl/r+eDYb+QCqHXtril6sO1MmF5A19+0vTDoeI1ChTVv6d6QrXV0IRlf
bWqO6XQVRF7ccgsaffWiyobZToAo2K5jBgMW0kIAf8g/h7Ei9DBb3LLZvm0nXkQC
nUNbm9IKQBAhDHu3JH9IhbQm/TPghL16qWrdJbxLsSdbMzlj1Rvu2mZ+Fs9ixWdM
ATXCm57YrlAwqBj9QlWDjQ6UJSMJSEj2Z7ymbTnKyFFFLUNwZxMUf8TBpTc87Qnr
Cf+8DZiL06yhLANoWszJVgnoH/Ea4+KejLLuO1Hu1JkGlLSYwV1ePsiAHcwvHfmL
pJvGLml3jX5sTSuWejXoKetyR86rccGqYB9G85vbp/0nme2HtMGJ5uoIpRu+1MXp
TzyFsURC0bILMzxq+MRNjXOPA9puXb80Ln6mTx+Lz2yEj0CsCno7wgFgmKDcydCc
lSYTWik10P0nB6R32l5gfMWerWo9dYwlIYhEdkWdoBT0RtPd28Ti/tJ8QZJfl8YT
Q9m/w9mLks28ilv0WiIQ57SE3S0k6MhBaAaKW5pvDFHi413iNuiuvMLuOONQOZY1
33IwkNN06pDbJEdqi6jOT5etiCADCJ/EPOYtW03YbTa/azu1Dh7l3dTsO2w1CeiA
y815T8ghfIdIbWaZ3mCcf+ssOAtdOccvO11y/2XR+gbQA0UwQyTqQwbZ26fJGKA0
9CNEufkIoOsVjDJppjBT9E+l4okHExtWyjn8bMXtd2kuAs7LTRGOltBbAFxL2/uK
n2IqlhKD2Et1kFt6MwJ7SjSg3rai+icI06Fse2JKN4Z1ll+mtsrN8u3CRaHsdU1X
pyYoG3b4iiRed53RqZ9CqB/YvvHakmx7+xa1fnmRQq2L5DqJ1XaX7Bd+uzwA1VB+
o+PZOvDbNqaOxXEpdY00+F70fOg9OB0C295HWC/hvSlD+IXOc9bYEJEwAekKFHBC
1gvLwmfI0YlO7c0SrglpkSzqKKioeoUrrnX8HmK+YN7fpuLDc2JY2/HfSI6jno2J
ZwJzgX+58Fxc29XHsRBbinnpE/R6qcc3knBkfm/lvy/TfM+W/dnt4i20BFyEndG0
+VJGDgbiFXbN1h447yIsJYfcokImfoH48pkZ+z5A+cRP6Ork74pWTFHeMb7hXubp
ZXKIZYOwA1zGZF5q8638gU3RewjQEGPeoMZ7yLcyud9ObpmqJ4OXgZl97c1JQa2R
2dZyRDyH93hv1PWhd6AS0iYD2B5F8D3+h9O8/WTxanba0FpyA/aP4y70+ZmDWP8v
yr59mvyNhO3+C8ausR/Oj5FTcvJPH/QQwvkcUPC5SLjh24trFtKLWddZ8DJTWYdT
MvZoMvQOWVD3qwgetYfVNtNELe36H+m3fPITkoqkH2dST7Pu+J3zvhlQWOcDOmSD
hOdMo08ylXWuiQLOjeOwZqEtAofDi3+b1E7HVNZYxPOvqUlJZss/g44gY7YFWMWc
NuxPPdvJsDtVv0SgOzid8Ofsn6xgB2rmfnDr3RqgmwpV7HQadFamjZURxNvkWH5U
78vhkpDCNcFTH9z/dMj1PHg0zInFCht5yj9vBMal1LoXdjBFTNM389579EJICriP
yEu9gQJZqXbOYhwF2zMIlCTfyzO15floXDl5bE37Se+re75a1gW1kHwHnF4gO1/F
UbX3EWsbCrvGv7uYyUzK4jEFneZVJ2bGnU7ptuW1ovPWtIjpHWdJewy5YfG4oQgj
vFsp3gLxRAFQcPTvrZAr+NpypCMTP3YwypI4K4GRNLZ3F2MKQRnpkF70U7oaeu3N
hGDA8nhUewtrtembOdQIiBGWxldcgywjIM68KFku3vK50qmhdMD/UBt9us9a7N0F
a04KCH5zYJr1w6YpkdpG+TaSMlMgE8PZinRrHEf14qHTCBLCi569iAVUCJswa3RF
qDrxgs8m6gHsHH/9pnPpxhLiJmGQoZbNfNcKgVPuzxWuAWbggq+h6ddpKgk0Z23R
F8U8c/+WO+KQdIL376xh9qXeaeSXDPgJWXKTx4bnPit0yTle0gmeH39LH1VHEyUN
fLjgp38zGSREBq5MuRB4OFQtn6XPIQxbxMQDMyLQMAlH5es+gOO1PG18I0ecbtcg
ovwBWmqgNJJqB0gYpPslloInCTvA/vtQQJFrqZDm3Pv6u/Aon2Pu8Q7ynrbnybCe
ww53/BGyXo1x/aWXQFpQJCSxFg0BJjahJTSOUcGXNFyttih0WCQQbgP8Qq+U5yX9
XjChJXDIsCfbhdyyxQrRXrvfd47cZqb95xZWLsOpBoSpNJv9IaKuhjGAt/YHmN2T
O06Zed/d0gwVbjv7iCsd44DtpcbRDwLkXWMchA8W8yDBIDn/hYojx5IkbEt3RMpz
65g0B74OyLt/xVXYrgUEXcKpZw22NkmmG2w/jJ0EGsHV0YnDz4AlOHQ0kEHV94ds
pKqyZ2sWGYiPgutYMbTNHJDdFR4CRkT7dF5y2ZBVm0tE+KKSIbTnDGjsipNHaLBW
4hyeoHm0NIWDOMvsKZCNpjIu5L1HfLTz42od0Lr9+FVQoj1AuelC8izpW+pG7lqG
bv5DjbmOVEumG+nsd9xkBoHu3CVS7ykrn3YL2mn9zi+guEIowt06Au1RHh/kLwg1
qorLW4Yk9f9EqHjre1cBnayteDggeiwVmJ+xRGDz/Pmg5nmqOTJpiicD+bz/prmU
zdBzD3nGLt+PXHvYn+6YPmvUIk4BKxGT+M0vU5OMLrUBLvHToYjQvZhmfZgEKjgk
8SI18CYUbSyJIiajHmFJKJVq7MHjpVNTpxqvdRwu365+84Cv+r3mNKbB4gNf8IXY
0A874+Ope7zHZowvaCpP6Z/oYj3PjXFSb6l7x0uKskYn8rw76CGvf+gDhuWvH+rO
sBLA8Qaenw8ltYY2+u2z22bGt9NITAmOTPE+f0i1JsySayDzr255Ug4AUWvReHli
BZV183igxCxixi2gZSHtey0X0C8J3ILX1USRmPMqclRGrAUXuMg4jL6Y+dX5Cwvw
LqsgEXSawTruK1Riei7HkXSQZS7X8lUKnFsjjwCzlhcDGPSF9OCm0l3gT2Sux4sC
m1EwjkoymfvG2FE0f5BcclU43/exwYZb0C9oFxNu0k7lBmAbwe+h8QwBt7iSn9Ka
Jps3BWkX/cjaNmDZphw3JdDwdlMHnG0SSPwMOsgHEqyhlzl7UCuTPYqG8Oz93ZDc
+BjBLhfPSAe1E5UcsKI1VkLp8a47ZcxBxPIr8HlOVEq4Yf3mMwwm1MJgV8mPmDAw
w2vV4XsfhwCMC4+jY+cx0EKj4LH3IrbJxb7Km+MNY5S1aUhZy6wbcYjS8wFhPnr1
2TRBYwqIw5w9xYA0Tyv1vQ==
`protect end_protected