`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 4720 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/9huKRhRMtvnNqb3Z+UU7TahEoHV+T8U3P3ufru7l1O
3DlgtZzb9QxCbOjthp9+wDkjygH0eUfDrEl1ovhZG60kznglzR4+t/YFiU2WE5HV
i1DdLfnmZCC3aPl5Lt9cXxigmb/XC7tNMW7ozmQMSstBq/CJ/VEnx1H7rFjudgS3
n0S4NxnrCFEQ41tXRuTarmADPMwsnT7N+UihC87O+p1hm9LQEZsd0WTwpdsp6gl5
IYOov6lMNY4CgBERyqW7Kcm02/uHdAEsotKdeW7BVX3OXw7uxFMx3dZ2VaAF1Yp/
o3TJ0YwNBjpvzEDLsaFGci7T6b3bI3CiRMb+WG3GKb4oZ7HGtqKnomzMyIu30o7q
2kx1Ys/13wCK+h602O519qyRCNLBPY2r5GnwlC9WBOg1ALkO8reOgci4RqKRTW/9
LFrAo3RV4HNorEK8Ey2YURMwJLQHKhXCjv1uZtHPxR1Ii61BOznJ/YlojU/gQZDx
QDTOCN43Gez2rJQxCgKwEqImBxh9a3zlzCHBROB5EqaAOfIeql+78ES2TfqdkGnY
X6uDTZQUyw4if+8R1Nt9fy22IWIIS9T6c8nsszwqorV2rQuntDWbbi2KdubVHBWt
YHxGtsW1BYTJcihPNhfUHr+RJPLYqRXGat8NAjRMdjGxh1DQNT3TiR1neNZOPt97
wxBB7KhaJyBdiAATB0AnFi9ZkRVn+JAQIzcfLKwe6y7ramc0eXZDH9YnllCHTkHr
2mQoBU4QVvwtu9wWUzG2wvaHiHecztnSKMgFZ1Q/n+at1brF+9H9hTSEZeVcjPAi
b0fhMeYtuFIeBJ4TSqOgA4wj1I8zzv1nGoiglmLertvY6y0C8vW6W095UBKRGYjQ
MsK29CN8VtGPUJX6shr0aI7ippATi1Rm99lFgbFaV4L6whN2J7OdVyDkJt/viYRc
WIbsSuJ90IILl4qfEmPzNnNM0M9wCYN6bD0cas9wmtgRzvQcv6li55kMMPhRuy6b
Rd22Lkvpulg5KSTqF2qWl9HjRRpxpEPmD1K1dbUlYDYLuEGrpZVkFoxfPp/9zniZ
PdmUJ7VUdBNelRDZp2zgoPibqwJRGTzs6ZKDSKxsJZsfHhAvtb3VJTq5nJYH/Nyw
vJ6Z2Yi/lEVvbUY83duMW9Z/jPBknQOHRRmKNydwPsSIuCqOgZHCDgGrJaRQO5UO
CANqKRWXoq2P5Tj8bIf4PvVDE60xQZr9KP1SuDL5c+lNv6jW9TYJ3N7FRQC7CHo3
ldQljtN+sKWTX1QAd/m1MBaoMFoUaJt7ZIe5vZsXkalCacyRYhNrwIhOWlqDRvzD
XfGKmVILBpPi4vmHCP4BrmVUPC7+Kz9vmwn1LjU2O0sBx3Hyga9niyyxJYUFRh7X
yjovPBi3FgEj3+O1bmQAwYmfOnixxd7nmLFW++9L4+LVErBkD0FTV3BdtWV4tJ6J
VSqs2SwkvumLIV9sbAwQrMxEPgCYkTfeaE39y4U70P1gP+ihiJq5Z8+MRFRbGDg3
8qscEZ8dFo/aX36HSBJ5k2/ejviG6TOo2OCuEH2yas4RQ+2jS96hM3TO2+B2f5mI
UzYCjbxM3+9bzzpqaDE/3qLAC8/ntwkPfY5TN6aP7kbL44nSokZXeGVXmxx074dg
MtcP8233eqaTcDDgQIK/f9+yiBNkqhXZ4wsLedFBSyHcWDRpOSumlw4Qm3IRRBWr
uL3iwoBQ+OKue4lEhAeySRhEWAdeKRMR53pdbqTOTyJCkwcmlSLffbIJLrCPvQ5f
AcrZTpgdm2eP3DSZjTPaC++UTzfEY5krgxBqDNdf6ddzC3wfbGmtdmx56jaHeEJX
eGvhXhPgBR5vsaD50TwrgtTWGkk8zllhFI+KNiOKZNNdjeHR8I6MApd1BuToRJk1
xVbZSaX6EcC0WLuk3bdnS41A9H3MVmaflZxSntZgVIUVYi5YzJ2C5EB8SI5nVIFW
CyPVkfuETaKnYHGd2uF9T/dv1jYs/+nkY0DD/81rBUVBVP6Hxlhh95632ST3HBGx
BJAP9/Q7nrx1LTpOKnpXPrMziS0uCjSXyEQa6ORgzHYdUDmrwzAcFOlKQxHxNfi0
5S3aXck1817NKv5JO6S+nkdxMWgI1EAjZzosnaIaCJGzrR3zYzPbcZhOTaEvQgpW
ZxbNC7k1xM52hbwjWwpoO1hzsNTY3HvEBcGWZK8upG3Rj2aGL0edYOglc46WMJJo
xUo9YLm5ETAgN03ZKvcxV3ohXwa0VgarIciCa5WmY5nY8jThlnkqvkx98SLTnJT2
M7kNd2EQBj3TiHXaw1F9zCkb80qmxOm9gQtN9heBz/6e7y6MRuoiVNAMtqfJUTtj
BkYZkKWFYhwiZvS4RjkCN/C1A7JAatYbO1g+ZnnA7HPOS6Wmc48D7lP2C4jlQTCQ
YjrUyupByGRRyejEahbUFrPiKdHgebkuTcWUuddjkJbgTMwLtWFOCQ5apz1UKWMH
OuRc26wQiliPsd1mGpFKp7dnvwWNL6nybhc0mXyf7Iv+NI7EXaX3xpPhxYABaNt2
fBVyb83CR533C+FVK2lR7JgVhCylw9IZcHF4pfjOEoHv97NpgSmIDaI+G52+LQjK
6RaAq7oUFyKzJ7wge6j8oIhWpxCjV93/x59tElDnYGMrAPlFoXHDaPo++Ukq76xw
W/jPeC8NVKmgT9WweWPUMv6X8FFGAb8nsZ1DMzIlp2plSRv+uEFliuGjdReC3pFs
ZcCFqvqxLWxjsdJsZAK+nV/TVpbZwZI8sr2QUolGgxfM1uAff0go8crBvLiSVY9R
P9glYGsg19JgBr0QutibFx3LYUHXZeEhwCKJGUycG1BYZDtCXiyTfRqkfmoiSbYt
vOuLo6dIajKgrsnfmjidnouQVNOjX+GknUAdA2Ojc+f+vLCAoRnaEoYvnZIHFN1L
A6Qup0leJn3/NoMQjn3+aD05mfaT3kzhHNroRpqE2GnFUI5jNPF+kWN/fQ6JnQUJ
+rooQ4bVSq9J9Q8GrrFFddlIzo59cjxbvoUhFw06il96oFrMRNRUO8TtA4bGylT5
tpafVfOTruFnB5U2UoegLe1DS93PX0UelBuZafA0ZDUmyf1GU/NepITMc7NpUifH
ee6KeJTLynwaHe6QR7voqNSntxgZJ5h36EX2ajjxfzMylq+8ZS69sSlnlS1rnHaQ
YfmBEjMHce1PtIj7Ndkl5Kcmixd7iWFPLKIR3C/egMTeUzOn6Nnsdlpkdj1og43P
dbYpQjqwxzX+izotpTUYhiwgOeh+zObplSkDLjlaplIDenKyCvOy8fVVro56leH/
hyncLdSscyyip4PrWew2yo/GZoHdtM56Jd3/GYPdg8O9GtpqmrHmTxGSAQJE6QbS
BloWf2x84ImwUhVQ7wUvqBsIQUW9zDPlgggXzhSN/OWv2ymnPyvIGsLm+PU6sx4T
XXC/5Y1tNHjvV2RjQdFZubkQBvqTz2KpsV2VkdJOLMh+tvQJdPcxvCXyvouG4B8E
vXjW41nHwoXTFpK7A9EX1p9M+OCrYDYnCV7/0OLwB+IGhF8GXUJzI9jYFG+1ghuS
820fFIideKxKBxt0Dw1dSinvEcTmr9ywI+uSChEBAD1jAr180Ca72dR2CTOKPrsY
pj+8OUWT5MAV10IDxXO62JKJjh+KkrGaSlMWIHbCQLQMV2/3dj7pSWewcXdvmIFK
M4d79SoRMGLHx/rWMbkB6MxzBcmdmhg9hQGOlSahhFcE2hyV51vOR0jOwCP6Hf1W
UROx6qPCyP6bPQeYfqxfaJADLZMG7Yvc9rM2nMaQnSrX3aD38OcgCtEJTJSmjDkh
WrW8nfD9vQ/JLp3LUv6RhQKdNJhgOMOPKXVk3dY3Iz4GxMegYTN6DDwIojzKAyzp
7veTjTl/me4Oo3sExvobWrs78chT9yC7SJSuavNv+WRSbHkpjoR7Hgn9J4RMAvDa
cGhQGrucCRuAMcBlmQdS9yGk33cSkHArOfdTk/5f9Mr4ed8VN5siwZKRtt4QYqJ9
AfF5oRTQLqZk4vauGHugk9Gsca3T5V67jAknVMUDyOAlpCA1YfOGqzXOjlSSf8mU
5zh2vTeaINfH5/N0y3iMgXouD7bGG4nKPfTVSGWVwbHoIjPUaC5GdrZkGFJ3sO5h
kdX3bxMjJwrzNEv8FyhE25ve6A9qldODd8FE0/09P2gNUamrJxeWKVGl7qEcoqzB
0YsdHxrzoNp15VC6apYg2k3KZJiqmNG6AuBj4b603M9koQddmPa6xvsVR+BUaIIk
zaTgYYcKM96ZYz5Dy13MZHCXtSyxTwyhlBv8atU02elux125tDlpS8zPYbF+yQ2u
ap4zyUCAPFNEQQoppka6wjef5GkOewsudl16y8IBoV8gUhJS0vRMvW83uz5UgbYL
RL0bZyOCuRHgM81eXaUgRKw8fSrZ+pDNLO+eh6vCyFacktmBzXi8eh7S3ejL9r3+
ULzrSamXj3rIx0TQUD67axbf8/UoaVK4BwuzxEyt6hMyc2ZGdth6FjdxXizUq8oI
l6fj7owdwD/IJ0QP41Fu0uBKbPa4uQtoBLv4St8So1zI9YG6qDojIiNomcWytL5q
fSwzqNaiKtjYtyZlggY+NUkp4JP7FfORbWGbtf1ATznXbGqgI2M7MmjYQsbqOWok
Ct02zBU0BQmgKGaXhUtNo7tZGVs7zKKGMqEworQWbuSlWUiw3IjRRpulmfTIJH+E
No/2WfYdiHhIHnO0iRmzAgHnf5gEL0QHCJ1mPkIuYf6zFbwPLgS5TlZMMNYMb1/L
C9E9Di95Y1BeRLarhmMzMB1oVPeL3o7qXUhqgJvy5VpSyMLON/Bxko+ub35pc3lG
5Krdcml9OX+M/ckxUit9INnqhzSRPINaLERE7c3XvIyHxFNqI98H5zSX2g7K/Gff
s6d4cYl37IYYtf8RoQ7BJietQctEOnqfPfwfaJLuPWiY1xv1JeetWI4KVhiQEsCs
Enf4s4209WkMaWkx28PtqJfD9mYQXlWz4W9/H2lKfqdplulzVganc7hcXtCg6L0/
1r8cPuJHbHZbAYMCcx3a39habqbhfvLFNs6aQ+2T/Enm4IjbEG1RAoIccev2ONoK
PfBtUyLZUnTtvWSwFp8YQUhWaQHyg/R7JpHln2hBY8K8qPJNfkWiMZblR2pphBap
In/GfmngP+Vt9iTfBllnyt1o/Bt2GFyYHTPiWRv8f9Ji+OsJpDtrwwSAPI61q4F8
mxO9ryHxVubT/ipm8ktS//KCo2uBQYIESZJp/408ITDPIfCIWgM0KQ4sol5lMwnm
QHoz7MFP3Kkd9tAF/gwMh5VBgBKRtgg+8bvOve2qsPXPWprc05zK6iMFhQzQ+g9A
h2DPCqXY7sC+oaJnTBvcAUezuWZGniTZOUaWXzw1+9A6P8ClZKK0Cvn/FFYGC1Iy
g7oIpI/WwbroAxVwGQQEnqce2UTjiniCDiGFFqBE3xR73xd8WiIceMhY5Gf8FHae
MbSgvEXSHMwESLhMXM1I0ND8lkwh+5p2TrPCgslflQFtFQyOSLvruOPHrY+dQLxA
ej7oMKH+vKeSqzoLCSVHG9SAVlZcgIjGR2+yHKmpqcIxu3Bd98/NijAP3ZvPFHZ0
j7yu0snJFc3rsNMxsGlGEk1ILZJOvWWltuUG39c9gNJYe+7KAqY/B6lEqPI8Q2Jo
5RgMSjN5MX3191KvpRvlu2n+q814tuqZjmag5IOyDIcBQ5YhEjF/63Hl+1X+MxJK
set/rlDmPcg1wmFk7Icr5Nb8909flPNCiT7rvtwzPrPF6MvaZQ3OG0OoZugKQhUZ
InFA72lDrVOl7ayNgyz5AGlxYFaLUoHUqxayH2UJ5rLsxPBKy7GlC6lL9SR0od0T
WEdv+67GrNlbA2oEINVyMrDG/m8ddf5df3Y32tks61qh5uLajil8rbThf2izB6wV
yg+ABsNFBEwiZyWX3pE4M25UHHtCehdf0M81ArrIYPZjSdBtQ6OvAGklqM9/L5La
QgQZ1Rc6zbiD8WPtuLF6u2dGdsXkZRECkHRDapwFR37hK8XLc57cz+aAqQ/Oj69s
MHUaKFBqLVZxLh76wvFvWmVr2Y/PIbQVSIpsm1C6eYcVMdNtZNj+MomG221amlGD
7vWLm/WmHL/CizvrLQSHkj4GvF5dQ71lkPJehMF27GTFaKpnLEQ7wPRBDKPYPqdx
zi/adk8X4k0OrtbzVoRBgnt4EUWSNec/5wLu0JZ555DTVZ9W2P5h5ZTrNtZ7YW+O
0zba0urOuSoVAkoOPLANCQ==
`protect end_protected