`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 4960 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/9huKRhRMtvnNqb3Z+UU7TahEoHV+T8U3P3ufru7l1O
3DlgtZzb9QxCbOjthp9+wDkjygH0eUfDrEl1ovhZG61gsVzKTOddJNhhskPlY+A1
nj1BQoBmSx8LC+TZFwgcPO2Yg0hLfq1bJnCGUcl3rth5KZvdgnACgPjBtG0IqV+g
hbCtlGcqgjJEbAHCFaToixfMDVdN83z7OvB64wuglLqn8rPWVgz3c9tnVKBsBnt9
nj6uaYnn2cU56dRtMqO0994H2BeOIh4h+UDwQ7AvNN1ivBCCe2x2hX+rR5EN1Jyn
aNT5KuI6iGElz2/fxtNwU+Epqgc0K9Ok3xrObnlXUOGvUTPA9stVcFubEUYC0J1Z
QhIgtEOS+jaEkEuaqaT9dJOOTfO9/4nBn9V7CQ9P/evlUMnphjQE7QxwA6/Xf2dN
eAJsDx2POuG58P6ArdN0BOkiVYx8ZwytDHfjEedqYvSQqgxpcrJT1p1XeGdIy2R2
VJn7PGZ3p1mFuXEQIvRZADVMPdjOgkM3xPEI0S9LZRq0GikjJ4X0YvRaGrDObNac
3JPhUV8K8q5852mpVjca3tSNFKGzhEQOeCE4MNAslBBYw9vw2+AmhpBFokE7hjI7
Rhlh6NuhQh9aV0pxCe+p4C2pXeaYl33tAyb/N7NHD5okcXVTdi/x/ffkfDdORBZI
H5xezXfWgQ+5mknS/d7k1e5HKoaW7KhYaNOtlIa+ITsrhu2aJNL5U8JTUs/m+u47
xhHCtBnhtQIxm/Wcb/4i/FoM1lazyPtS5MwOc4YUrX/fVSdotPCTK5lW2GRmqSg0
TcCkmiGd8/yc6cShA0b0eoci+fPaiFA2C3gTn4cCNWN+D3qYJTHGsyRX9CoeNslM
I6yPHbdybfrjooNJVZYzD91fIMFgqjLH10kak2S94oK5OluesLo5zOc+gP/Px+Kp
K+XBlMPExPEmtLSRkSxUGqEDcd0rEy73zu2EcE52BG55kloVfu2sCY740MCCFruL
TiO7O/2RD3nxMnbZvU/8hgt3pcZ8nq4vhUxZFYRmFGAE5Lhk6zFCZF2Q5JcZWAk0
g68V+nM8i2iGTOGdtOwZ8mN8z1EMgyQQg2rTBOx5Uef1Gre5o8o+rkEZgnQLIYOE
yfV9j2bfTeHVwn3kd5T6//xodWw0Q5KeWuHkTsKAyaSXV3eaizl2NwQzSuDl47It
IZit7Dy2RNeX7U7cqFr5I+10bDdFCP1EzUg4v/UarNBev+03um3Uku2+vpiA+pdU
V/y4k9NgMz0Rq4KZ2CPcFFpzCOUN0MsxPy1EkL0PbgC1kAQr2JeBVUdC1qN/zduH
AxYH8yez+rUMrCDPH5LVMx+sguo3/IBzdCjZqdQzG3VN6qka7grCVB6vhQYCMriY
pbRatnxMA63kazzxCWJ2oyTzoY4LDyDBqIVPnyfnAYQyz+Tjy29WNAMtzy46JXif
upuYjMkq5r4oMQoLjXdpCUxurqR+AWwIxE8oCJnn016M7cZQzDD2qw9GAqFzrdkW
E7TG4M/g7cN7CM6xWGWk571AuEZmwDd0ykvxyk7nXh5WlFEkhMJAkfJ9gLsw283W
TYJYP0aly9gQ0LlIBWMWP8ANvHCcXxJFWSwVBLuYkK85rnctuwLTFDV1Syy32USk
UxDkI2G76Tf8vUCmRW0sjiVJH7ktbRzoOiCnFLSJYC+K1/cGtFsrWUtphSu6IbOg
0bNpcjSmOZ0QE19xT73jsWceZfg/quTGrRW0pgNm1j8VlNvwjURMeprUmJSyhFK6
xTc/15t1fRMBao9e3p9R6iNK2k5LGsesn5txR6WOlwW9/3rjcMOeESlGbKIZaAJb
le87Ej14lhYuyDVKQcYKGgAwEHypx4afa2MK84cfopYlFkpMPD5Cq3HcV6LhTfvj
TNFXUzqxCeIvHHh+5qVmD4SGdtD4kKUvVkKihap7Bq+SOBYMdckVSR4MHZhriXK6
dn6Zp2iG59a9rVvNO+DxUg+H5LXqsrl2CWHsFlm/pN+lIkPkbpxseeyuXvDwdEgp
0l2ZgKpX6u0tBDd/1C1ZprQ+FOSqzrxXhyvLzSki/b+kRyvNc9Y8q/czTPypvP+s
T1ecycXJv0QzeeDPiQnkC78lHWrYl+gQd2mD63QeRnK3COZQ4rMDGRWm6w3eVJCp
ZiYHST+hHTwprgZl2/Ld5RD9khzUBG7zhPKu0l8sKH7si9QNRJWr0wSZCi0tl57q
lYvbub7WY5+lVl1HOpHMHb4iNvAmSfzkt+EeGMr00Wbxz7FpF5us0S4yQeo6QxHs
MAqAsY75TLhOCmXdI0tEkRoPSVhM4V2a9qCaIL5iCeOXMCC0K8X5FtYUGiZomRHb
rJC3LQ1nVSLQG4w5yWK0h8boZWZG1VJSBZ8FRkhFUpZKBPej+llAlRIrrf4RofsB
WjP6MOvv2Lp0RKe0JqzPQyxzNJJ0KgxTNBjrbik9AL4OwZqasZaujjTkWghU1GTi
YJaI9W6MLG94Exa0wi4pBvtktMiSvOy9cFAPTnRpPsF6TMBOPZS0llYFHxvkoszS
It6NublSLclygdutt7igJ1mdEgJ1VWCvyX2FWCqgUBqXtINkjcVmI9enscN5oh67
3Im1oZO7hQw89K76yRrVOIyGuLcLOy0O2LdzDFOTWvpledj+BvSPHmOYUqkGZDlO
CNlRep9ndykA5lxTfbtTtStnDa0vvAkxtPIFPfe4AuwG7qEWHGYQ5LAePadJQUxt
2Lj/7hhngslZimMDj0f/gp2imP/8vXFNjoE/on6rFW+3Mj2LEd7ONDDxBf3Ix1dp
H6SLcSqjjxRbwnmFpmKmWr/OVHRJ6d823Ed+MOCXNNihwW7G73pnq27HmJ4EkWOp
dlafqSIPeBtWZ3zjbVw9dOeQUF3jF1rkmDxhr8cWDYM4T9lxqR3pLhLQl1Dc0HT8
g6a7EUr2EHumgNEn2Yi4CyQ6MPxpg8lnKy2DZBc9N4JRYzhJJ7sh0pwXBlxfDGkw
2QCv4gJ9C5GHWwRGOJjULjJu/Ibag1JMS/Ulub+C1LCbgLo7wsXK0m2EQ0/U5Abq
LmsGCQ6+Ymnn/VzKW2sWRgLmw0kOXYbqTjKoRqG3UyUI3JMpwJuw0EKPg4/+ajJU
8ltXUzPeadpWyxTSVSxC/e5ovLNM8roDYGKTTtoqSgm+k/XABhJoiFFdWeunWmrN
IK+p6LZimtC3G4PIvf/4jED9vbnGTvX/LS6d1oNSwCaufXKMu9nDTWhe70dyGytn
2Sft0YxOYtCpWRJ50PK0kAZYM+EnZ9TV2EmfvDWtcBxplPQGDlamrwg7UolpePdE
1F0/9tFQWIhDmHQ1N0D6VDs5FOdt2tPRBpHMZ19DP1Yvm+SIqI88kNibGq11FKao
WKIUsvykZvSek+XyjWvvz5hO7WdwB9ptxfQk63mHEEHXUPJZAjnj6s9x1IAi+vUn
uUp6khNBpxDRix3JD2xNzattlAra8rOFAe872JNJZ7i9sohg98vcNM95/DxUwGB2
Mh2c8gF3VHjYcX8OIHdZlx1mrwkWZ95oUk/86sRJV5UZE+9kW+8sEQle/d16SKrY
F6tBX1WUfrQHXJ9tmQkZYSrbNN8TQQve+sJ03LQzKCPDhqqYLkzoFhheBn1zqpd7
oab1WWFMpwjtoSBbZpcAtnqokmh17UL0n5TvWaf8pX+bqAKNrHD5YH2uWyN2MDx/
8JqYiqYyEpuQfUjv2rHYEur506G7hIyPhopnoWddlCG7E6naPsHdryVHqIsS0LwK
E6YY5cydQa8L1CNfK333hdUbIHwSU/eNDdfALzPnGiz6BzAktj3MiTfP+MR6rHx7
mnJao4HNfOdRbTqr/naUq83i9xlQByMD2VZ+6RRaLtMkyLxOSRpl57+Y2PPxF8/z
twdPRHfR6CjX4bI8fldnjetuWxwX1JzMoTacX/YVnwziPhYI15sckQzXpDQEKbkf
GDocpc4TlKXdvc8t/temULHjeAnJBV6741+WYtcWUNZfXOaLfoXvSx5gUAwwVjdl
SteRR9wb23X7FiN763gK85jQYo9dCHFHK1CAmeOJiruoFAxM4XuqhBOtyKW37F55
2cs3KDeeOzT3GhrmaYJWCTfGo7+y1pjonzp4TN6e6uh/N6JJvsJ4cchJ+80d8Eoq
F4UiRR9y2wpV38j4fgCeItk5S8Qu1/a7jtfDFdyhsdJauxTBJveAD3PFQNom6b0x
uJUY7KthIFcqaCHNW1e2vIWgNuV4vCtcf6MkKwmcJIb5CWXyTs5M2iSfHMeuOgb2
sfeYrui+lIIfOl1JqeLAbMNRpea1BYVj3dGtiT2Ifran8Mqeb4CXVgOZ8BkpqfI8
auyToJstB705rkwqTL/4Rn0oxQ/3MNDiMnKncKDk7MFeSQXvqF2ZKT4D7+LgHT0U
9lkkvNDyjyMGGK2sO/kdH9LbCpp+GuJ45SFTCjgm8ZAjuT61yBHZ2MjRvWlL2y5I
Nh9JI1S0macMe3iIEJy9dVwNrEJTiByYN2xBXgZ4/CK0vl9O/fZ2eW9IFhNDBWfz
t0+SlTT4iAy7UBG2ZLWU1f5MIlfVbODt5GO1qomqXf6nXS6zba4fp75Co+cdXAro
gPY2eWIDcpYlIXwqpOvXPTMimGMCVhMondBAySrUrLeCzszAz0iIbv3l7P7ENLpx
VV1T0rS+jGAiV+k4K8wqTUDHEtOyn/se4T4Jlfk1YlUGBleEGLEVifv/ZHs0b1MY
qnpJQ2FdVHqgBxSu0DJ4K0vJRidhAvhHYfyK6TQs1Alo8gZqsnB3woLHoD8e08ui
N4jAA1MERBj5WMbgk21N3Naek3WELdd6B9Xsbao81pC9LR1og2T6MmEQGbhWE1Fb
A94t9rdl25pVXdu4f8TRynVNrPhFUcaHxyoqhA+0FVPDaWArHkpCn8IKYxA1Uanj
NKsNWDq2maDpoGWYTj09eghjnkZNd4vGQSh74qeVed6+nSzWyClfF0M45e4XyqhK
sTBQEZ+cB72JS55OXym2rb+DdHQ4ixA7LeZ5Q3JKna+PS0qg9iMkI0BEvzwix3WZ
2GKYYC24iklGrslWKecAe66A+Las0ukJSZbGHjXsBaAFLraseUfZ5kKa/1/vqLqJ
Svah3HJ7BlCvxhxRIjp/Ukc5JsLoL2IyKyr11awJR/26yg2i25bCFJcLOQCZT9VT
YRXmpsb15PRgzR8x8tIu5fwiXH4LGEeWe4Ss6QKx8Xeb8pjRfew/cuuY4tFqAK0+
vaCIxSrd8KqKvPR01xpf+hQ/aMwtuATONTpWcYVy82/zXPr5V4EqgVbdYKmWZjWj
d7zOvI2vVHcxxDhm+Ea7z3DfzQOZnTL5pFhhnCd4PQLEBCrgXAy2quAdzozofWlz
AurKuB+1o7TXUFZmunoRkxsFTaC5R/+TDERB5z1yS2f8DrNDoQGhDSXQXS0HvniI
SLocq/e5Dq8ZLmJuTeqC4YUaUyikUeBB9XWVKBlJ5HdnYSYh/rSOSyHItORPk0xr
47E9FcJzhg2lzf9WbVO257vbCOIUGt9sz3AG4BOCbCSartXFlKpEHKG6aBEQ/oaS
5wzdXAq73sUCjPtjuQiEU0SbzXyW5m8Zmj7J3KTPr22fddy60X1ZOyqBN25EyD4P
hJMCoTA02knrx0xej1QQjHA9hs+xepvYDbBUlNGK2+h9hrICfFnOKC/7djPp5bVc
MhxhyHBIKgwR3Ra6bd+kEgj+tvzL4tEK/mBU4KTAEoIgJkmsNBTJ6pghI9fot7bQ
bUYbQhRbmODMzdeg1K0901lX+f2HDbmtnukOzk0f8BfPk2l+GFmdnNde1Kd1UN24
bXYfsHSA+0/pnW4E1IZ9j6ybGdce2mYbhdGrsBUlk3KJ0c6gZQTUcPYFPlSMLf7T
l4WARDOo2kkdyrAjtNm1bKNnG9pGGSOhbYuXCM0lsRrKy6JX7sw7/ZFtsVjw4W1y
+VMMiNyPzk5jV970BXlITPa5jyqXUQ3AHTtTybbxMoCnUi0EUcnf0sBGCWeNXj06
RPaiYrqAEKwyUjS/qoNF8KOluXlvzq/EcmEATPC8utRQvCgwhOFNJH0xPznNSNKd
Xo5RdlrvntIN5KzIatrWLIddJkNm7cqB1voGs6aK+RqsgKYqAJItKTxoGog1MU9p
sijlhYPD2SKcH7noe1MI4TPvVvbNAPmoQnZQorjhAVy/1/2ohsduQqPMpt5SyqkM
vkmCfXsQ+cs6lEpN67RziqFW7X4KFulKOMPOKa/uHJsAyl4srpn7qHxshZNLt1UV
vSQBwCBrsS9mJGPvHeGmwcGU17WYs94+DxB5yWg23yMSNB7GcU8mQJ6rTvSPfbRC
44sDvuz6h1oK8SuC1yNq5rF3ZOVUxyufwXu/oOiL58n3m5F8dgujelcl556vAtt8
GMC+QJvtSQZRQpO+fEW89XGWcB6jSc8PCzssfSRO9TC3MdMk0cqfsQmbSc1nPYE7
5mLeu/gJ7t0Bu1YtNQZL4xblSzbXVXrq0V9Ii4Ac2WMtmhqaoO8/AB1d4Ho5wqeb
v88c5SNxLPFCxznvhhQO4B4hIIrEBaAGUjjnZxDhbqcssxB4wVcNTxsLt0FFpppJ
iDQcqbwLfjuLt1r14lVfIA==
`protect end_protected