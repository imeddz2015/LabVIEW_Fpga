`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 39008 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/59UwEX+aE7FohaWu0/8IpTj7mav863zUNIsgIH2BWb
Abd9opeuBjbGF/waQMI2vMJTwD1ie1YueHc3nSNpEh4OXp8P5ybZFY89uyGz3ztU
W1EsuUnchJoQgbHZ/sLbgtGRgsrAFn+ZoIeGN1d6RAF2wAESJmYP8zw+p00RvjZ5
cIKFp5nAtYJJL/0ymHGZSK2KjvdjJ6M61U4yLtrKI6fgqm4w4pborbocyXIo9UKM
lrWHrkjpQm0ucEOSpj+I6wuNhTV27GexFnr9aFojCSASgHY6tZAW1SHaCSRlhKi4
jBt59GkXiO3bBjAL2A1f++Oc0y88KhFH5qdGLZ1hyLP0LIUOH3IzQPPOGS1PthE8
JCdAFFvqIPUGEIX4lpuSqKcyVvW8IgjodJLhvj6TnwUlHMaRqE4G6XXUUicsTtDc
1z74TutfatiKv/457LQrXDV2CjMLzTUtpTBYCCFiRuiBBVq5txgIacK8D9/qHhed
Z/+A1aBS/w1S+9u+bYxZyuQJsIKaAM9ZFcKn1YRZMG1G/6WFyGqyaGhXD+pr8lTS
pgsPs+N4gLSdHOnIi6J38I+oaia9zwgt9gb0/Tzd0vGE6X6MXz2R5AV0cFgyTHvH
5yulvpWzgAguG2llROkCSmKKm2ruTFhCDLwqiuoafc+BEThESos+cfrsYj3CpDl7
kbytTRj2gEZu+Cq9ir64NvNFi7ZwMxeaF59CSRQ7vZU/ksFGljItiTGpM5tTtKCr
BJqQIfyaB7aPaSwzVe2RI7j7pmJMx2dxn/HNcJ7aZyd9nJmwYIH1OU8Y2MeojbOt
1Nk1SAMN1OPni5EkhSGW46ZEQ1ap7+hh3wX/1oZl4KOhTtJbbNYEBgL4wx2YXbBd
PHZvaMCQVUnSzyrCgYOrVTiPUAdRA+b049cdnOS/zGdoxHdg74zWa4PU4anN2Rnm
UCUfi+ZMywx5NXzhEMFa+WKUfYWY0JGzlNFJuTnFLVjUJboP/RvNZUsAIl8TixQZ
dnJdrkzoRkjAYS5kgMJD2jofvCMfMgR0RL8He+/Rr8USBp5JUz2U/Imcxgei0BcJ
bU9YkN1TBXM16Wa8jKNLmBCZgd8TjYw4hbtdrDBixHIokwPN42BIS7QT8soXhACJ
5BpEwrke5pELjAI0Duq2SQOxzOO4kXYjNes76ZcDtxuyiLgkwBx+2xzXXF+N83lJ
oS2glMeVOoGfbiGP82t6+VY3bq+XaEktI6rBtuZ1cmEyQ+WQaITOBfblFM16yVTl
BJyT/xs03C8w6PKuhvrZo5zfTLDNmYhjj4QWue73LEZSSLXq6Vy3ed4vxh8MTr2u
MutDtDNn3SANxdCh6KcwodkGy2J4EJ/AclU6v71Fm/AKtetEw4O9Aatkzdaqql+k
SNZrjKkYFGsPCMEm0O3IhgYk92cTQXNm9Axyn3C/OeJFB0r18UVZUrD/jQ9k7EKk
nP+AxORCX1Myubpz9R/EG7oz78khPzgeAkZiq2DspPR/vGXmUqEDzm8rH46jdKXG
Y+OaWqjJKSXKe5LAUyYGarszofM7o3cgwN8wY6ULbhbKHNUxTXXrOuoVQ70dkfbM
i69VUiNPIWxXVAgpv8DumzgqXfCgor7e2oEQiIlsGpauheNwQrl108JRhwTGEc07
vJpyZ4z/GvQNK2RjsvfcYxh/nrzME/rD6D4kkDZ597OWFtcjUHWS9QYGiM/+MeiL
BSkGWFu24PTgPLrPpsuObZ0RnwiexzLz8P7lwhIamaerjpNsQ77BkMKXfCVbdx1s
sJUIZ+yLGwN0SD5GI9YK+1vnPp1RP5UGJl0WPSUD68k8mOyZHZ+N14uAf6E5xoAY
fC3ocr5aE/K6SK7VJL718rAGTbZozoug0pEqvFjyf20JwgoY6r85828lc9mNL9oK
zDlluyhe4GB9IkZpF2syl9DeeBVKvrK4Yful4NOv6/tIKQKUEZCxPgp/xXa1Vagk
P5486mmW92uOAzmQkAwgWInlAOHkSe4gPaOHfT64mal9D579Rmehj8n0n+2bRaBw
qnfdzIe2piYkqlEzRUWsycR0iSeFpboA82BYrYuYirS+6AAt6wfr/PG+qgr00Lvp
phYRtyJXM9bB701qM0+ovYkzgyoJFLSMfucHduoGKMscs3yHeb2OP87MiClWYazV
Eap60/d1eu7plTwMfTIAnGb5smhI1ssSLQbWNH5KHs5ZHcGVKyKKO673z2POuhdP
C6qs4YBQdK33Ejl9Q9K1HEe3yJgO1a+SvAaO+pMWA/n0XB1x2x2bXHjHovxpha7X
j6uImMsC1rDh/dvy3A9TqQppSdeKfzE8nxfRrr+kOY1LepIfVM8nQyMGhkk7ggDb
fK1JmoHw2iO47aXZrIQLUsIwDkVsLAtiT5JzPRnPCuvvNDMc0oepdR9JtLd7j0Nv
QhyiGPglHVmzSgamUMjidG5khN4rshAIUeisAEliqu+S+yuMaR9tLB1xVNcafkkd
qj+e8ca5Ez5OnSfYyxNOHsbXuHlkuK4EB3nKahOjRt3KTN4Qt5Z6SX8IK9pKOiHE
OZtUu7veosKf2uHrPXzjhXT+ShXmq3t/n5dfxEwewjQX3cUMjJmGqajBLUVvC9az
ElEhAFt6Gp61TELnGRDD+cPSYyCnRm6T5hoV1ZZ8NtHi6T/XlZIjGfgSjcP7rLbp
YgxJxny+AUuSn4twOLiYal7Ixi/3F/t3uUrDizdJOV6UKt2q0SDOSuatp2MPL0z0
nbw/zD7WOwVsrWE4mi/tBxmzbuLX90+Hn5J5IE8E0ASmyN8yYqw372GpHCGpoALo
w2X4o55gKZxC7FvLD5T5PbZPHyRDqPDX5JJfECSMpDgBPHh+AXDzrzwpgRHBxfjO
shoASL1dJEXxeVAw2wFGsF+phTvPsx0nXE4o94AYhIvsprnJqwbth4yTjToryXgN
CbGkaYCKIemUvvQCK1hysvDlRmftglodje+4PEvX5TaYeKH/4sOa0iahs+XKWAKd
2sy7rjZdatJ6g5O8nG04RSc2kgJHyxufZQL/b3fqIid/AMj5BSRRMnBzcuZl85oD
G64uF/DZLl3rOEAAYRZ8CsHemO8wH2HXUtnK6MMutDvCBvf8VKR7UmL/6GRUKmul
RaJ4pnfP5VFGDQt6iJ+MoiVxBrzU2dwx6pKmHsmxrBaXaLui5i7udeE88XdsNEcU
n5mkgeVIA4ViJuBf8/LRawRivqrrrILZfgFUdiyCGuc9nOfC420mDS7Sv0+XcVHP
essNfhG1/Fp8KMlIMqkmnWWnyj4ueNHCOnrkVDMi8YyzVbdyDuv9Ih4L0u5+l0GK
/+/qU2O1e0hLPxMgMb3ts6ps7GUFYidCJybNTfMb2ZwqT8GTb8N++hobuCKyVbnB
ffncNHNDpOOdip0CCmoYhgB6AtiEuv4abkGpDc4lA6GxpCoXi4ufbMRH4esrdFmI
XKdYVJo7gzLDjPkAU4jwvh52rpjZ6hOyDy3ZYJ9zdWXOaWczY8pjwRZUw+Eqn3RE
ftVjKRGitYWtfq7OyOMMD5b56WF1QgdiZo8ZfbxtRAbs+AhU3Wrqd6B1BVDg0UX4
b7pQub3FTUzD0bUM3JFsaIGdOIuYxJs9wfPAEk2kVaEtXpQHXwEeQ9x546Yu1/SS
ix1DBmccwR2+3INK50Z+ipksjgHlQz0ZRvCkPzh3tuo1j3SKhIHizkzwVCLSc2N0
WlALyK62kR0JTkZ5T8LbEAoygYcvSdXrrkYMis72hS/KidIrcsQzAyMgrtiu0r9P
QFmD32XsXdJJ760TsX2g7I3UxRTMhdUJSXVCGfhmBuGg8KUxGQJNe7djugTI0juL
0pU1bvPM5nWIofDPKkiBYCYrzTarplVAYjApU76/AFdEYjHVvwzmYGBJaOJGobhN
fniuzcxKk8jm6yyEcKFugUVWo7R1mixSYN6cprqTdYX7A2Bd26awipVDBjQR063c
lzTr089bOvRoUOOdbr3AM9tnhi4dLZ/3ZPozCi6bifuxgDsWq2jSpW6qutz1SBh0
ahwzLTi9c1vf9vA/rafFalfaKbqzOP3rxP8pNHlTeLh8Rkj4uwTHFLgEYLfa5bq1
/Nsmv3olOXfHy1UNpbLlop0L/BOSqF/wllcmI90k4JrICa/gJACkud6TQ/L5R1lJ
eoFjtWDKV+HJGjICZKMJJULkY/XteepbJb+qfElFrD0SNHSt0kkpT8zdxv2OpBBA
kTHYqv6DUUCfMbY4dqK32KaGhzH9PDqEmMTUG831bQt2AE3pCQFd68D4OH1zRRuc
aH+IE10Bw29RV9VwjQOaFh08NxLDlM4xRS8Ag+V7+1Si0e7FEy6638iWeUyJscRM
zLqHANFgn7yf68egTacHGjfytI6qT1oYid/3oyGGWM4aJuGoHD943x/Tn2noBkWs
U2jY7tF/R2pWMiuWfnGNw2Nk7TEHYlfIi8bTWLv0RpxoJ6dVy1BkQ7ompltjoEuT
C+sz8YzG93SOTnuqmLFFm+V8jXdO/D4iujMs2XO+YVARHJFQEzBPUbBDiWmiBjSK
VZbFZOkYb72YNupSiSGE5f/HDDZu9jD3N4EBqfB2O3s28xwyB99+D86+b+g4dY5E
c3D1vmMvBJEmXp+0I6QkRrMxDkH4PICzHtFuQmRNYhob5Bd6G9vNI0DD3dLwbgYn
uUp7D0XagVeWabLUasgD2f7hPHUh8qfhwf7mJFziUWhZxyPPvcr+5hmTyFfyX1Gq
h5RO0mMni3wmZ4NHTV4N1FWGI8x3AokrmsSDM1GwyRycxsfkTCENsEW3jSJG76a2
7MpwtS7eKuOEUt7qZwfFDsz2nWU3MoCB9cq+l/GmX5NJm0PFNqCVj6rWIAl4g8sL
W2KiLNEUa34AomGIFVeK6pj16ktC0Muojf9EZYGy9h8qckfPW+2/89ljFe/FhEg4
eL7qSVBSeymQze9YzcsWgkmtLwJEAUTXsVLT9Npgm75OtGtUw9tuextydRD8/YCS
gn2sluUYrUx+tbCZ7zb3I2N7Lm24IVkr7U1hhCsfh7VfyHVIjbDacbr2FvV54SrR
8AUtYIow8K526qyNwypC2/OBLIXCwAktLaZlJbu+LH3Y4aDe2+Hxgkd8YmEK7fNA
IelSUhxizAp5l0GHyhktB40eA5VWLb/somDkFeJTi9frARnDnv/MiDPtJBzxSmJO
wxnyEwJsETFOCQiruhiNaWiE9P2UDbYziCAaH7XZ8Ru+642xgm0AYp8Jbv9vFzdz
PU/VAq5hZTrjOPU6URtldmvu/GBVHSGRqAtdvAlGK1KEt0KIpLaXbg67/DNIG3GS
VS+mmnvtLHxA94QZu+HpvDjr0tPz+Fz6mLWL68ZU51dRbKGmJo0soe8Pv7fMMmVG
xuraPWOpXY7ZZLUNrHeFvMWG2SeurS1S25tHsDkqfHzeggkmPfz/Po0dkU501o51
t0dDOh3xSrenhfjkfM8j16E+tPTos0hwvXD5RpW8IKn72lNwztauoSinGS3+0LUh
bFiD1KS5dD84NhwP+DIKENHL/t/A7PijywGX26KvcgnOfLyy57dCkLIgj9EAEvYq
NiKqTQvChx72F5p9BY3I4CYveHzxBj4JCptWbLeDzh6jR5n1IBci4mpoAlqLI39U
Hb6SeLBI5mZ5pjrMf1lQ5X5jdVJ8RswvdaiGtqLqdLuPI3ED+PvhagarfNi080Fv
1h0Z1GXvMHSmBPNecjtkKVSQ72QWtxPcs1nLHbJmLkrOPHrb2Nn/sq1OdhO5kIII
xihUMiHI5bBZmyLGmv73A6G7HIp66aYu+DMcYXGSv+vgGf0wpAY0DBFXWun/W7w7
w4uVMuD28dgS6sdgNYvRlQ0kVf0osGNXfj+Rfn9clWqj8zBDhno5CJE2mjZ4EE9Z
gZ9nR+zil0hZoDhfM0j95Ref72zAIf3SAdo9shZrlR1CjVyFJlkpp6Ky45WZ4SXa
JQqPszMnzdOMsIGDY+cEQdt+ot61FNhMxM2TuY09LhKTL5uj3Rp5gsaU4dsNQ6tc
aH82VH/XAr1gWUQykvzeBuaSCk8ug0XS+3A7kFdzCH5e37D+RUdcvR3C+12mJF7+
ZeyToRp/4Wng/miyuhzPjKX0i5d/owIFjZVtiufULgEB9fdOutxfaOInF+L8AkIO
qWcMwAAdqFQpgFbgzhdU4o1mq0Qly8uIRnUVbCK9gTlgCyiuEStdku9qUz7Oa1IN
rTrFLzfabs5583FQ6MlgvdRaHdhjUvTfjig7h2NBe9Hbj3DF0O9pbPI7okb85x5T
WBekZ38yiC4ua64ISZiAsOuN3U5u/MQhAhywgfPciZ8wPGUgI9nO/YR2f5+fmF1h
IVoRs47w0zlmWwUWoRBx0KJUDUppkZIizleYDvhi3ykYOibl01mL/YQFOr01twIw
9oYY2RXevaRMec8qtFdX8HfX7Ra0UVkrj/bamppxO6Atyz8hgHUorQutbeAr6awk
abjZHIC/O3Uha2yYK8HvnnxQBcOnG4s4KqjzsTPsaO0UOq0B17q6CXj4ntlpzndH
dZCTUj5vdN5fFJlmyQ2+XnQyluMQXXq8gptagsKlVRo1na1wHFDhkcdhBFwN6BC2
meVKeQuHuzPZoZg2k/Ay0rpMKXgp0lomJoTqyfAORB+im7S2RXleATqfqc2J4rLn
budJFgtS/95FQG15xS3gZQQCmj13NtwUGP7I5IjtS4/cUSB7KfcdlavjD/tY8D8W
Rl5QHIi8gMl2RtEAfAuFA/kWRrwCjMWbayhe7MzW020mKn48G1i70+O9woaVZf4M
39KhPIPFdjXMaRKVc1T/t1cTGmIaYs7arEfxiPszzUwh1MRL+6aRk+A+1ClZq1I+
tQNQUMgc/kP5UajerYJN8el2tfvib4FA0tYXrv9bJk/02S0tEHZOkxUyZFTqm7BF
T/yBmySYp3eks9aHk0D4rd4wJIiOqCW7ifJuNg6HYBb+QuzDC0dgZZSVB2m8vpxG
qve1xcnZmYlsPC/lnY24jmgl+B+O+x808ERMRhfqmhEPRmmSwt2wxQnM2d/uUaqM
A7d15uLgupWDjjeVLcSjEXarg/UkaNgFtWZJa1rCJhgb4DsuylU5cjCjmR91/gvY
8gL6J5zDOB7m8P0pTWmktVisDY2GM0RXfCLFueLPTa3Wl2ycc9e7AivlGqTyFjrG
QGoX9KCkAQSJjPTDBU8+p+rxXgMCAOQ7+w7yc+go8qElPEbrVv4R7AhsYtHs6p0I
iLTGi1wGXwi6FoRNWF8gsCTcc5osXruQ3k1Kn6/RegdJxyReGRRaSijwo8xJ19VU
TkPrVmT/eKKinaKpHRcR8mWoj1Q8Dp+AWZvtc8Xx8NU6t8NE3dSCct8ePLvOcSaV
REIrUQhDxlOEwVYt/pBXjJWU8Ul1/0lwjtINk7zmr53VRZOY4woavEZzqp9+3rOQ
QpFw3gPyH1t7RY82nVGiL0qtSionm3QOMC9tHm6pf7hQUOh6YkcU/CSkkKJeWRFx
M1Xzapjwl+yUpFUDlGFtjCRDuFXt/LWectZqDFP81Qj+FePc3d7zR2coj/DyMRiX
tVe6dqjJJjkyOUYnswsSSw4KL5ydAqTbT15iGOZkWGvwDjGNYBJSldPRQ5zwd0qs
P0lAYfasG37869gVojOGHDPLe77sj/GztM9LVWs6lrDIgg5VKU8SP05fDei2TrOd
IYI/7fDw/bD6l0/NK7wZrDy1xQjoVjoTJROyeIUpY1W4mqTbcdF7wVr+VkdlijEW
p30xeh3UOMDypXYbjg7bIUcIGpBM4OtdxdQ5BUZqx5hzwJ8wEUQeJW/ruJl5q5Sr
YObXUoPjUKvPuI7KsmIN94+hlTFpleh2d3ZISfjzbNJ7z1AVoSyKEzIF8jQynetO
759UxBtIA8g5QUnTYDqVQB+6GFYA8eNcUYHtFsMsb5ktLFpbCV7s/DL00Rb7D7Ic
t8ixWFu0Ejh64RzIjtjw/bK1VtaEEBPK7YGHjs2TtWh4de4MvjxebVMVW5IimOwZ
C/ydy37vJCXgN2kUkDMGGq9HCFlZJVUhNLmdrUZl09ys5toaViTVXDBquFo+OAFY
1cEGLTYzuBHjnicVNM3hc7ePFtGeA8cHuavtJIqSNRUQrjF2drJSp/9qs+XNPyEC
O4JdQLTmTDm3t6sKYEpWtgFtTqx/1y979ySN8IkjlVpgF0a5dORoprx+C0y6WgxR
foKwkJ14mn4SzM4+GKjKtiX0c8HYknI5YI7GF/eyDBssEkpDUwEsq5PVmJIL/fG4
yTSS/KmJrujnMpZoFiY8TMJFkyo+FIbRUolggkvuIj6uWNXkwlUh4PCOOU6nRDm8
TqHzZnjTeGMpR4ZINoJExI4iVEj11QoIEBiFa6wGxhnmT2UkygK58xOzmk1QLugF
QhQ8v/aOAT8LMf5OJFaw7IjrM/Kv3eIsDq8zLKGDnDPEzPrnukyI8MpLMA5qObNO
nC/cKeP8FpuU6tsVPtFfdKlZPI125wx5stIuoASun72GpVA2vWQzE0vUM2whtanV
O7Q4jbWG1ZFwQwnHOm7lSMKXhmyHgOm8x11CfcbmmjYiSSow7tX+UhuaqezOXgDf
gftYvaMRSiacQmAVbPy4yDR/yuXsUK4Rx4OOO7qLBjQftX/WNP+dazIvPsCwLp1G
vaaoNSvJgR/bYrU2RYkAP89rftJUQC5sYUwRm5PEEZBxjXUCvpd1I8Ih1R0JNkDf
Ui3MUUKWez7SZ0IFWE3neCMjBuwb4GZnwR0NuDZ+5sg66ul6i/iGezXbydWLa3rO
T2BS0INvtnlNSC/thVtaGVzxT4I4IE2VHvOuzx5YnTnTcDCs49PKiWYhJg/5ymKf
2ORSGyaMiEXwSFJT60/B2w93XbnqwJO9Dx85n5/75rvRdpu9V4CpWTpgvxhzdnTt
qJgA4b8HCx6Y2U4imsRdI3vukzLzq/ftyCOYu/8sP7TlRllHAgYgXaVvjgLNozJV
A3e6ouJiz9p8oHY9VJYOCpZ+b/x/Hvq3+ucH5nr57O/44pEfx/BrF/LTIDQAU+Ib
/G4GREf7NetKfcaKhvZhRCnRZhzveAHhrdN43y4LTI+N/pwiooRXIxxGSmK44FIC
6tOHWIjPP7AWNQJ8/nlwvHYeUO2JD4B7VXp8LBXnJ56xtAdH2/01Vik20+R8S5R6
xSD7Lh1MLg6l8UIfxdXu/SAviLuiXZmqVrAlkj9nMW5VeMzlnDkaGoC6Ng8pVr14
a8wpkbO3zCyYbQ/Vnq4lW6eOJKQuCOEhNd5yLGbylY049l2j/aoJNgTXaimDhsdE
7ib8MA+BPFGDOUaVQrw7W0EDrgxa6yLo0+JqDZQ+xx8z6teaqqSPphbP8FKS/nqc
2TdRJzJZaFcvVbH9He/+7d9O2Yb9uH8Ko4zIvO171DDRLWtju4W/cVt29oCHQlxA
YesJe37i/lmCuzm6SAsCTIY5vcEW2DYimYjo++b5TVtMwfGly2eU9lQwQALhS35d
pM+9Bw4riAN1MKOAoeRodWS6Qv1RxChDhuC06KIYWcOL47duAJqkx4kqLC2aWNkF
u4FmLCALO54AiSQSIub6jK7i/EhIejqSWeO7+dYRrgLiaZCo4NaO9pXGc8v865OJ
KxzQDlLUK7/fwrG8B37qiH9yvNxqsL06wf8/UXfGzkSLxhoBofbNk+h2EriQiW+7
X4LqCCvP2606+sYq51/bDDMvxvEH0JyhYf9n1vleZtbSCHRHt8JAZ/h9xFn4agyT
k2g/iamrAHN2x4DnHK8RVmKjhkfdRrShmbCUX7HfZr/XGSk1Cujfw3zHNjEmjuWr
FaOemFIDZKZ8+gOQSNRe1EGIrmmdEn2U3A80o8hPjZVZz07qQnokMe8XhtNZ7oxF
97+n8VdkSiELmtg8waSa0tuKJirlbEAr4dIkNeKVysAxRjhG7XfVo3CLJiKdIdxb
M7UQbp3OwqLSxK0caJ1ugtuiKAwLfsMv17u6nhARbMajRlkkD1IgPeurlyVVv4HA
DwCdtBrKUtUaraNj8tdAFRCtXXonH8sss+2hiGdR3xBu/ZuCxyWYb1BXu3ej4yXo
2gYM4enth841k0hg7iVx/1NsYwmIRO4F1VpFpJLbdZ5RBDvhsVBryCNr8o0KCW8N
ZR4Tm/fLKfdzB7udQYhHlz8P3QLlDxVz5R6VYV//Z+mpluIqyVoNqbOBbmrPrvbj
+bvsFAFAQME5BWPiPurM7ijxzucS9LErKsxKLDPOz85f+jsfxZbXJ4bZlbmwqi9y
neOc4mqjHZU+sOyW+WGCBaz1IBXSetPTmUBNZJRMxTdk22A1WUMgqIiQhRz2ZTR4
wPJUNGxYMv7pZNOSF5670kAS1mY0DkLf6dDKTqP1mx8T79X6VFLLH2G+vmzXASRr
cpuVcDl/8kDzoocIsFdnSCcU1zMlQzbiMm9dc/oVAJfs8WS17oYTXG6E7PKI6HK+
R6heb5pq2W1qdIn5cpqG4D0ulaaccbA0VZyHqmW+uqtenGgJ19XowqzTZFLoRRH6
5ysOEI/h62d9Bg58hvU9xaLipD9llz5kDjzeDjZ1Z7goV8LEQvT/zCK9KoCnT66j
crP5+deHBWhyxZAX3/nUmnyFnIZ3EUivzahYNZ8x7S3Ma5+QKrriFKay2tQC9OE0
H7DtlPHEQdha1pkB5rB/jdqGZE5TXCabg5qyF3u+jInTX1T6nJ5ylNaEPjtCaQED
SCfA3fJfPIKhQkhC+owzHs9vl1gT1ZJBa1aWKHV6gVEhp0m64x1eXuAWEMtITHsg
9kp+ADlQxFJXLZsD7xPcoW45jh6xGDiadwv2+LMAoylqvNqKgXV0jHatQk+3Txkh
0IXsQAmg6ZtE1C6a9JOgOv7Zh+/WakTAOBYQzgtYVCBFNvbczbaAmc42mFKc7tHM
GrHZYwPJValvOw2SIWc2BAc8H8BFhvEH88viowmYAzaItBNf4UMb3Q31xzLt6OVz
AHOHKwu+zemtIMxyb7DwdZubvnOHl4Ii08+fha1K27JbDftN8apXY3nXR2obY6sJ
2QmE2nMyGQZ9Wj0X91eGnLMLnYJ6pZRERpxbCgtDNZ4leylaeAne+hIBtnC6rVjS
QE0v8Ngd+s/V3uuds7aJCidx1f/2Ne4UifilHY7TIRSnsLVw1wLuyHrUpFDlo706
dUExI6ms7exDWIIwXtF51aGmjOt1+Cd/kw1H3vTBLqgiDxIrZrOfpFjqn/XkLyqi
0LUqp8AvQt44M/xB1v3NVTa2xA4V7dVgQTGIfJTlSU56bMjzAjyfx60o90yZW4R0
DHTkPAWJHMwAZDG4Q/qamjtOsL41nt672iTFgEt7bw3Ae2VWLb4ainCAcq5teTy5
6QMjRDs8L/m7O2BpMaeTCGSlnSK1G+/y0vKGpfAdRgLQ5VfJ/3hsSXPwwg3sMjfa
n2AIbT6KQ2CQu1SK2bj0fYfOAxlr9Ruxxmir39JxUKqZBYaJCj+BOoM14X0YePGo
UuDhI2CPGPdUbB5G/c5vQm/efbfaw5fr2VhLraJYQeT5UQfFuRevbck6MM4qJ+q/
JOWnvE9svqsSDInB3bNRY5ksOljOq6mFKFmZPWBp/JQmGdRIOpEni0xBKDpQyf+g
cNmD/eUhKXq7gWMPyJrOuUOkSJ+C7YKE9ValwDU6KgXjv1IgjDTB7MeXtVFZ950T
mjbtojPzF0vBHwww0fWSf+ADFsURiK+yrpc7K65v8h2Wu1krptu+SokuxirJdDer
vWMTnKhIRTORld0rw430RiH+y4BI5UT7uf+87pCff15OvYdF0CcYIt77BuH0C3hq
vHYG4+xAA5EKnKYX6m+fEPYX8Nfj48KKN7k1/Vv9B+SqAGh5nZGzXAUNF9DCM72G
dmTPkzT8BojzrcOdFA8AdCxMzKL+1Jk+q6t23XN2erbx0HTKss8C4mB8c5+xFz8J
MVzSgs3bCkzeKXRCXjIub61UTggykgwln+FIB1NU6JLh+LdHkRVNJEd5J6Hm7Fs4
DxBfM0ItfoY5QHZ9jz7PpKf+76skWVAleZmFbl38jfUYicCT8hALd06icLWyiAGY
n0OQGPDtqdQAOJ9b8y4bp6eo+PZ+A5ssNeV/HMSQopU3YCQ8KuFyyTBtJhaoiQOZ
DfJctJ+bWJeFUYGVpwTX5yGYH1m4uLL4wjk9mIhTX36yMA6SEKE13vcgPTd6A+uJ
h6MfK0e7oxjVwVx+ijlY7/skcrtAD2qRIBbqKIj/QpIKBk6/uqBQPP6NCv0TiEba
W0mseGA6Q5s3Lc7JxsbceQ3mldNy3q3yMRMlwh6IFMRl3fmzH2T/KMqGUlw0zFCU
chbddnNAtcXwV3FuK0P++zvxI697sYITC9a/CyvG0UA84RqdTkMbLJBRZrHOJjZR
Ktu6UXfiTUUFDzrPCBHXSs5PZBOM2cm0bwEAex0o/+XGzccvUNht4aljUWcbE8I8
wHoC1caNZp5x18SAgJdtVxSB+vJv6Ru6HDxUzj9SWiBRt7QiBsgcnaL4guCKYDCi
PV4r3DqUpEly0Si9DcCEYrVQDVp5pdphhgxAGmdBD564ExN3wl6TpA+AWAf0mvUv
1Au3ygyqPIcPlwiCDcQHqs11196Qsb0ZVnFOP3UipZ2ICzc0bORgX1IGTasHovfs
szhOs1OHvSicu34fUvKmnF1JQMesq8+rCyAfRbGLFqMEn3WpniyuBweP6LNOJ2MI
8sJaX/GR+KvsYerip7yKSGYwUPPoVDs43VwiQS0+lJyzOs1BvQYZEYlZeXWK+/cS
K3KQb5suBDZf7eE+6xZ9g3sq/LB5X57WVXlC+7spbTbbl6q/Vgkv1JilFH+585Nh
5hsl9AcPP2wd3pBI5tJl9qK9bhO8JQcEROiMj2tkH84OTXak7thI9BdVTAURYpBO
XATFaSk7AuwWEuqC0h+oXTvNNgSq/5GkWWemLZToBH3jz/7V6M2namWmvnRWqVUK
mTS1g7nQ8nkD9X8MVrtjtbnREjN3hX38hMI8HnzM6lci73iPkErJllaldksV94wO
ksGxTsY0e554PCVNmHLG5RxN0uL2eTGSojXeslTCiDrWUriGWqVC8JG8CoukljcP
Txe7oIiiZeeq4Ua1RGWl+ploIWNxp3vQOG4AwIqdnXnmgZj2uItXlEkQM7Ao6dPu
zvx25ABSQ2ScVYWKy4eZ+CsmojWbItlfCMboEkcLLpNeyBbZKFvQ1wupS/t78fEi
j9ROarGXlWFkRa8iSN/5es7qq9zsKdUi1EQ98LxpdSWTEbWY6unhM7XQjh7C4UNt
Mn4dGUHF0OIvLAMsW5gb3PvjhbSyx5Dc6gauNZPK81XMRo3jzwk35rs9MnYlweoV
7R+LcmjpKxxkGIMovR+MljH2LLznqyVabAxFzDMhmCnsRUjwxSuE9s7LByG5jRQg
Qc0Jpibo61qjjf/pKAQxJicmZKwMEcp5sb8N0B6hLG+3Jy0m6qhEP8+4f1nvrIUg
CRo72WXde4CAXDH9ns4ecALX0P8n0e+Vb85O41zjMBbdy2qRxmRFkDlKy4/5pge1
J35Zu545+9Qkjol8UENwroRNWWe2K8ZB3sbXxgrVuqi2HD8yRsRzaThMbH9G7oNZ
qvJ2oDVP6KISGbJo2/36xROz9T9VCs61o1dobtUHclDmHbR9iPnkuk/WWNc9JJsA
yoQHBbNex3FKWxHKIS5ARt5grk6dMX+bqsQkCRE4kqG10rE63R1bqzGQ+BWRMPHI
NtwbDqgD5pCIpozJb4ERsvo3h6hjSgxoVKJuRBn+0ezy2a/lzEKRmWFt8xcb/KDQ
MKXme0N+z2Nyae6qZhq6ejmX9DghpdIAVZel4hH01rBq5TGcD90p4p0bfI1Ak6/n
eOppaEOTV4w5skUAtC8SXg1dkgp4YRnnG8AfG9GQgTSLHjfvDIUQm5fzmuTf/BD6
077TGiHSXvIqnOJ1oTfL8zMkNRbhZfj1/IwP169egcy+VMzlZxawU8fzJmaM+u4n
4Qod8J/bOyJ5u8upzgCEu8isxDcYAZaXc51jRC+iyqAUOIOJcJRN7gASHhDOZBu0
FWEty0aNQnp/V1dutYzjl/1HPuFa47pqdEaJA1unZiyFrkng6Jxg/I9zxP+9U+dH
RWBJVwrz2N1Ci0ZlO9qtO1Z0iE1TNbwivq1s3mCv7RzcGFnwMl/70LDwxZYx2anH
IEDwycZh/WLwhrd8xa9gYG9zfB1LEoIW6O3suCycGyIY56XzD1kPJshP6jl8/HTC
kuA1KnIZI8SrUnSMJgTzqeLZqHfk6oC5TlZarVH2VXCeCRPc6+U0Iv3QuezGAAuK
LsG87TnWuaUpeJfVfcJ7ey8aqMwYVX4nZSJSo58DIpN8koUebzJT35EC04rYKSTZ
5nqwao4uL/+CJfgQC9ITJP/rULPb1DCnm0ci3cnnmdb3hdZTHEoJDeizRmz2TwMK
saWMyRK1fmdl7d6NrFuXiy452ETywAUdKpOeoaIRH9XkAVVdoiGQtI5eBbNjslhm
fZlrhJbzeAYoYAFjl7qbEM2UcmWMWC2GnZWqvJjKG24646VswUh2PLhGdRTldcK8
0ETWzZJDm7FQHBKEUkBzf8EiTmTYzlKofVvukmrWCcOD/joRPluW+KerWAftPePn
mzMiuhaPvPVWqtrNzpe/cU42PMD21ympkNTu20hIYvm89D5QgaU9MoTvGeuIBEJu
neovm7jU1UfQk9LtNeF2hDXXocAdv38eUA7boi159QwIDjWFDn2HC3wDhL5K119D
8Y/sEuT/hCN1A95u6NBQ8f1FLzg/6p0EIX9vO5IuLC0iaygLaLMFjHdUI5jw1X3L
0H6nhZ3dFVhRvxRntoT4uBFaOhwXWc3yZLXXiwW9Xp0YIfUdIv0WsgmJ8Vdf1/6f
rfuIZz5RwYJ+nw08C+4COkYj+W8G9vwCGEMDTXVkVw4isbcRKX0uoDeK7hDu1d+C
HKfUTiZBeqxSdy899xtbaufS/4LpjrRs7Hu3/Zhhv8lK3Z/R40YdXOjFDlD04x4Y
6VNJ6bXMNwRq0v8U8Bzva99J0dA7dqrjRRYIQOidgtyiMRLVq1fc3g7Kgv//uRqw
KRkEfD8AiqxiaAJPm9LpB232sswLEVpTVw1L6Op0T0kJ5fI3wvAi5iWMWqceRlVz
5A9EJTdsFMIoFd/t7DEmHhfm24KsEdIx/Zz9B7JDgFYsJrf6mghzwb+cR6Y9POej
pvf1sBmNm+QgccbOYlNQSnh+WSVvd3s0kuis7ZDBsVuc31TRKz9zd3BomwLGJ4AR
d7CSbezBepA9mEB5VGHboEkLy/PT/6bujaKhTZZ2b5nhkVdE5p0FuVI+Kuj7fLxa
GSDnZRhgLLiciTA73WKuMiUNqsj3WrsxBCnJYemiZqk/VERVkS6Dq+w7hciHVpK8
GbCvatkCWbcYRnv0V9TpvFGvHcAY6SXLBEenzYtwVDC9zPA7qwT6YvI/SdQNNFfd
NxB2NWzyKnSOc8pzZXtDBjHY3AN63NMIDYGuqQZ1IfjyIziqg+HeLaKdTV8/Dzau
mOCl7gKBuZ0gXEffY6dZ0fb6RmJUHNgeDfoQ4irsTOiXpjsfIrp8hE6axr4BFz3n
W9ZOg8HICp4GDRxKZm+OEIRmg4BO+1HdP8ur47H+LNt98+qPXC4wBBDrNCB5mmQy
KKHcgprCP71yHdKcv+h20wnSUzo6VzYZoICQ6XEewRClMMAKWXZbFHQXkwkvcplT
AKksyfNhE7kmtwcfc/H2bLbPm/9jRkirfcY5JvQEXyiGT5yvjl8fdbxNGRHcLQxJ
YgrTvCSJfv4SNGSr7GJxjovM3iZ40bLGU9MkgliWOSN57L9aKTDHArJrqZn/Sbj1
m7NQEy/7eIpacaWEr6h+lnzFQB3Yyura/W1JWoODuX5UBBH9BB9boIAsOBMv3CcG
A558vwgGWQYX7A7cgb5y9jhGRj8iW6OKuP49SzXQ90o0F0ynT4BQqQDtBO3DnorJ
wLBPC+H2Ev0AgxWbDJ87A5xBOwNXPa9tUDWmxc+oQArokhpqGuNP3SxsdaKwFPbl
7avrku7QKizwqRUjCfKNNixWu+IyFIrqXMEqpJlTtf6wPNj8GY2h9NsysS/kaEr4
KHUwaOmoTjFVJtQgiHFJy87mBOK00Y3T3pyjjmgPlnYhO6W2wuj2swZcS3dxMDO3
jhf/lGEkGu4dm61QtCSeAA4LRuXmBFfunjD3Z62pQ1Nf9eQ9iW2rW42K+dmoQRJr
JfjSd+bfP+a6ZOOGwetjQbQo9P9ZNTbad2smTtyCLVqZ2pHsAbGBR5RPOQwx/23z
b9Umk0F8nCjGQoASV4xTyDLdUrJBZMx/Kt+JnCekZBb+UpfW1zv0HInJGLjOUoFS
TxJmiXcsubOeniPWRoS6W05JuD6reLYUlkIGKcLu8ZKCl7MfO31vDRH5w95+ka9c
25bHlX8yv7dgtCBOalV8q8N2BzfzEL8rr3MNMc7jPActFroMr9xINg6Ocy0PCygA
EopASPFBqK4QQeg8kq0LGNR8ogwmItERJn1Hq7z6dJfM3kYCcI5VditbixsA4xjf
/UsA4KINpJh8Edfi4XQspfLn4UzwwJRwz4UthLB77EQpoC1xNA85JXrxSvoDFa9q
qMvkBQdWK0pdVWO4DraG04MRQLcR9gahsfgEqrd2xhIaR2dgEbv3gR44a02JJJ8a
3zpFkgfexL3OskW1143rg7RDH+2CW1ii/ZswEhuWEJ75v7hGSIC/iM5rijLaT3Kq
QCdICQFEsDFh90f8CHmj0Pyd3P+NUu8FOQ0gbU4e2uye94VMQ4oERgKsNLQaHLAz
vknXeKgCj6c3BG9CWCkGwMcAKXRL7ePa/8gVezOub3HNB8klyfOl974+ZLZjSOW2
CQJtiY+fBJl/bcK9SZd8T6q5VGvGppaWHJdWdgnhd62AFPeIDmAcZX09mNEim7pQ
5DGMQG8stWIeCv1enJtYgNxzAYSHbyqYo+qMuzjkhyHzWMn10iC8V6WbfaK17+0E
A1lkkIEry8TWOC9sOOGDhLfTRSjRoJP7tJOoWLz00YscowDPAkjwQpNGCkwVwbUK
fTkBj468AAY2sN9JnArxlyGHdO5n14FmS/UkNS7y+x92oCmCgT3PlEcMpbd5Azam
qWPzMHlahfD41pxOe6E4dUDXe4OeyftQzAZSqJWeJmYbsT7cKilzEre4TkmNMaX5
6AeiZus3L1F2C885UcWswfz7s5MEqESBY1NY4BIV3LR3/ooH4HnRTPfwhBM2rOA1
Du/SbsMHWK9eRUlGoHKr6JlcRzJ80vMWZLTxHm9I4o3PFNnxaA0lvmCDnldBWTt+
3wWuU2pbnTGSUdIe0dHN3U+w9TykHbuR4VqMtSIrelv2YmvO6IEajj6O/jWZoPOg
2Fgyfn9DdFoU7JNO/Oyw98eDbNnKAofexeTYk8rrQcug+W8xfIfvoju2+oefyz/3
DVv3fkXvvR0CnZc1ur2cb9/WgQSFpkOduAdc1ldHVO33qkKz+VNAZmcsczkvWeZE
epVZavtq7OY4UZ7a3y2x0s/6W3/UPlASbpfOC7OmyGFjEjDM+SyOIClN5cSttVQA
guapqNqAYF2Gl4nQi/1LZZbkQlUX8zl6FZ9/TWCouKWZ3zeGqG2b+7d3McSdTDyy
qSFwET9Br28J99iVPmOxgnl7YhuX5LOM5WO1nUJ53owiL89Hqd2m7UReytq1W0Mm
ZTadb/2e2To9xA7n83Youm0evz3cFAIVTiwyJiqyPBm9BvZMME3HpG52dljHtoH6
UUe3EU+90FFgmNHjebBgwU/yVTaV/WAziXCyApo5jx9ZqsVCiAN0EOoIILdQomuu
uzYS6sA9nDnwaKZY7HrjcqS7Fq03cOcoK5FW8kZlhHpfSaj4vuUOy5Vf8jT9Ka3t
C5Ian6RrvdQfzkf3HbxrnD9Okdpaynri7S+L6apLow3VWzwQNqzspIYoh6yaEo+/
m/DyiWD1Sv3iG+outH30+PSfcqHzhv5fBDMgeEoVl2HqJVPNdg6hxaaZBYCAhpKU
jHN1tpluc1i3T3b4cmj1t0IEmKnIds787e2Xea68dtpYGA8rkIUjPHC8RbFB1PUi
Yj9QpGx68w0eyfmbxMx5OFu9ACUqVi3MGwGbp9nPh78vm/Y2v3m+J4guHWiGIj0W
jMCI1BU4ptQ9ek87jGGDBoTvJM/e1pbuRar8A0uLwZGcC0u5l8hxMlnQuX/ZQTQ1
FZDIVjOdycO7nPpiIXRwt1J6FS4xho93ulByTqU9AnjnsFvBQVyUoOmTVTX9LbDS
XkPdM1NaPHoxebIt0Wt3yTZIU/Ic3CLwS7Z8ytEecJlmyMiRkaKUQJ89uSHhe0sp
6rPiZq4fkPoZsD15o+gUQusMNN0DK7lKf6WzRiFQPagL6j524TP1TGwaaT/JeQTR
dMetT3y4MF4Y6GrP+dBmsVFbLYue2rOsCOXrs9Aj6v14gHtS9jkwBKqCQchVvq5v
2Mp9vvmHO5e3EwluQTReSiNtJM3oaKPUNn7Mdi233+rV0fw6f/gJEbwWEBW4hKYF
N15MWKuLpZRo3a+XroDIt4a1KEDnIJZej/tOFDHwhEgBqhH3jQztN5H61dZYWRTL
jUiLPg0wrKdHF7FrUMeucrr017OO0x1PqOSDRmvoNRG2gghcKpFqRQzwdAIUGPrL
j7Ck7Qlsb/eBAJQW7pASadH0dcTFI103Lq8SwNWepgvuxrOFA7TpBf4vgHA6Hpkx
eetRjw6wCyz18Wg0xdvuKp79Lus4MOtlNWDCpmXBG/TjFvspw9YlNFN1uKbvR94h
btqZf/BrZARuQaLQKQ0u9uLpGCv+bCbsq0WBr/v09vIW3VKdFaF0ONzNGtn/evho
nmtApDiJXUaV6oPB2Wm49/3JSXqLHl7qQE4hBs+ymPPVPFlJ1tazmj1NH1LxKEv/
yuZsbSe/I5GZqdkUX9Uoo7r7IYsakj00Ix+GWyphgHZOv7wCOEX0jsCd1PYWicRt
4nV+Ac2UCb8duL9/KBXy+U8MSZEOAJCz0E80s0y+k8nE3t4dY86zkaCdrX+8GrJa
lmXSCeK9MeyywSImRUuTT0qduTIodTrBTPP43L3aUEgl7Fpm9IxWXBY5Z0urf8c3
EQeJcThuIvfX6tt2CMhobxda9oDhCR54ZHvJ99coPpVTnjsHO4RSEa/YAZo/Zjfn
anGeduMXpXVKqEdtrBZ3s44EhmDlRn3Dkk0dinrl/k7CVzZJQrnfULfPdbQ10d3y
6qpjy8PveDrlYotfi9778kdqFd887iy/ollK+Xn+bW6efDi0FoCrX7t93PCzi0Ce
MUnhh+WIxCJBnY2/0jykLYxDGo4VWH9RaEx2JhYXerMIGqiv68mY9L+5oqBII9aZ
GmtgbPbc3k/rESrPZvwWmTuh+XylF/Lr3ys7TKGNlW/Uea1Ea/F1RyXzLjtfVrKS
FCTveP9uKB/U1N+CF/XLwpg8wRqcYMDTPBeB5gdGIdmLNj/YKaLBYLD1BdrSNfLQ
fp44Ee5yerinH5GwB1oobjykrHPy1Sl4nN6QaznkIecSl+htNSLK1y8t262YoIGi
+P1GpUbGJR+tTXl3aJLkExCNkQtU2zkbjOkWLRlVvpgZkYCocNzmcHZPReWbYO32
zwcj078gTfEp2w0ZvhI68c0S43MuJwetALmFqTZZG34YyBEmfGripa36lSEUtA71
eFhVNuBpqfLKMsR5ixxHYdTnnJGX5cRGU7+r5pCaZie7PtYA33VVgoVphQxxjzl3
lwoSnrcqKIFVUwoxbxf3LjGnnB15SmwT0bkWzDEAG6uf9B870BM8qkUSq7j80Tdb
lENL33PlJaF0DosRZg8aeVhzdRxHWv3j3IKYL2NPIE+ajEKsX9L2sb60r8ighloX
gp2bMf7sNGkZwTuJPxKkGeAtO2jcC8IXSuIcE9G0So6f3yU8imwZarEoD5UTWD5/
/Pwfbxc9eVGj73tNxN0dOTSQwXgZ/fhQ/W4Hj2+YLaZ0nITsOIOmDQjXfFizgwu3
+mZrWxHsDdBPU9LqCO5qih8CCrRCa/q7oXmOLToxFNRR5Vq6OlH2/JewpVgvZllN
4HyA4abskO1hN5akP1DGZjj6LS53iUZvrQGhWlgsqluqTB8CygseDPJI/d+8WyrO
NRbbZM1zQGOl9cyL5fa8075kKc5CGjnJiiK3hmqrKsdeLFmCHDGk20Qqsb27M/Tf
r2IcaNpfYbfeguoRS8PvwZJX2ENDdi2xuLRFu25DSmz7CfQ35UuuBzcP3ocJTKow
a2h9UjNAiCshQGcdme4z8mmAinISTC7seAfjJjXd54ClPVPBL84nOP28L6M8hKT6
p+QALMlOc8FDaWyA7R/DCdRGZG/Qkwor1LiWBggRYfzxKuVjzYB71/1OjiuofPS4
k0gRNpS5aIo2XWpbcEYUOzKa0J0De4trIhn4Kkz2dSvTMcqCFL9eQ+3VZvsS7lln
ESq0PWtLYZpcyrfWr2GawzNKpXWDCQ5Qzi3EhytT3Xj6vkvx3o7AjIVbPdsweQx6
ywbvFAiB8KKg74I1GkSSZ5vET/B2CD4d8Vdkw9XCQgMWqkFN60DVhPu54w2AoexG
OG8u7e5tgAj12lf4x9ZxUAzDuoHfVhTXEF2atnrBJqsU2INpAQekiojPqFuVmhQy
just1a1Di40ZjXICB7ASYGhDUP15eU0Lxy4NA+1FyGsW9XgxlhuWsK8e2Je1UWwq
RgvNdQ6S22o5enwjUjKXkJ+0Ef2I2NNEzfeSueqlrb7X30NOsnTNWejI+G5B516J
5HGYfrTFHxYpBRDpr3JiQFqwZGZlPHqam9bGhvm3RDWJyDb/h3QNnw+wP5bv182w
H3AqV7dxDo3w6HKxTagkh1B261RUpugtWQMBPagF62yw4eIW2dtZjOKePsBLdd0b
28aVHlLtgzTFiQRA6hVPj3fC2Qvc0eRMjqpjUYuxr4eLwV8LxyFxNRmYASnYbL/6
LpTozBJrLmOG2JhplLugfcC7iePwkSzHOfc1o3lqC0Tcqwx9hZGAp6gOLuS0h6mb
KgSs/tOFEWuuwjlqyLqr69dwKKXlgF+gakFWICr3HQn0tfGISn67B+8/+AIBlSBs
kO3ofqeiyCxLNKQO8kA+JpMsmbjIpQYKss6yjhhKzaaHz2PQlM4OnJzI5Wqh02Bw
P7Ml5xfQ6dAnTEJOIeZJsBPMF3zAYsi3ezzTmwWTADwGfC/gY0MDJAr3JHehpRSE
e6DhZCPTU+IneCf7+zqYDA1JECF0x28QhEHMy1uiK4n9eWoLgfWaFIHe51tw9IT3
F6r2ZTkVkVjqjGWW7kjjj2A6x2iGgN7I7jZ8xnYqMkkcnmqY6Q1+BBNPQ3cLIpT5
H4CS5CB16lSAkK7PCmurscwjLVUo1gE8Y8H9uTBp0saEVTGOtPiEykV0ghIu53PB
zIfoBhnZCB/YWAe0SSclf2D4ndWLsvn9ROtzQhfjcDUJu2v9GpL+ZQ6xJo4VZ1ZB
ciuZ41wANPoZKSdUU1VKSkJD3BQYKnc3shzLB5FmX8birs4JzDW2aFX+JKz1L7Rc
M4Vylm0rupye6PPqRKCjXo4OzQA4uJ1jt3bqta/RpMrLEaipuLKVCrsKZOyaiID5
K7Kj8hL3UJD2p+5/2DBf1kh5G3IOmi/e4UsQ0IQHvyfAJpsA1SYOTpjFUVM0gykf
YZKDNlf96YIMjf2sJd0Qz/y8fXA5JjmSHtcgMa+3ONyRDkoCY8s8/NcIb9SLaZRN
H7pzctwRIxfxf/DcgMrBQRSW+jFs+0rutVX84yzCG7fZpCcjV2gsmfamsAhcbNN9
riz1iK9xbNmCjlzYbhlMhdoIT+M6wcVLiSHHXXenIR1AAuxbToKe/mOXS1bBoxBR
KIxBF7Wy0Sf2w7fdja3RZqh4oRVCUfq/oUI5H4oHYseoHcZSb+PFQKg//meZ69rY
fJIWm2mRVZGB1vE0tOvjWfqXFnUiwIW61EBItduc0hBJUjYyOnjj0LLbikkwWTgc
vn6L1rdLl6/D+SIeb9nPta4yTIEigPJMfkyHZMHAPYaSH1TaQmz+0wsmtb+CBV3G
tWuE5PHb5EuhiPRPjZuusvY245aExue93g3Q3R7SpkVuTF/VssY06KN7wALYNS1m
UewJLwBztr2FlTlORZZHe1P6npdnYIzS23Iz0p4tcNJKk05iF72pyyrQd9qmSFnO
NdO/5Q6NUkDRQBqpXKQTBcRCWKkOIUjVnvQ2f5TYb9MiWmXw8KZJ1CfTXF1wkwef
lltkDGW6Qgkjzhg0maDISUdMXk8AQu7ebHeU50AUnI7S8BZvA97KLtfvWuPzYUgG
gjLXa8svURfGwKyYSulEoo/Ro5J5WA9SytyTULwggMUunHYO/lDEGi77Kx3RkcNF
kVql4VfY0J6R4eqtGhrn2Gp7BW5QgRZxLMrnboIuebkbb9RhHr2sVpwUhLpwJYwn
9bB9gdtJ/opUrspQexuNz6J6ktApnkml3efUkOt51EdQ1g5mEGv994IUlpa0HU3o
eEpSTTq/qB/QQj4sao4CDwHRVUdciIpC5mCak57M1CX4DEj6TIwoE0FQmwDYp/rk
k3wEr5l7q1wNH4iIYv86S4RF+wEvhIanet1oISqgTL29B+0rCDQqMoybTELYOmds
+ko0yjJ8U2NDaXz04Kg0sK93lP2bq9TE7cbbXAxifKyhd1hgwXomLdy1n8HlAE98
qp/vxMzdyOnr6zLclbBN3sc0BvVKgMdti7Zb1JvOCNhbTI/m0fmJf4CcHw520Wcr
YwQ861o/+jAuX3fds4t2IKuwtIq/ABdyKBeSocJX5AUEqiDaSk2SG4/Rx2KPmPgD
3/5rkbkjAgXH+Cju9TGMUHvwu7+C7RZGcbVu/MYOOwVT/+GUMzZpp6PDJNohbvYW
zsSdBCDbrZz8eBW6u9+BHadIePtxbaSkQ8RIXX9vRM85rA5xw6fAEh7zs4tybSv0
K0aDueRwyIoHmv1LjzLSE5Z8J4xvCjVfgX8RaBp3uDQ2QQ9Z/lDbWHBkEILAO0U9
ppBT4eFNJpohgY1hhfiPRcgXPOzkLiSc2ZWcAi4ciY/FADDsRQOO0jV5vOXW0sqH
YomupWN4MvmlyK2wFDvFHfuJCQOI+rkG1fLNM1/WuPU72EB/thdCtfcRhX6/Oljp
0sAGdDgHoBP0Uk6MIeo3iO0rzqEq7n1oFtaxP6HRgwCoi+ppu81jvyObHCBqMOcK
HFI6EPH6KgfdvcSBEKk9XryxwMZ/locP2yFDyat3HDm1mum9lUljw1PfI7CMnpOc
NFstif2JRAVwP8w8sQNVQ8zXMLMPIG7CoqJmeyksftBb12O4YeJSa9PzAb7LaNlz
RTal/4nwIasfHZc9sRVIyUCpT6VPzC7RK7FwmCBk2+l+wVQ1KVRN0mvzo2Q4jXAS
sOmiwKYcS3Mh+tgrn6ctyC0rhpSpQNYjgNhJ6CrwCNU6glCTAV14Ol9UanB3Ob6Z
B5uAFJFq8g2xAbZn/4p0c6QVFOqEXP7rNUYNqTpCBUulqokbulMw76iQ+v8whlzS
MZIv2Htbv7HfGpX0uxEkh95t35i9SySx3rYaxUyL5T27VciX+LWxvlQDrKCnoA0z
c2VPN1UuaFRgzjKdJNUyQtmoYXStbmKE4tC6Z7ORKrFKC8DHIjqG4HteFGpW6rva
Sh9bsGcDB30ydL0SDi02vb2h3OU9YZPL0HIMSJO1xTVuzm/GD/Vj7Bu3uBI0HWdR
SKFzP9dpMoqsgGx5irMZ+Bdng9sQBOH27xeCjm6ycemvZBB5jxZjKAk1kCD+V6fG
cbacc9+WNlhaIKK7V5o9MHxgIYF1qEerZuq2T/1Yk/JIWGTxC/MXXzifriNVUu7y
ziIUk9VKWu9Bw2E6XLiWvlwfEivla8tTkwtMnOa3MqbWcS9uEBmIIkA7HQgkWpdc
Yt2joxOwNzNIUQn6vcV4D+XU7FH140quVh5U97jVEau4TY6iXiMramCfLuHDPcZ/
CNaH/R16eDntjHCVOcW1UZ0YNirIVA5OAnOUx5PNbCBrrG1C+at7WoSCysizXuJP
Tc5mJ1jGLT3fbth/BKBk+1A4xmn+eby3BN357XF4HgkbqK4D39jLMpcK6WpFJRhj
Ink9peJ9o6astWlSKOIDXQ5V2t5/0E5ZnF9pLfY0M7r2yo5tp8fD0/TThHT6sgy4
rTRFH+hzLqkrq71akyi/5QB5Ymd0C2OmbiyOHTKT3VPRX7cGoNqTtC4VagzBcguF
jy3qx3oRDZWCsRna/LXCvj5XtLn0YWMJ3Rjx/6dn8P41bBRdiuKkGX1O3mbr+B/e
6ZQoRPq4Qr8zd3QrPDHff1FVOKYsAcxy4TPnAsMdpN7S2c5nnZGyz+OJT5D+ZNS7
Z/ljPYqoVuqIiWXkSoUhEeWpGlxzA7q03j2daizi6/29Mf3k9tpPZtGBKdXS4gDP
sn4Pa35pJXGGELz+G+Fn+KKASiaIOLyZSnzSoUE/AP9Mbd265LWLaK1vP665K2sh
WWu90srH5jJZlmsxSoVu7Xn1vB3MLyEscoKdwN+wJHwUtA0lBNtnZW6Za9CcuSvB
Wf0D88grQJ4QRvc/MAwpbjqeLGgyT862NOxJlgPtyZ+AKx6V8xnAi+OLMTyBuVL3
/CKFtjbPE9cqazXWoClAyPCGrE3toSjEfuVpfShWQ/hdo63A3VrJzUoVGH72O4t+
WbMLqGckbPmNy59DoBnS5tjkuHiKtUHT9W1evXk6dVjay5IwCI4SWHuzHOua2uSx
X5BcXAr9eP1pnsdinIG7YbldjvQ9Gtm26XqNJNJm3r5u94/R+Fn8oXPYiECKl58g
UJtnrUKp8diXxzbhSAIDZfcavQ/+vNbKBNHHUW4NypcvUgQIet/MXbXoHey2OPDy
V9SI6Vt/GlHD3tfVhcfmhus4Iclez3lki3SXwt1FpjPfwo2/hbO7SUXRLaQ2ndBi
VczM14R7M/l1gIi8uh7kNS+HBvgWw3guY7cPCbhkMxislAt4Ek2t08aRihAlDzGA
8rELLA8pJ/35iJPKH+AvaYSH771xv4Ha7vkxNy10pvObYnEwTwz4WrwJuS28RevO
Yf/sJyJiLqfoJGUqjSD79yEXgTj1Turv8+KTWlr3kn9xFUH2UV+UNDbdryYfot/o
S7bbUmGNWRT/TpxZr8aVIwJagOTdHSJeMY0vJfgOfUZFdVJ9BatkJ2CCKftIL8rz
HezuQWsMf0Ku/XQtN6nC9VQ0JsGqIXuWHh9E44fGl3N40nTk0K2thd6nHCTqj/MI
CJAQnnqODa2YCOVOWE/rJvhOYf3j9KNXEFilnqMnNSTFtUbB2XClxYGLoxi0t92W
ajeKqc+prR87Nf6Rou4e2qMnr/M4u7nmE4n23KgSX3RTPFh1TrQjUc8tVb9dzlv2
Xwzi3Aka5KSA97u+gvAv7WGJOBaZOwJNBhE+kbHT7QmclnaqW1k5V52OeLBAMoIB
LLO3EgaqrXQyBhyQWCjprY1xvbdMg+0n3W5q1Am0u+I9cdmKz94YvT124/9OqxUw
UdRctOIWXCx62anMpgz+RRGQTVl//AzXx6KCdLvB9kEK8dsUj+5J1iLQQ/UofrFp
5uLVoTLmMGCl6weWlIvoNtzlAPKHXevc6xwSZzikgCYW7fbphC84DokKAN8x1j4P
1Xrn5VwX81ISfNJbDX0dQZdwBDHelhP0rifcuQj81ccOcWWd6nql8svARytuUYtN
5R+mQhm0zmMdcVB+OaTooQCtoFHbjB/JUtImH8fkIJQMIyyWt+v/rCtgOwanJ1Bl
JwcVgxKj+Y58+Vp/hCLe3aOBUXR4mBwa3UL6jG3XL3k2p/QJRdmLYMlgA06vf2aH
hRxlcT2RmnFHqCgQKMB3o4554bXf3jjWeVHUJ568sw9IqQh38l33LHciW+H+ZsrT
0+llGbhpmtS//1cd6crgqCd47K9UjTbyU3IA4XJGznZ7aBXKyA3+GFoLmc7MvF4C
dZjxIFmKh6EYKf/O1xjeOmlvMhIRroK3kssbMwHrZLfFrm5uZFIKmbg5PRmdIjjU
zGu/3bmscndaxlKLolIV5MmKjAYyvXzXU/ljXvcf7cSe6JQjlhby2TfyB1E8Lr4N
52HgDJixYnLzrvXGRNw9wnl7s20TdU9NgnrIqqItbD3lAWhOBBm23ijPgUYr7e5K
xUOICht0EpYNo8+dyRZjnQ8OYlbrkIuZjUsYSjuL5aJJg4uVVV7rRe1ESS4EHe1y
CbMIcR6nkm8q1qO8SoagBx7qF+pz6Pd4Z7p9SZILqqerfsV3LPdo4lPBKezmYv5j
ShCejMJZnvM73glIb8R9BEqA/EcF0DN8bJurQ0YM8rrgsKY3No3pR4Y2MyaBvOSH
j/63IxDCX7S9TuhSAoi8Vc45dgLGGFYSQqgT8GTLjZEz/RbFFoh+zLLQxNlF1f5a
7F4em9fqk1f6tOKu+FhgU1nuiZu4qVaEiQJTUMu5YKH8szoSKYC4i1KcnCj41qgQ
T1vGSr5EbMgHI+k5cxNSfwBGXMmF4SaQDquEsAi6B7gh7T3Z6HMM1Cs+Tk4Kpfd7
QUxir97vm2Ds/qsSJwfJOGzqBVvejof7Bv4j3QaLg5UjgkeUjF7E2sESomXG9tOI
HJButDxR8WVI04pj/T+lcs3kF/ne8T5onFTbEWHl3XqvYqkuQA+Un2LXRhJPVjZd
F9KkvXBzvbReWuMSFDOpaOTz3n/VxgKdOOXazLmDRL+yf3jSjGxe4ZX7Kurx/C4n
cxo0Ud2HWp2vWTt9BbQhlzW+nG33C4BB/NvZEKGlfCi6Cn/A26G1NZ/Pg+GblqYj
nJDX0AwfnRrS3F0w9bfNaaEWsXFunP0OWvMRPeIurXqitCXoLPIU26HYscPVQWO4
CJHIwWW4Frwu7bzSYI4j3UfPpKjVTsi54MaZIZVrjRZwfqY67ijNvIqVjkm7V9wk
f4wTKQJIXtmTrqtUDu1dogP+jJcV5hNG8dbGmyH+LRYk+sK3vcMAH5mP2liL9AUc
4bKoOi/I+ll6NDf6r1fYf0PkH1L0Pyc3LePmuWlM5DIF93+b2CHWGWQtmYlRhrdr
wS9JlTUzGILkI2GutI/QiVkbxz0pOsapEUn/rm3TfcZy/ss5vqfQEOMkaJDgKJkS
li6L/mlZzVGj5vWzJDNiboMADZ7RNG0e/+Wf6iAWDxigVCDXA2YPtoR+PN82Re5T
bl4F8fTnzDd1iNR8hRa28NlqqhtGnSRv3PY7A4tjDs7g2c/6DmAYJMCmbnGRUPmJ
1RY7UtSpUaikrC1i2G+5ST0WsuXw/aZMCjLHI0MURTunc7bApb2/qmlxIZoKDEGC
ZeNaOaAM7tFPKqbuaWPFUHWDt5mg4YB/uAweCw88ncd0sJ4Iwu4v7513tMZQH4w6
vILpoUnaUCUqY9aF75yAa3os9kuuP10QwU61BC0nyXp6GGyCUuEWyigmUmnpni1R
CJGn/6aBpcig6wGBpEGNlu6uLLzIwpOdVpr5rAVAZ+FAKTGf4NXkSfwB+j8xnNQA
oHH2jl/QngdYE2nB3qsp0Kjflj6Zb3XueDBb8n8yblKpjZkc/JfYlOIYgrr00GcX
wUrwnIoDFPq84segK9DGSGNGRyYFoIzVdEqaVZT6nhGS7+lS2VchQYaAxANrm2oX
wFA6LSgVKaoEO8/N4IT794aZirurPgb2Q1Q9WmlAkDOb28n4Og/IIqrURdsDiH4D
LR+dwL/6JVJPaCKqMv1w9m/vGepeMfC1XveJJPkB6q1SKY+zqmJnhINlSTjFEetm
SZwPvsJJXEyStc1P8KtKGtTjq923z6ju83H2KZIvqMWieu0Jzjsmb5mKWjRj5TzI
E9H3adGKOAsUZX45JK61OPoy9REIg7/KDe4oyIlhPWOYkRxJJwHso8eo1RbeVHKq
c6LlOAxip0n21aBzkoZfNTJdcNb40jkavAejPME/86IU+eFfeoxqZNmL7YKY7IPb
Jb+Z64rcttNlhIjNFIMs9UckyuDqO2rdnYo6Ej3arngQxWIGhy7LQYyotBakwzF8
AjD4wN/TjetJZPfZ+U7quzU73oevCypKjHhyGbIA07E+HHpoxnn3ABdZSCXPhGWQ
/jcrRMvREYZkB9pNEibiboiWlbmhF37uSzu9vwJmydx1oNvXgyNd7HTeGso9K7Mz
GoT4Cyf6YqWbcXldDnXvA+a+hlLu3aG0vCgCAmhGcd0aJ5UPj15gCZF/q9JgZAlL
vJNbATFpOi1l2vMV30QKDxIF1BDuTmzt8iXyljd7LK/Fi0aMCwHFiMtSRJxq/u9s
JOwO7iLJ1o+Krv6VyXcER4khYSoUxIg5Tle+6kdYvffx4ueHZBq0fthWH802jM2a
tS7oDLHR+gNxO+Kx0NwoihrqKgQJMX/OZ0NzTJKdBAKulTF2pcA7PZYFpcz7FpwA
5Qj4aC16Mm7K78psTDY4rAvzcWjTtZZZx3c/s7cbSjDuZfJDXNii7jodt/NTMbaQ
LkpkzO+STnav0xwd2yHu/NB50hZ4Z9Nq4IDgEUMu1Nc6Wnj/W9XdGQ7NFMgSZt9e
VrQBgNzOskN0XCayWCZhTcFXmqyAN4wwBxjlfo+/KM4bmTFNDQPs5q1fi9mz3aiK
b0JSssWmyy0MJKMXqPwC2Fovmzrnx3ZQupw0i+ChcB81Oi47rIx2RD6JbIOKIOIO
6/Xdt/J37XHc3kKlaQWn9unAP0tnZa/yvGgf8H9zyy3rMCXj8ulipPOXyrL3hWe2
nwB18UxyVP3XLYmqQJwwW12KMy8QI2UxVIIj+4m90k0z/g9cHZPAD49k6H9NcoVA
sSJswglwYpsE/9ZOe5z5qeM+rxgB4WvWWA9S0TbRPKZV2phXm6vlmn6+0z3uq7BL
03/INwHQKaO6gsLtgYKKR+//UeGW8ukWzptCRJOXeObzaNd4fqqs+zzb4+PBKalO
Xp+5RTDIbl/9U4lIB9JK6ee4eQKzKVDUZUZ2R48x1p+NfbIHgGXsABCXRXMy33mT
6rSyEilkQyMOyB3JinuZVASILBGpJguQIFTExsqCRlkZ/hO6qexQGpVte2VBGjDV
iKXtmnQSiPmnmFf5bYNpF/NvJPM/ByKQ1h96dpn4QPwxz6nDI9g+9YHbWsn0sHOl
8GSPRTJizoJgwMXHAEiqRu0k6hn8WpZJgCTxqCqPltMpm5W+VPvf0iOYTnPYFIre
UDEbT1Lar+6fFxSK5pDst/ZoFIebX1BSFqAs39Td/RecMrxUHapQJoEd0xYGtk+G
oF6rrQyucQwy9JIQB5ro0BRATFUOnGADDJtLgWKvmaO131IzN4cexqfLf5ZLVZf4
0OZZjaW0FBGlMgAOj8ynjGlQTKW6dWvYd9wuIRIm0xE3uT50xg0iiX9xxiaKoESt
y55xVfNUgb5GZzU3e4upk9frgl77TdAUHTydY1xbYX7cnsywmc+K2X5NDLciuPFg
JbuOZsNA50X8+o9gFTFIERv0gt4vi7EEI1SEzzv/unJ9zDvnyGth7kfACQvyjtaZ
6xNXgHFf40a7axmfW8thIeZxQSCuYx6RZFW81nbG2mvYSdTipOk0DYusvhUlM8Sz
6O8QZRZ5rZr5xOPTTKSQ0SxZv1ZQFFChOdRuFxtTCYt0OrNCDGq21mo+KXDJOyPW
JnKLlmjXE722lawFza4ojfW+uLQ9A6HVZZNh7MgF9ATZLKQLLLRdYiaMohqA2GVD
qq/2XUENhRz2luA2P1a/4z0F6TTo7cWlsjkcAysvZ43X8M0jQZDU6GRHbDA61u0J
gyuqsXfLw9plzmKpdd2UHSFHAJWwfnAshfHNOoaDhR/+yo77zl9xYeVFU8mje/s/
fLw2r3M/vsCfUJH1A8DcapJpIouS/LU1X7LPGZIoRfFBUFTFTDxfjR0fgynk4FdP
/ZAwGGbgz3kPPYNPUyrVhyqyIrEwJrDGSnNpfhtLpWNpExAT7qMNdZz1P0QbSflQ
FqsfXC17FlC47buJl6Iah/tSYV5lJGVYOlu7PKxNxz+PuHIQ1nvQ7t3VCCWC1SEN
QYWfuw1ZCnYykllWZuAykWhlt1JxswGPoqf6bj8C9/Rf/nMtlhXIkZWtlrnY0unP
X+beaMWSdF5t1pCG7gvp58GdNcNoVtzUCKpy1P+cEcy1elRRmOVq2BbT/147oQAg
03mkkJxG8LqTS6hRaxjoiPnxCl6zEX9MnotWKX2H5yxA/7T3jqAcSvlgYYX5CmpL
s8Yokv2Azi9Ggx3VZTe6USqYzIGCx+9CWkH3u8OKwsd6XGSoL/FktWriPwhyKcfS
YqdVyBYWIITfdVh7E5TmBZefydo60eR0lN1YeB1bYK4xRvVndqHh+oF5JWdv8wLA
o6aXDn1ZnN9MBi2Fh7l3JaDlrYibRv0JbJyWYSSukxc7XrYAfqQSJYRte9cSDx+v
+FHvFjYwlTa5HbobkJTo+S6FFjy4Dl83cg6j0VbHQQSj8JHTBjDJ+zjuDNroFwx7
WjNrSnXpfJPqqjfMnhmm3GOF1jyaYdy/X/5LL4XH/Psn2ipQazxOB6j+71Soh9Xj
AIFZvXoo3oWHZcMzUm/Oo4kIWXW7rMWD159fNkJYl10348OGRbDNYgnBHU8A2W+0
o1y2qAf/xL+FuXVPWMdfh50AA834/22OQFSPtZGUd4Rp3KPY0JqQWcZ4KhD2VNt+
UcZ2Wlt4RA/7jJmKww1NCYf9Xpel+0Xqwm2mfFUhg4Ky7RklNNn7bhhnv/HPCBI3
kSC59FnXGi4wWjRX5f4urF2/4nvqIOVXb8UpdKsPSQ4t2YhZjhC6F2Em+4/eJXPV
pHTvP4to1bjm4nq29A0pZYzwaykaiF9vz6FObf7ruyhkrvEFq/yw4l/sTIuPsivG
7CDNfjqSXTBBbGaIknvSBwj0kEC2IuLrznIsY7/AeQ6UxxXXUAo9Nbl0xPgDeM2Z
Td7+gmBgEi4+hCkvaecbAmq4tUeX9KHTulUqNKaiJrZ63o1dBY8DFXWGTk4pfash
27IkS0fyyVnbksN8OvDzlhCjClwMOUPGejXqUHmUcSVZapF/TJKcwbUbqE2FENZL
9z+63a8cyEvpkF7N+BuzbN1r6h/Gnpskqmc4FL8VRBxZqfLSE++3zA6MDIVmO6nd
H5SxkDlJ/mZ+T7eRKtJCZckOCqCm6b/kLNpWD/DyDJAHokwDnGaOG/s2W7xGigNu
Akc25CGU49zzyVKnDEvSAKd532BjTCsEgcEZpEGKbYc+flpeBWuOmUi7jz7S8YkE
e3xYU2b17oz/davMdw0+5d4B0pnQuN0Cbdh+znNFOPp4A+VXM0fNc9vCSLQZEu2X
aFs6kxeuyP4vxNKmWWf9eRX0b1535REFWp8t4JO2AjAtOg80JQLbwxZKsHcEubhE
lECjrJQXefehUDlra+i1/7g6+Fp39UnrjN42oENxt2PXDNhOG1x+8QX4O/mwz+TH
fDWsx+PXxMkUtv7pniS5m6g1EKyNj6w3ZNn/rXfxxOxXHVwGEFr+y/exi4Y72oQG
iuA/mG3J6YtuPs6v0Ame0gxhgqXjlELCqFspnbOGdGSzZfhng9L1OOiuwljWBJps
J2alOhhI3cTy0Zfy5mGz3kSY/IESOjdH9qVasH2Fh+BebRVcZAOIL/HmzBuiXpU0
Buoo6yvGjEHSTNgQeKNZoeDWREFNDedRxQ3JTiIaWMPimYlSTo/EqDs9RHGTkMgj
HpOcvYwx8eY55GPeTV7xPfmPyWNkEj3r7KROUaVUPlqw/75MPb+pc4EEGKiBpeqB
07wlp17njpbs8mC/Ai/wgu8ohkuYK57orjtBQYRBxQt+3EcCUC5v++Z5ogdyVl8r
BnegV56yhuCrDzgiH/JHueEoZonXek43/DFbt4YiZlscI1JhbdHVNnNxpcDHnYy1
I0OgZeDcLItwLvrWIScrOcLoHS8M06ZDCYKkV+8vqOLZYWXoK91Q3M0XIA+6xSkb
2RkqovGKnSK08SZr88S9G1lCm343gn+S/66YVP0kbmd1dKfrqmghMvQUUP4WaHzy
zgoTTGVyK3RAFv7+NWhvLs48pzrJ967EhrD7MGX65zic/JnCPVuuRAB4WnQSK4r+
6OhZDFkwd7Rk3BWfXxp+AOV9H6Pzl45LxeonkLlBKJN0mbx9INIpGtD1LtO3otc1
2mS8z1FHQb+r9omzJIi+yG6CQCt3MPGUKraP2i3Oewp8CSLYsF6QMZIJmPBC1NQH
pnd7moyj8SG4N6cWQBVlL0ObVRAfCEIZw+Gc7xyrnE4DJ+rjvsE8VZXhp8o9/HYe
U8eDN4Viqi8HQpaWt3lSicLH2m3wBFcGYwAYJxb1BAXLqRgbl0+a0XxCEApMESka
IWcauxJbfckvvRjDi0lLFOco+e/S7BK0i1nAHuDJcc1QDFi0dlVRWtNkVdTK4+0C
+z+qK17qy4hLZNqgj7CwFo4pb9OmDnYtw7udeZciEDRmhe18XIn8i1m1udPTfele
QelLbXkDww2Sr5eSad7Z3pPqa5EnE+HATFz0A7sNKW7irpzRQh7LKWaD2r358RZj
v/UKe+RcVwrDH0komMxkkWIHNcbS2SuqYCMsMLseURpm9soX8qeyzPVt3q+JA1da
Dk/WNe5sHjgCRnPcliXIj0zAFDuDdUycqk5ntRCAN8sCVeiycYvC5cXhVezDApN+
5Mg3SAfn5xLojeY6qaiwYIRyMvQzDPp20SlHNFOKtsNX73hqd7Q2kugSnKdC/aBk
J7LxXyF5bAVgYMGn7AbmkhjEPEwkeWi6fHdsuQsIAFxwhI+kZNxxSk6p+XeWoEp1
huuxoIP1gYNNRsSZkuKGLAeaMQaFx/ywtrgPYqNZwCrLyyXcJ6X+d3qv9rofb5I+
0hPIS6WnUuHWSwr6hds8JHnwn1Uhp950XoNppHidMhMCJDxy9eFSSVKOlKDze3Md
dsMadOWHVQCau0eZ2gqQtevx23iB7lm71pzNekHWhbqt3uUtzJ2Rf8tPDa13BzAH
wvQGu/xjEJW1KCgFRqGpD1sRG4MH7xTVs+/YiK6Cv4WQZaZhriXMtY45OX7bdUL8
SBfUD2EmlD0I+txSd/BKiKt2xIIBS2kG+jJ53XLa4c4Ff5iB/kNSYOjqcUjcIHXv
Y6UZfdBx7s3J75X1Ye0OrBtyOC+ms/HySnBlz6d1pQzcyXmVEYKyS4np1rvXL91N
rL+pBX6njmRM4tKSV1q+J4I4RkZYf8fMh2iFg/9XV+L3TndyaQaqRn5LEbosBmzr
MJsFWxTLK3kEj7rLmZNL8V6BRqId+lgtamGjjO5OoT8ap2SHylu7bN2nUaYdcDts
SH2jKEFxiucmShL55+5VIODagyS2SBYBcZm0lC8EQNFsXBa/f4M5vQnSqBkHNqme
rAtuZWP9CmAt4biniw4TWdnZHPYoJek0X8oA37OVJE/03r8dgPiKX+jV+0bNg/H4
XeXHfWDTIBzni5bu2yA0+tRLIhHCXjLBQccendAdZfTIReeantmnW4H5dVS1Bedi
NWd3DtzenJUb2AHpI1YklSLIEeSOn7YXnw0TIQ4LnOYywHtfneKrF/avKs3GTjgL
WJoF9aka2zCP0wsLl6J50u5Ta4QuZq94VVTHmqeB4b1Mb+Lr2VIDOnsfDBStyDxi
ozrq6Om7eMk2mPOfhP+4Omk9WA3ovWiRa78PkN15GJd1CEq14sP9oD04T8gwZZaS
yv2KbrUF75wN9JfbUuAVVYmW5IrHu1cy+ueQa9WpCOBZ+KWTFjDOuL6azwHYyJgj
7HH5Puz4jErPWGyazySsu4ZgcNc0aGtGt0lzN2hQfqfHd/A3vHH6Kt4mZBP2CuFb
J2yP9dOxSl+/5eM3MBPYCbw4z5OCIt73m4rpZY+7YAbk9E//IvUVjSGqF/kxfBpL
LyASQRtsaGKlet30/V4xwEswn/ggF2flcB5a2ndY8Jw5stfwif48734SMIs1JJEg
WoVYAEATaXtEQ/w9lFXaYRD+vLvQJwqDbGhJIDzaisnvyj9R+NZoKY+swedyDqzO
Wuqd2o7foyGwcEoVDw6sVBQevat7LIvhtPIDgG0YyZxuYMUFsgX4POucGigPN0E+
QY93ihICMx7LSFw7XocqfhcDy4TrXGClBjW4IQOF4vQrEVveTKB+ILcDZS+p8zsk
X6vTgCcobrb5190BYvY1SgNOe5t1xbHdQmk866LcE7Tnhbh9HlDwMjZvTH/SBFKJ
saRyx1k7ODoeVjsQesWxIZAzV2TCrqPzlCe8V2j3L1oazW9W6boYCCK3EMqWOak6
su+IDgSuIukEOXrvfhSmvoEtSRGUZQri4Wqo4p78+6iE9wEbi+4V6q+I01mxrnK9
NgH1HUZaW4UMjydmEROrsMVLXEFhFUlMczDpaErrKz6XFLyuCObbqkJOx0FKZI8S
yZF7076nD+XW+J7xKjnCtKiNgYrr0jnvlAuOPTloOM+NEwK6QzVVGJenLck+edyI
+FG1iZlzyKwjaeh2+ypt9bSuRSnfuwjTEFOEk+kifd87kP4OFTWY8khhjKAjYRnr
g2G4vn+cLDbHkzDBAumzlFkFLkJqdoHc6UILLQ2056e3RQRnTyrUFpJYxkalyUje
QZ4/r7HhPEW6dOTEY5wrJHDZJhygfEfxSxIHYbC+4AcS6Cu70m/+yerv2M0Qk8Gk
jrOCy8WNhgXKgdzN9sCXNn7OVqfzcFeqLqaWsWBqeHEGy4qiqcLpNnwVdDJXoNul
/uUJOzUWzN/y+GsKCuTnM+wopIqph7WMMMO2N2NDBAgL9NOyXiQAqLvT1HZIYCCt
7FMd0odbCACPoIQqwofrWkdljEQkdIzMhcNaoKb2wYO26pEfMjAFITEEKw+pMBOW
V4ttcXt1Ktpoh3ziq22uejlYLDd8v5oNK+qpUZy+gEnGOwB+IU1KUVhexbelbxfh
5g0c6lhWjjzpqzn9XZmyW5CAQH6EAEJQZGpjPvkngTFZyrpb88ab7345C/AjYVlg
d97hl3SPHfAOWJtn8ZG2Vbr+4lpfkxwS9cAhSOQm8LOibN+OoZYHG4IF7CZddoOX
AWWLmC7XSSul1RzIeTkJgIYH+JjMGkmn7PVqzaRSbTSogwdpWRAmUyqE7Y4VKRPh
H/P2qtyLpymQkApYbpoWRRZu5oM6Qasq8dqYTi36AiAKcmt+xczxGmtgivwv2rM4
cOnYKj9c3XJBIHTu4BrywIcGaXw7p0ufl66Y7nz8LZyFVskC8OkTSF+ro5y/LCNt
w3QBvH6swvLovy2apnvYdPG0fFnaJBwxNu3lkbXtb1YvWVHdJKVleN/EmHhzNSct
syZ4b5roUG975/z44FwoBl9Rj/Suz/q+6ZAM6rUUvdmtL/WrljuUD/6qqdw8yqxx
gGJeVsadnhF9wCHPQvbCdfN2a4C9tcQ9eYnxxEGhlRJSngPp6TA8BBk/HRqWMyIm
bOt30XvNYVuw/9w5bumJhIXlVBR1QZfKkPvUmbl4KiqQ84ZNHmZjhJj91jv7oZ0m
fHJ95PYuDpOwRvjVM4ISawGGEMq9kRBY6SrAzMkWpWD1n3QpG6I38paVtizZhxC/
6fwPu2RTdgs2PqvFjFK0Ljbwg3JwqwFn9dFP5P7AAvVH356lCmZlSLAgtsR22Qy2
HUd5mrmEPh8EyhleSYBMB/uhpDeyRhHn7hTEZaHlT/OfEMIWa91e9FxoURc7Zlmq
TXUpTkouAndVDMiHn+4HaSEF3T3+idE7vthPh0uY/ZQhqn/XvmR9ipAmn8Had2Gt
osHCG2e5HJoAomPy0FL61PcElA/LNN34AHb3pGqpUVK86SujwNKbiOkXeL1E5m6z
krVr43RU+nqvDGK22e/PtVBI7olnixA28weKPmSlPsXwWC9gRKngKeVIWn8S8DGy
u6GU8kDzQb7XV7Y+fBGxIOzRVt+5TCqqfi8WXSGCaZVpXdos+BFHuh7MFhLPcYK2
Cbyyac/9nXz9cCRy28QMCdwU/7JBCfms3Ca3zxMs8JXIV1oR6iQSZ7sbk/mw0jpS
p8u7eHVlcChcz5vDcFfNQYETpSF103RcKUVoktyDLPQi7xBJwAd01g72OCHFnXTU
lzoEracDgKaqcTZXnolR2MyXP02LJYbny87qTnvE27LgF2MFpToHupeRT3tRogZ7
EC44lR1YV9MGyQbuoC8SpjBKLmVqrGrMaMPBRKwVivrJ5io5T2zG2XZryRw/uTBG
PQfahL8389griCDuF3ojEzkLdzYvwAyB3Tzw5VrDYBd/ZKl20xUhdRjePqyUMyEO
xCeaU98dIUmySh47+FKH/keIfOnKZ1xuw9OySGdiYQR4Gf8jpMjoh0YAUhD8kDP3
xQC/Di3MiEknojz10+9N40dninQY3ZuFceRngegrtcY6t+ny4TguF9/l88NLl74q
33Q1mgTQKfwB8UmTrxT2p/KEkk4x30ozGAuf137m3RZ/NFPMpXmWiFyBSF9/5MM+
CxFzK4Se7ksWw4TajQKDQn6bkDdJBkMrDjTs8MCQUrMyr/jf+RR5Jq6yCTCFhFet
z/UYx+hSJg+TazoskrzoqGn/c2i+hzsjM2fp9qdYbdj7HgaZfAP3aG4b+eGD3448
RhGS837ksUbwY8B2fO+JVmuLzAeRt7FFDkuCPBOuIRXWa8igy/+ePCcL4pr1DUEA
xleQHH4Bsg8EEQIeQ7mZ2UjbQMjcYOWH6ydFV4srT10AKjf6Bv9f4BxbvkdkfKUb
KxCPrCgjDcEi4PCDU7ra7W9goeDYv3oGmyoMySAaFMoaRzmmqezlvXztHjVYTvNK
wy9h0K+0xtLCqxI8bSNrNHE7xkEAQjCOb5+hECUosbnwqtpLr8NQ5znIoe+XzBCS
ZuULKu/CE6AV0lX2RE295kKm1w+2e/TMfqIbKWVufhPxL0+3hs7Smx+stxCARQZv
MpECJupAaotf5iKiXM9knCQNGVmR9BlZIv+2d4lgokQwGfNLENLmm8q6HfLqXE9q
gw5ShseM0StALcV46D/ZwBe+TtAtttoIcY3PeatC0w7VUIZSQLh5jg/zDb7yhSrN
Cv3ANr+6UPG6hdC/hKzGEgVy09Lebhw+6kh91z5ZK4rpkTUK8WStbphgznjJc+AX
Ja8uSBIBACHjTkFOKZuCNhhPubvkVy5p3HOMaPHYSfwpFvNTZCg9vNw2Z1Dxnx5e
xzg00YxFmENdhLH6wxQMLmfbEM9gGYgkeG7JTZjLirYT7f2jfALXLh1DqsfEFkQV
HkdhmpFosAEJerhXBv9U0DZGgoa20/bNjCEDqQHasgNuaXGX9PlLNUORuf75pHCK
HOc1/dzG71tyapXzATqp9i9ELNyX6VRE09y0p/GGwnVjUI7UhhDLlBo9vb9+zx+W
YT0N1abhlDmoufAj26g1ZlwX9o06mU4cEuAavmPmjMhkb3qVHt8joPdaB32XNrtN
skEcfCOnsNv7AzDjm++6HQkCXlvGd0rFo4kLpW4ANnwOmP+HNOhYlzm3t4pex+QY
zUip8S2y3u+lgCd7SJbj8cbG9/vrul2QPdRjHquF4PgnhOO0l1IX8EQm/VgAtb8W
Oh0sQQrizEdQ0wqFS5foL3uv7JBvEYiQRm0xiCxRS6GjA3QB5/DWftvEDPcKF9pr
NKPeh1C79MaCWHwWu/XJJR4umn8/uVJP/UHWyjgnx+yKsx6s0jwvj5AKgByQNV4g
INGvkuwZfSSSq/Bd1qHVVG4+yIrNfQdzozFxGwhacesuKpVe1VOsX1bJTtf5XmSW
T89mkNetzSfElKBvIHzrZJSw9MeAyffy/rSgGsPl3A3+VpGEIx2n4/ONlIqjAEAI
S/AoIuN6UnFO/Ugdjlgwb4s47LwDYXuF7L9pYNTKnDcc6zmj9ui2UGJmE1PdAgZz
xtf2O6l7YOXKJFEB+fWBv6lTEGFNMYlrfODB+QuhrMFdDLzfQsBeDRQvZ0aQnFPp
ZXdcutVT/zBUaUhGobdsFrRY0YASqlINmAUrM7/HDyjpqfg5SuQhC9lTuq+2MX74
yoNBy2A1ouy/2TmlkfpA/aLw2O1POAV7prpo8p41wCXpAxAzpLNnyyajBUoxiRh4
6x7y9kbV5dE0QhGhtlOg8d9dTb6I955BEdXCiZya1TQdODpLUSrS3wIJ+Bc4JX+M
5tSsKyxVhyKSYOL/e8erVEku+fd/teYihQAEr0rhvf5YtN/n04utZ8pzhqj/lYUU
nKH0AdYHFVLd4lZO96xRg0vwn8VQSc0PF6/5JDJqnD0rhGg5Jj8aAK9F2xldXOea
UuxjhQGqUiLGV92xwWH/i82RfWt5uMgp8K8xMBWmsYE9Gl+Lac9tsa/zY8/EtKlW
+JViSdUOI5zK5SxTzfEBjNWi3fXV2HkSIBAY/EvsIQGBFVQbeXR9E5EQePHZvZhe
4IDb8J5mPIESefCEdQCIWXzmoKXhbyOned8y8BPVeP60v0Ep0lI3L6d/rztyp78o
Q/zK9XZOP3vZz7HPmz1kGqmorgojQ+O/gxIv0LQnUzI/FLcMUM44b6n7WfhpNNdK
tf6a6YPRkPvdEpv409EP64InsLr773fB6Wi+D6nlJ1nkWOYV0ObllT2VODq2OXHf
fMCptrP4KRDaUIoe1gTmGimWYRNgLXcoKpuVUyW79ZkiwZTq+Eyf2hz2xE5xOwar
IOleoom4pM55l3dFi+U37UNbgtYiTRpxlim5Z2CS8zVA9D+Fmb8hg2sb7XqR6yfw
PrwqMMtosPdGmDmXfr66QRUSEtUnJYq5jI26APQSvD2TdWvHoSWvihBmB8Lgvw2L
QHiSutRsdDFJAcmngCMwBQg1jYkkNAOfM7iY+zAqY62/OQLjcHqFIHXcyDwX3ATr
u8+oFj0EAAAjtO0xjX0YYdk1QObD6X7xRfuURma9k3hgSVsQU9bdjf3W2M5Vng0S
nOre/IjBb1G5LROgrcEDejgT4vbYtTMp2a3ILU0VuDamciY+Nopct65+thS85EGb
0Ec9nLED+319/6i3ihrZTeQxX1UqpG1EcTUI1d7xhAAw2miGvZGb217h3uE3yNkB
XdY/wSVy9DQBrJEth+UOVYnuE+iXRYUK4R7pLBKNhD0h8CPgczwD3aqMI1qFevaU
DZpDxYsjd2SULWW/ilii5bfglrYPIyFQ+NlS0Hn1l0D1u34BY0Fm+W1lBge6sfm2
Z2h+ZfRS93qqJk9/iM9vbA8xP6iWJLqJLJViDT4XiLqrU2Rujy/KvLXZMH8XGSz5
USzHkK0gi/I3riEpnlcj53Sv6a/D3/Jvq1Qq7b91g53lLCxkI4F7W6TqYHeRrg+e
CQH1eGcWCLjNBY47k3P3HTkY3x5cWFe2v8xcOyTrJIXuFmGD0bmljCkdbWSMfWm/
ZB8SFfjvzDfr5Hix7SbqemIHJl2UQQrtnbOrwiUVW+I47LBh1mdjzfauSfwV4kSk
dOyWKpQxQZMSh3aEViK0aTyaBdpxlBJ5H1as2SPHXFfQT0OGWge7sZF9ib+vk+ab
yDNxAE2wkjZ0avi6UwIllFRx8KjNsftpzoLIQjCSvHU0vf8ivtqCxGfgCbtRQVbD
AtsZAGO5+lslJPQdYdQ48bHz/k+e9K5JGYml9Q23AU1hTfmEaAyQRqvUa9fJmavp
JHH8AgKjyYTNeMLl14hup1dbDFRXK7F72WM9ddZWDlF5J3fJ1u9aPqSbA0YByw4n
uprzE3kTgx/R6W8wy0IWmKm2Hqf4ARrcj9BPsraw9Ua2NBO4wEyfJ/wxnEzgh4hx
y9lniUmm1JrxJ7MuMCER2HNPv1O+lFrd0kM1XaHcwiTZU7EGi6IgMdx1Z/q86mzK
xQTz7VFgmg4Ap1V2WTYRZFZd0Qgmt1AS+hkD21dlCLqtSdtkc0hRm8f09mpGBZgu
pJFkid4AxOsAHEgUA25WjJeANLhZapUoqWm4MuyCPHqyCt2SFBg9LRPf/PDF7P5c
YV5ug1zutJuS5DCaR/2ni58Pnl+PN7BLv/DeOSGUNFG1nlA70AcYAny5R127P3pf
33YMTxNRjUX1/PGArmtfJSNqSmHNgaSqx54FtJTSdX9MWxUXdp3vSJbqOmcWz9ip
9wOQhAlFFA1jmOmvujhmjZZ0aU29MvwBTnBChU+yiDwXApjn130+1yYISIaJ0a/2
wJjoIFVDqbhfNlCpg2W4m4Fq7OyFkjS/kZSEWDwzUjwfYgx+r/f6ooB2Y7faaCxc
vG8DvumnXAuGQDGI7ZW/6QOeRzjjk1UyS9QeiQEiwa1RkmQI0C9lyRn29ZsePXHP
kGbl7haUsjveTYVvtO4h6eMtLl/eucnGKa9OpZJiv/qffXJSzP7DmagMl9aJSadk
iunGKeOyYvLrgnxHv63ZDzkqxrJEkWutzBXXAylZYaLlM/NC4PBfk8iEcUaZ+Ea/
xGCuVas/mbRJ9i3YOfA+yxlXeViEIR+AWPBd2IVKY98elHC9IkzeQHYNSF5mJI3j
4x1qvb6kXWsuFTzVomOcPTQvcrn1yUhk/Iyj68Se7D913om/H6Ya6hk/WeQIDVmG
d2SWyh8vGfmfnFF7pesFPUk86cj18WnXGwt2i+vNvNYdTipl1Bq9wDIcKz38Ym/d
OB4QiSnkTwPPa8VUmsnyhqIVIxOBYavR5Pn6iLGefP+XF5OVZ99d5fy0HRM9wTxg
zHYEHxksohKdY6FYPCPob2GoQcOp3AEVVR+e17oHeanO5yDXZvrclyiPLDrR8LzV
S4afkkXcgbb71NnK9QfUq5BnU2sgZatUWdCVYThRzpnxTfM6fRn9cUNUVSrUnF+r
7R3l09P93ij1qE8ljN1u0P6sCDzcP5H0mQf0hvYmuxWP6u7B6NEc9VOwlxbuvkoc
geT1nDFCqFpc+RB0ZUnsXTOizcPCeOmG/EeRtGA2oKN17wEjHlwSziwHbr5AfMuc
vup72r92ikTWNj7VrUTI9mKjdjHSXpTWWf5C4xIHYemO20Q2XJX44HM+K25cSKRY
YNRLnoNc+VetJ9Bo4A+d0155q3dQmYbDqiRUXW0Wi8/dD+xr7su9ON2Pb6LrOrL6
sWbrGYDttU0sGP33QrYZmOL73dP9fHsuaWqJEXhap2ZnUE/cSXn4ND3lsENo2IFr
Pgwt9puKut5u8VPYZnBVMaFSOhxbVSbkoKnTfTxTdQ/zFDmsA8WFdw3i7zr5RIol
cYcfywYlKMX68JSbvIzImM2BH6WmxrJ2CzsMMWSkzW1WHc3WGPtPhuWRovLreVwS
ptL8Su2EvHRGa/n6yZWsKa6bXhEQGxF48LOa6cx4P9y72nRHyd7PceGzf1VdsIuT
tWN/DznzYuns8kBiufI2qK1acfVsnCM+9eBXY7xb4N2JQJPDn1L0DxzSPOYxVzBr
VznPJ3sNVC5DuTIGscdd5k4DEIbn6o3sSm21l7Y1g54zLlWLLA34LQX0B8vXo46z
+r6aUTVU4F7raG4EgJa+qStujfsOPWSZaVBAZ1j23HeBp6pdZMi7zm8P76ts4fT9
06eORfBTh3fFAPJpP2J6fZArqx859W8ytCAykSsrHRHBfNm/uqE8u5NsALQItcCF
mmLxbFLfMaN2dkpYv2wX4Nxh8aMJvakSBHcOJCMZBnZvX43Y0vvV2bwXXeFtc6br
TDx7+56z7Hpm7VyMYF1iVTBFvYz5ulbM07c9AqbT9n6wulsFRfNYyXbc9cEyjJAv
jSl7wv9wDd2tPc+KsiIkfCnWhoGgcZE17XU5lxNwQNdY651t8TNE+EKh3rVYwGhp
yRoKGiEnBQK5u5fAT7ZVdKQAdCM2mdRAt8LspUENHzd4gMn5iDTHDqXE8Oy5DXrC
H5BRilMElw7NbpeZlGhD0KmVMvcx5tRKEDt1z7B9SGK4ilmc8ovlUS3tbFKe922r
Ush5o77brZHYBLQrQyZN2WzM6qsCzDdoULyH83J2Wan/zSxv21E1tzBq5SWHN9Pn
s1xcK7VlNfgauF3vU0pkLE4492Pc9QDsfc5bzG/UiL+vSIghaNadrqclHlNbPOrU
8JzVYJUjS3mYq0T6WXEbSBl8s3/7UiBWWb4abGVXCUcnaBSTxe/oNf5jiRgqr+Rh
Oyw+9DwHvZtgw8sbJ2fotdPGCpoi5XuZaFdQkKsWi4ry0YpMLXwtzhPriZGdDpvP
0p1RlYsdsTKstA6BkGuHVVz8LJVFrlm1CHmdMLdGe7Azdlf9adkbDCdB/eZfKhgN
7UtdqKi+gwQnCKr4Sz5h64c0OJP0tQFfrm7HrtAaL8Nf4BWCkqDnpzeagBPUNGox
JeFDLNFsa1cnT/UZfy5NB0mmVJunh1mn/X26s0hyWr++97bD1DC7Ois82xEDS4P4
PYdqBNUAYj28d7tcxrOirGCxsPjRW/OMaNI/mQA3WZqoAZLUggTPu1wQl5OynLY2
VUUHHgkqQKEQvhpjpHWpysgCsRNbBln3fSNQ5ZFsMlJo8XKqK1XpViQEgKxNaOcx
1q8ginJCCw99iFsfaUFrZrSN+IbEAM+scZ89kmMsLiDR6oA1iKvPukntnyXs0H4i
O0TPTZV13+k7iVHLfwsUe3JxjoY0lU7NTypHnbwAXjaJp8KcZ3Mt6K8AJ11qjQ5L
BapkguUrNLLkGcZlvj9xs81WJL+li8HbMam44aGd8AQSw6rNcdJj0HJH1bBjZqrn
pKcLC8s4GvHz2IerRfgfyeFwEFckUs+sE3o/ccMmy0FR5ye0asWGa7CgEmSlOSvm
9QJeNH44SU1P8/1T/aYcDAOp1Ucf+kPJN7an1GhMuK6UBW1r8e1peiMo/w+wwyrw
IUiwlaQtS3yTr8hKLWX5n3+VmlsgYK6aV/+2YweXnEiz+LyBrl9s+M1vri2q2GZl
YyBzLjhDECFS0iPfNwCP9r90UwDdwB54qezlasS8MQQgJgDK7f0Fv/5XEXg3hMFI
cyPLeUhNWNb9lAFxs5rnZwHR8pduqtDBbTAENpamsXTeyqHADTgEcsIwAUclPW1R
DWStgQDOHpK/Ndyq4oM5XLKK89fO5BO2P1j/auWCSp86QzyuFEFDnP6TxaRxj02r
nef9DGvIs3bmBdx9WOC2R0oZX4ThrOUf9iWqx4a82dBc3h3roe7wmi3WKTwVxJFG
KjN4qp30V/0btMH7luOcg01UXJr5OnhEOBmXBPt6iC4z7tx6P3u0Yf8CLS8q0abx
MMDZlkxcBaqTi0twOJPT0ax8CZnwV9j1AFJ0lPnoolvlovcREod6lPO4WqVjvba3
jb62P7Gs512kGqQYTXR1CGLIKroHcjm6xC79PINDnkngy/7d/CBkZsthb9CFdm/6
YYkFELltVDXSVbApFQlau3G67udbUESJne8NVQaqbPdKedY0r8etZvlHNXhT5qvX
kA7AoQYWSq2kfOBi3yMpkwC6clKzUUhecLKlA+ILJn4XjBzvPSWJ9kEE4TWMqm+k
oAmuFdbw4Yr/SL0b1gp+rhtnVeyU5dv+85QHoAYSGfepf+p2rc9FJqB/zBZtruxk
u32OTT6CbRjfbU+/erTfPU9d6uScV5FPwWH6Bfdu+5xLXzFztYTG+8EX9PyyaZQu
MK2vUHAFjNTEvhZpMXyjxj3j6NGrQIVYk2Ag1U1HBXuJEJrc2HxemwdIm6TAIg99
OMy6RSj0fLbLumeBOfa3Y89X6/pKH9U5dvl3E0B6ZsPTOCWQSUmGtRssRtVO/kVl
m08p2HRKZzouWqQW6n1XDnbPfSuflJXLlqa8NvS2VobMPX3dO4lvMe56hrpJo6qj
xu0N7Z0rZLVk8sYw3RJlxEVsDjz8a09/QUDVjCxl8lqNaGVqQiNerAVujXU9n6pY
vW8M/fD9fh3ljeqGbegb8xwrT2tGaWBLdNEutUdKnhqcbEovWgm3sfUz1oEbzaiM
vPa4/zXvcg90XsDEr67XQBVaSsQSEh6/nEGcDCakUi2UYW8z2Oa7qHv5JTW+N39B
IjXf+K932Jh0sYNh8TNoleP1g00f9SWXZ/4wh6Ot+lLCxTHgfzBDLpciskawMeWz
zfgyA30ENHdqfr8/Vp+S4BeeLsFiNIkCbE5F5WNBhmhhjLDULZcuMJZiZ04zu6MY
VTFII8OjOfnhvOO37nojW38JxH+w39bCu6OhHGxxQDriA6lRWGN3Urd5SZX5uqfO
IWlys7YsZ9WmaEBR9SLInFK15guQpLf6M63uPnDDbjjA6sCH2Tc5FS3pdzwEUo5L
Sl9XeoHhH+0tojj8XSjXf+fbbtlobJ+z0J9+P8QDeosyzdoXz4RTak2JRJWnf1s1
iv+05NxMJWUlLojNXRq0W2Y7qN8ju3csCCNrfZ8mWOzrgURyHYcBE+la+A4Ao6lx
BKAE9rv9vQ5ZAmHL8GExCtFDNCOayEESy8/wonZvCZ4hq+/KI9lMV/gQ64vD3OV4
T6cqJZc5Kq7JXrWcZwPj7DNwLPuzoXVxRpLw9MApj1B/4HkLfPgaS3ErCMO7TSrL
oZTAuDIa2DwNGlOjmEez8x737wFDJhVTxScZGSSyJBAx5Oa9HD9UAXGJKjN47tZV
7liuRxGDSp/8UO0hAaS+j90dCY2TdUfm/78zEwmB67A3PLgRQHGbQ+CUOOJBeuyd
t9v0xOJ+IebftG0VBTwNfsGRWXEN9uHxd0bIcJmaK7N9QlbCAFovxjC13VpCTE95
CZiQYlTrCD/GmVDIPediTQ5WB1ylCMXy816u+/fjajv1uPD+F6jkefJeRYUUol9F
HT/INNn+v8v2cPsEYMHS3I4MYy4/e856S6BE7GQ5TAHx7axUbgdDni/5Bi3Mfd7C
RKJHS3nH6HYxh+TS4AG70OsaSwqF9BCvDKvdwpkp2QibAJ4THRXgyhCtv+hRYE0L
k7CfkW/acYLGguYT1uDnfwgJHsI2nvj2vfuaXUcWmUpZtWp3r41WN8AqPfdSsxB4
KnUYBp+h3LYqTqcNrPkT7BnhtVyErkBWjqfA5FFJPOm8Yt68roLQ4ddV9sdNsKqx
hh9xlSVMYcSWlaU+Mj+6UcO0lAPM4UxKlipNTgko43dQXWgixbqjUPUs/XH187iN
rDbtXlB+sLfOTCTh18jD9QiXucNv2YpJeqDG2/Vvw4hadRxl0zNo+FVTXFaBhyf8
Yp6zYW3sCmgYIg7G5GGWQjylTCX1lHUuZERQKRDTdtR8Pfpr4LZa8JpL+GE7dG+D
mJoimebbI+qoj9WxgZHPVUilzu5Yo7saTUnu61Xu6vBL7n73StMyCJaahCbBDRY7
jCGqaBz1XzTphLH21fbPTM4gEOv4DkyLJObaobEXN/TraRj1l2XLqnyfTsPsvAkh
SVG/FMi9eWcsx54+OBhlMN4rCYcKH8YdbbPzQKa8lclVCvoqjV/A4ezaw3gaqRYS
UWAFm+WeUzeO62ANPUPgkkorbIOqUDedgNwcR7UwkIv1qY7EvrlUhECee9KuI3JT
vCY5gHsS/tyDRwpe2PoZVqsK4/w0H2dauI6lmHISR61d7cR8DKP3Tx7ZsKi55Zfj
hTLo+0+R3IBw6x87eCgxBmO2iY9hd7RDjd0qFJUxoVN0hvFXbzysA/3fDsNZYXrX
wiVNKSNBWamYivzRs6X+WmgK078gQzEiV++9Y4pu5WKdpcaP3OVrS/Sl9ZBfACQX
9jPkGkXmfJiJQB8Ru64z4B0gQGbvee4N99NZsbT9t7ItGJFJ01ZIRgZygEdu2+em
HBYYGhUVsoNpM2h8TbPiFV0AB3ldYac4YovxXapTIfDVn1AKn1qk0Sp6d4ULwZha
/J7ciwctM7MS6QkMygD3JjSqg/Zpy6zadWQ9eZE0PFmDhdHSO0j3/7VTp0Ed9Nwy
c5XRzgv3MsczZBmGZQbeGpSxXuapFShA+akpgdU2vmFlTplpm9UjM+HYIbdWGVhq
PMT74g6H1FKjiioSjYOj9Tu6bGEriCXhWDZfTdG7nZIeGlnV6Gy0/cOxmYBveHz4
6dR1tDdvh07v6EFHjP2FGlNFPEvixmkhuJU7xpD8HW4JfncmEE3LTAAi4QfM6Nqt
fc5OZkzeszQtR38kHRRFsXvvx4VydRgZdyPTPTtFbPWCOT2paajTbdp29Whbtd5j
GBnX8/KUKMdOfq/r0aA0Vfqh8qed4flVAB0qo1+D///EfI2SRzWu90/hqF9ZrHrh
lFLaa6uty3Km0x4lM07Ju9GICxvreX01+/nM2mz4Fr/3GSLSbmtXnmQ1X8NsSnok
UxPswNI2sSvcORJJsAPVdWqVf52pGnZf+1ziQIVhShUQXzHuKZHEyh9ugAs/cfgj
6lAutfLMz6Y276xsH278SIOEGvC2PHa19ErkHp7SsU6hTPNYYts71PbpXB1aJRSA
QY6lTclTfH4vgmME1CXhmZXR/S24RgUawjR3+XIVHmqlK2uVmRN0fOdaRt+Mi/30
EqjtN445ErdJZSv8mhRJKwhFiH5ndiADNKkGfYqhXSidtaQmH6ej0ipMn0FPSZhe
NPf+4tGYcLbLq1qRfk2lURKD6YipvfJy+PCOO+gjAo38Kx+jK0bOswnVAul2qQFy
dkDoiLmJn67bw1hniefmGwJkw7aImkNYRi40t8yoQh61f8t/wAL5LbRh0RLXiGfc
LrStJqo6je/8dlNRj8+ZPTxY59wlhTC2bPJRHjK9TwPv1kxY+7f+whgqX9hyzpuH
YYAdDVA7sZiUbGYkeh6inZGr4f795us1sHPft7BgE2HCCl7dfvvAby0qDYxuWoHN
SlLRlc5lmtbN8MyJdF6bS6bKOri9sOEEbeGrjKzzNPpQ/0a/ZIOLVCYLBcoPbm93
5bp7D00wlvQ0qBlmT09xgptkv1o124N8ui9Ea8GfmVQoRW/SwpRS/Q6lRTsU+EJQ
eYHuXgGgN2F8pl/ZAjKmS+wzMHKswAi8huhWjIO8Sk2vmlHJoTKPEYgOjC+wcbUy
0CGjdZnkq95dkTAXi/KbzKqahk+LLGaIcOTc6QXL4LmmW07B0znsLUCMNX41i/aa
3a6L7TfA9cSyOlV2VgPZ9HJy+4tmjuQKk1bDFvSnPoUe3pXkEVX9d6lUhjyp4vBu
spi5uPuzMxqewEyNkxld0l2ORbh4HuWhq1b5+NC1iY21mnEL1AWbYGobtQqIRbND
R1wv/QZsetbVZs/1Oyj/W4azlliuYmcV8xk8NLiJ4hNt423tNBRDj1XGgps2Frk7
AxfvOiKjzj69st0ZXGetx7YZHInSeY1EyTNjHyxztVGyBCZuwcD/pO4NhIfEtqJO
0tOendYoi3RNwnKO46GawSROhyKEn4wUGGS/739FgoavCZxukYAUEKWoyh+clJ6k
/WJYDCMLzMFr2fpBc4J68FFAFXao697HjCB49f9wmenpzcj3Jq+f3LiPy1ahDcLq
Guqf28UmPEppZsCRnynrDSgKelQ2kmtpfyK3KOjmgOWWhbGyydC0NKn7vzoeNT3q
CeJFlj4PoWMhIDJJl/IBpAF9xGHVcG4ZvyOCyZzdz7QapZRaHU/k3aGQplIcm2ow
6o8UeV2/h8yQPardjlg8TeFJ5sZKU4AX8NXgNC+7R8TyyHzF0TjgEEPqUdVtreXD
h99ptMz55MzQSAfZ/nZ4c+N9GJwDDqyy650QCGzJUqaAs4tcbdT6SdwrxBhg3sh2
Yg5I6YzoR6bbDeZS5WFpt4MGGECSaaelzuJ1RTk2+8M1u7rRwkUNMUsCaKk9ILEZ
3XgTpbCVgzAxKXqmq71OUxUWY7C8iIoUuAPiJVjZE4EQtuMUQGjbYh0WmJ1XB5+u
p8uP8gn/ElFQPUcQuxtBb+z32LUua3p/7Vm15jI22V1TnDj2hiQ1jLKMGyElkhO7
YX9InICppmxnUPUQ8jGU+mKWlZLpQSEZM3yan7geDev3Z4vHoH3o2QljtBd8ymkO
XEqbCFFqV+6645ZulzN/mYJxnb1mingYHo+mf7RrcfJ2abNlV1siST78YW7hDe8C
Vq/fM20UP166bOMBdp8lRNjtgN0WiCPAj4KruZTiJ73vcGpfQDroTLNUNysjUmt5
zK9myODpcVKhFMjySUPe7ZKKC38czuE5fz/NcWDE+dQBPA7jAXXezBTHcA57RsfK
PF48e1mdTGi8TddVL7BgP07DKoyhs0wi2GtAJhbHMNr38FTd8cBnT5qAbcjMGfuV
BP1vvvXlwfLCVU8LHxArK0/wProzsdZTKaciFW/GfIjFsxyW92gq88IVYpbM3UDq
6UawowsnGuC12CtMqn5zXI2KFujOema2difPAHtq8PAZRaTTMPlnXMyWLVuS58/H
koh9n7LLleRAtnRqjR2b+kvgdA3YIVmgtF3WxXEW4O1XghzsZXPcfsvExIaLBoqs
OPsHsxjvbqzcY+rrFyRRmSWR2RY4uffhmIw9GG8y0x49CwkT4Pta3Pn6Qw8zIjco
ZZz3xkpVz7LorP9AtkEN7GE4BfVvKCXK0M3FqaGahAdTX/qZ1rnCSk15DabFS0uc
3PJBVajoGypimQ5EniUstloSvqo4y4r2Hhg8LhFZkVLZ4XIOX8yoMzvnAA2Q0+04
WQ6SSJQfRMTx3PzVBSwy+22McqbzfCDeu75RJSGgC4NySYKua/8WdbneC8/6oAl8
7y8vtNY1JstoZG0632bkfOFOJZgoAN1fnbYMO8BObRgOUgFey+RDmJNRvjarhgTS
6FtmKM3msvftNzHlycA8FptkC1OXUaRx9d6n9b/kFXLvqXaACeef8kndcQje/Nfg
NVXxaVQdxgIu0OfmDN3SwuKhU+GWa1ZzK76mAbycKFrtQWHtXy47e//iUyDdsPRU
grGMOeRlnsbiJrcm/wKM31g9XMVPv27r5/Tm2o4FyQOxUgancHz8hN9IjEwV4Htb
3L+gzZZbqBuAixBFf6Ys2bBvICUWTWdbwAdY6xbUY4i92Bpq2oM7OQg7O0YC69rr
6FcJjieCFZxqhLgZH+bRcAfR6TzaLiFM3CsPXyWRpiaSNqD7LPXU0KurZnh33OwB
LQ49DOA5OAworlO7lGHmnYM6oByY6uPrrJeZZwjm39LUfJnDIqgcDVnxN0e2w+tJ
03jzCvl/FnFZ+Xv65ctNVxVLnp6EUipErfuPk9Usze1FXI+KPWN/jAk6cdGyzrY/
LH8SNDv8g/UyYgQM+23eQZZoSNSK/OAcVRv8bRqqmriSblRA6idr8o7tvhYIIVk/
a5QEWesJlSqJDv9Mh97CLr5rRie5LuN7XMtFgPZTBQOKVnoU1xqiYUI4luNKdeB5
pErC+Y9J/BWGe4uFFBUbXkbygWkQhn+DwpRL5tpRlvK97yhAO3Qy1h2ROtkKbZaY
yTlB+5k6CPCU6a9itNfT8mlA7ug+RgPmltD69yClqLIuCC9AEKXKc28HzaZN+vpC
FYbegBrUdZHuU8RgQSSGu9E/d6iu+JHjO+bbQTKCfJW6QxY4hU4pn+tOHXOwOI8P
Q+/PO3din0upB8hG//qFXBo8v/e9erE+//HqyJ+aEL9fDCWAv29ZgNeNZ/z/JRcq
cCO+Yr14uFoZuVybAv/9TZwGwTH9VglVTC+kp5ZeYSqZVIciKuAFf2fYvkKq5vn7
e6WtycyDvqQmQcQarKALcO97qyH0XdiksXxjlycDuZW9D4drLVvcNPWyimzb3Ufe
/TixgAzTkkv25oXIf1k9rVV139jiuQNMdYROFis+lZatr+MiuebQf9dB+aIQO15e
nGKutol26brCfuWI3pHGzr5aItHefo8tbTatO+OGgrj8evtEw2BNhx3n2AOK8yle
T8nBlqpHT31v+RX9oJTbSAxk00fBv4LonHlQUIRCj08O+CYne01aHxrc3a3dDMYL
01BE13I1/8QiTvM1lGhV7sv+gVzohl8aYrgHB7UrODaPmZyzZnzJps/S8kIhyu06
WJsK5WmItF0SV1jF7K2vJbv+VnlkJSPj8hTjBmdlJ7yKG41lg8NK2bOTy5ARjf+b
EwyZpOj3xQNHl5YAawd7HCDdOXtq3++UXE7MHf+bs+XrN/XMOuNBsorFA6lQD7v2
R2rGDxLZyCrUSOKKmhk1Y0UY6J6ITdWv2ewUrFCrt74yLDWwoca8G9+OyoBo0Tge
4O1hnF99iyth661YvmqvKRZ+Hu1Cqup7dhrX9aicH0AUPh7KThnZR8hSjL8hn0sg
6bk7jOZDn84K0Aft9whO0ZviFJea34QBBogro1Z1uwC224yyOkpuhRkxpHKUfoMM
OvM8/QlwcBGnaJ5C7r1NeDbcWDdq2qWX7u/NSPXPI1Kat34X8k5lY9BWTITlpB/+
Vfq3T/Keoc3VMUAuyRMyKf+yq85p2e5YylcphkP53MncXLu20kzVs4nLMvrfFcAl
e3St/ipY3Gs4AthziB7Nd8yU9rz96o3JKpPBbUtPX4lMZ8DHWCCU4TDS0ee+I3gW
riZE6e7xeaXxMIdEtr4zqnWMWCv1QtCQ3brH35XVVORUihzcdkBrj73/aMZlhbA2
8L2QTinFGFEWtFHiShEo0Yu67sh+WLOZ/D6LxDotuVW7Sdsm6VOwcQrT4F5UbtmI
TkC9kxFFcpkkAngGCYXBkorge0asuqwPE8KIFJv2lxlYqMmTR/5EtYCBAbLvW5WA
1T5KJpVHF0tbDmrXHU4fyTxgiji3FcwmEWA34MykeezFEwwM9a44e/837B7D3T+j
zqO5EJJ7HPbd6bkEFLffr3LX0VaZvhfKoKLL6Cy3eQleR1IIEUR2MOYZw7Gl8twy
5G9O1nwDQ45dAqjRuKMTfptHO55XKiivIIZIq/iMzDq36CR10SapY4tlocerYTxG
rumNzC5ty3BnuN00pHE/pJ+PQEXtAe/T1E9DMIKZ0UWDu25B+hZiiJr8xsmoVor6
q4ihYE9zar9pbRu2r11L0zEsgewPMnQtoJbAi664GbHuj2nYar8tLKXaxETH+QM5
w5ygsXtx4Y7xrW0x6VPgaSaBFWXwrLtoeHBuaflnxZCwf8z+wsRriywM8l9TVZd5
7geNEdrnIRyLrBtgSWfknWfeNWdHsWUoD0+KoCJ4AVzmxPCk44ePPfm7Ftq8Rv9d
SO+GPuKfFb/vOkEm2UKuWFYZxgpGN9wPn5yAd8XNrZfKDT51fA0oK/xwD83FTn7Q
hpzJwlClXRA6FDqIv2aREtypdTOdsICK/futURsbH8woal6XEMAPMs3/vBgmCY0b
o8CcYiiznPTTApRYifP0uxy++9hwFptBiRBnNgN7FMwhMpArYI9eovYytct72Vyf
mLklndn4IYJf/HHGSt+8xgiPfJVrQ+573qGt4zuQNg8F2Nt0B+6tgyXxf4ZVe0s8
pRFR2SgAllKaRVsCCbOQeoMU72qcpQhsmbAKihPwWaR3YmabBEVhRmLOdUXRcTXh
S8INPHqjMDfCOLv7dmUDR166GDEcI3Z4XPVPhDVYiQQsuKDYx+1f9igttrkWBVy7
G8oe+ptB3gaHJrmrO6qnivaqSxTNTNX4PKv4dZSon5Pa1KZ64iwwqMxe4OXGsPnB
asRNzNQM/gYVsKBf8HQdLdr1MWiynMmtsSqscsDkzb6KseW9d0KvKFROsSZCsSjC
JHl8BuGg4TwHlzdaMLsD7pWj3ChkZ54FLwhWXlXhfsK1mQTFks0si/HXDr4Zg/n8
LIT37+r0vKS3NAd1/QDs1SIoeC+KwYT9NIDBWieP3BpcGLrVpWPAUmFOXVgB1oQj
5LE6gIhELCgqYMID+rtbrFGskuDlsC//MyqkULkwp3z0iIvB+jTCKTspZvdJWIyU
2OZFn7Cfkhffod99T649bd89A0WWLkbxd4FxJZ5aMfMy3XgVibyZS8uL9ZnRtVlA
fcq3CF3YoV7J2wF3RJPth7p2IhK5BcNq878bCoLQkCirNk2ivFLoch7At/EPonT7
VHY1NLAbmdACOM1Aj+jZoKCuPLGybja+XpfC1RkRsBym5GP4YHb5OKChTVAwolzb
rhJd4rOgTmX5+pgBguIHznhm8OpUOEWvCTtGHKuC4q6IPsFhSndptBpQYX/pkWLu
Khq1HIJp8tlnuiDXCNL5T1qHy1gW6Ph1kRHEpuS6j7IgDQ6rsvnAGCLd6st+w6kt
eQZ0Eea3ys8SExWBPfhjdNX5B7tMnuBrzIsyp6HpXk1o78Mig6U7zBUDf1qXhel0
5KfSP7h7wRrSFFIJLSCuULvuaaIu/uqjy8WIrcVx9GGR+J1zPNkNlVhy7mH29g6V
jvmjKYPq4Sf8jXZkCC3Vm6Gbq1SrTDYex1GnYp28FKU=
`protect end_protected