`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 52128 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/59UwEX+aE7FohaWu0/8IpTj7mav863zUNIsgIH2BWb
Abd9opeuBjbGF/waQMI2vMJTwD1ie1YueHc3nSNpEh4OXp8P5ybZFY89uyGz3ztU
W1EsuUnchJoQgbHZ/sLbgtGRgsrAFn+ZoIeGN1d6RAF2wAESJmYP8zw+p00RvjZ5
pBGEHX7wooDexzkaqKS5G/Abg1I9DB+g7tix9utv581SxQU3v7LlTg+m6jJJPLud
FcM0zOJs0TQLJ+XnZZnyt9RxJNBEFP4cXb/vKzjYSAQ2MvZ1w4GXqTu3bK8uFlhn
e8amhIKmxlvK5iI86v91k902lxyr98AwXEuEZh3FTomIsW6A6ArdRgrzBd/MERVi
PhluWbZ9uNL4Bm6blt3lAWzhQy7vE67BfCfT6nIHndHnKyCjuhYR+awEnSBDffr8
b2sZz5EdNIqYfitMyHwNiIiuk4jlPBbMYm5ejPEjOsMXhCj+6dRZ+rtAyx9NVhLe
r9djxqsBwAcf7lNB3AY1CvojVkaJpRs9kd4p+8d2ICQn85SJY6N5LIEbvBAk6Uy4
YkMRyfVOCT6f9TU+vO6K4DXAG8FtGzwpMKaTHulQAOITdL+5fCWdbmIoZ5RVkf32
zaU2ggK3/WH4c+n8DbnY9QXtUkPWRdoXz+eX0tZozrMXCFqMmdmY/STmuYn/CjMY
x8dritNEHnJFXmuFX91FSKhIR3jse0rjpaMVRZP99o8tyRjOu1MfiEElh1U0fzqr
vakullAyzhbx0booB1APzuq3RCWo9+smrnaWoM3y/+YiiR9/YclDunz2bqdedvaE
Uij3QSk6mT4EoaPG1Dio7ygs7IFEfKrLGxlDcUeV4haAR0q9q4p6+APytPo3iGVq
IMW3C6ad0BQuI1qm+xBhwJmMVNPuTTLvYe6+ZvVuEQYHlgGtXhKNVx5wrWL8tdVB
FqNZcR/lMldN746+HTINGm6//+taDv2nVZdsHXSAzbBqf41lUE7UVQk9wI8CtJ5c
Fouwe24ADa0A8yq7IUq/O048hb5M6bT7hS5I2/wVW8Nw+5F3qUh5tk4ix5voWDtJ
n5oiuhCkl0PPAGn2bm4SZJGkBbqLcrYhJn6GG6fBFUQHEA+/sWN+ccMKEpx0+yvS
w9hvcBto7+wWRMlQuQvh3+yk1fZtsxaTVQrr3Xu6JcXg/aMv+NJfAM/Uz6vAEY9I
kUl6imqnQnMB1FSw/A9ZQGQsiCvtCvW8CuuFvx73T/KTtW3LIP4EKUqv1zI0zzIl
Re9Dedz0jHJ4nEBgaP/ofXCmLRkXM2tHKRd47NGOTQ/4fL3IEqB6jwxcFxitF84T
Xg/dX9HiLuDPubb7mvgkEwA6vYK0Ezh2Hreiea/rtrHzKog8fXs9NSAddIlxjkEi
258kCIYDhkGgxakEMKpceL3xTGvEpWxou5DA3EBo4+jCr11mFMElpp0cIihZIcSz
1XTrCTBWS5E7OM9VcCpAhcsoKVXai1nHAat9gynBHYT7y8YaNcNCcK9WgnIRWpS/
y84JMfD8H0y/86OzTZiX6GpuBBf8U9WngRvK6aqh2++aYTpJ1CS/qrF/PkF/FWhZ
YwNrGhYfByhtBbZfpXQyrEl4yhhQ+9i4pwWVLRXgUfc5HkTE1H/NkKDfRo0aToqh
QPiFQjZR5RNIxVTmkR5/FE+P3FUjNS9slhAOVb0m3rd1YbR+q/lAsxjRriA+501u
fAkJj9+eqqxhDyRlBc5w2TfhXV3Oy+1JT/OXe0xfois2ntKznG7kSxeHVR6NMnyx
ymKHYK3Sqc2A4vdn4vsflOaREgsRih+Zv7RJ6c9grIm0iIqcXVd4MXT4uegMC4W9
GR3i88xfJC8DItiKH+tBx4Srt8mxiWiE9vgbytOk0xfgazVGX9DxTzgDZIQXjl2R
mP0pzMkK3tUALPeL82fu4uIGYUvlkB//r4rJh1o7hr0dfsduaRqkbHsHlt2qCSJp
5wFNtaui1z2dgOsVFWZma9fxzgq+fp8tj6x+I4etI3lshaMdl4Il5UhbJKPUd4LZ
uF4H7Jay08ReZ2ogftI9PXapTnU7FpeE6YwtTc9GjpJxN1vRURfMpr8e5Yc8qNGJ
IID98CtBeasqcHHZ0umbG/l0VatSzcJAKURHndIk8eEEkbJ1rpveJ2N2/M7pz9pF
2KBvaI6T4rzO9lMozUDuLylYBccx2dHi2MCsJpBLrcBKyvr7oWxKNDekOrTOPBtc
X5cnaRNJDHfSaUw2P9KnzCIAJS3YDIOQTzCldv4LUZEcpaJPNpRepNi747zN5kBg
KwayIkzTAqY5knyRWskJ1r03/3zrpm1Xj+8n1qR499rxWoGtXFc2j9uZerbbYGmt
wDET31NHJd+SW+xFkbYfzjgSskJkRTy5eSZSFpEXzgOYDnxlsfK7/tMPocKsV1OM
ixbMgOh6mCxs3O7UCn8w0qc2T91YUNnQAvGYBejIGofnj3fwZ5W/PBBSc8HHO3A2
bWyFZlDfWRBOiNTyisp91GMgkDBsVuroXLClPYi+1ssdIM2PxBrV4iQaX7kFg7X6
IyJJ0S49T0pMJrg24z57JLBEACDQEos2WuaJ+/JCdI1603o7xSsGqBCFnXSD03I/
gW+mzDpGggziPxIGj1x+NpZVM4EWRwFO9taHrjp3LzTHHFOuQ6mL4Rz/pca5Kyp1
ewmDaT3CpMBZKxxlm1c/krH1k0hiEv1nE/T5jzQZwVb7QktQ6Gi+3lQiGE4Q9RTF
ZJu1q0TYIldamFg//5YRh8RQncApEbTANzJfXBKU6V5FXsvWEFt7kMukjbtgKGfS
NNJk9tMr7KNEeFMMSaSiZh+TVfx68guE5BN8KNwZHPUnhEkqdhn3bh7P0dZrIt52
DqHApPzAoM+5MZ5uoNA9lRxIwPpYEELH+MQ82rg0aVe7spvIGPZQrelCS+/+aFvb
4WohpN80Idj+X2Li1QNuEnVPu89K3IFOAURQA0BapQH9HtuG+k3Bge4v3ToaG70G
B4YodMBnC0Tu5jNccnXl+8nQIoi8/Z4w6J9o4x0RCTBBWtc6Xt8PJiaFQwdS+gZ4
uoLbfI/qHjwfiGWR8z5TPQQvJx+dXpsC6PwDm6JK1QF2ftf1B8bLxCnIh+fO7MBX
GvghISyyDoMMEbhFbjjsG0KI9P9MFAvkayqXqd14VC92PJFRuh2x8DDFzaMM3xOk
rK2yqp3CaPGwhmrel6TdHnsYsle204LOOZrvzaMKGrI3Apip2ya0eiI+VCUzqAki
ZPQ5b7NHTwSmhmjuEIwc2E2kmszBmil974H9AuWtEteUQd7DE29plUACoWbbqMZc
kdgSzP/ni1X7Xkl8OZ/0L7y+Br7bqBRWv8jJ+6Z44WreqKK7X3XYlzzyZQbgauqf
0ESR1iUc5SnyWqnR45jtA4zetHhm+SpzreciWxdAqCuSdi+xpfQILveZ8DyIRqle
c8swZuG2ba5v+7P80pnnlkjVT4OChFKqetXam6hdm9fqgL2dgwPpXaFZ7zqc8Xp0
a5jH/uvKFR9kyk8hCqsq8DK9/YbF5kbKalfjXSwBu66TXbc+9u3blpzZNeoHT03v
4vZS/fJkSBw+d+f6OD9Z+sncYD9pvEsEUwVAmXt3d5u0a+1IMA1hiTlLb/jPSk3l
gP4COIp/jsbScQPLiXmyUSepGj74tnHRWEBPmqpUrPiLRHu8ntr2EK5VKn8LMZfw
ziqiNzwizC9Q0gyF/a9T5YwL2PTrSh5wNsM+56BrOA/CrFJbP+RGjMMP4VPTZgLF
07N2gAivPEwxEeezHQJAteLyJNDbbStyw1DE9o9rgg+S3U63F9WQVVpoKbv1MDj6
pVfQfn53KrYDHc2p2A+5hekfuWzAWeFwvCI5gEqeAhHehv38wYwP43FlQpw3Cbvw
jnzDSJu12GMYLai0j6aGN50AvMEMYJOXN0zKNN/8lc1NCyw92JCPLv1okM15sd//
PdKUajmZuBrUT6eKgeRZzvKNatCQ17s7+op+wgUJmSxeE3p5l73qLYNLfEa+bosF
mMDbOX6kx0P/Vd0cqHaKGtBi31qTL50AWV+v1XnzjDljAPCdoBvK/g4ZpGKlQRFV
HgbhOXDyWUb0emKROZknELwRlwgmTwl6HE8YRBQUUPCNBv9YbNcU9YoGJQtbktcI
L4/1iV+BbBIJ/Z1IjVSePNrqBu2EB6PBy8X8+PQHqzvnAxcsUm+RAr5Zp2TEk0hd
Ps0QpTaTfvXMuGOqnWJx+aXhmfOxAttVGHEhEHQ9raeLCwN6pwTogPcQoNo5oGTp
7I7naqMu+WdFLBPiS++/axtYqDBErykjTH2q56k1vDh+uo8MMM2Ez0h5ooyXS8P6
V4paNrAfiI8lEwPXYH1xw+k3SC07TPSjw3MNvncO1oL+MfSwQwK7bb1sgzgZHhWI
Dxh/NrbXxntODpme/QjQW1CYRthM8ALT3tUXS8hB827nfthEWmiIR57cxw+p3IuE
1SdoTx6d4DelsY8KK5PDQ5YtExGHF2VvYgIDr/l0qmg0rBTA2RCmp6JT5OnC1ILl
pubYsQynIXg+UGJFL0hbxqcpohe+Lz10coxF//eipryEa6hMqpBxxDy7C0iERlwS
ebBfy5FAh8ydrMagit4EYDMgf3Ue5I0rVHfdB+ua8Mmkv6xOvibhhD+vZ9y9FVS7
epIZvxPc5rDBhKVmUNXsY+qlLNBQaOKpfFdxhUSYu2JTslSWNyIMcn63uzQTCi5r
GebvuX88EsRNCv5/zHTqPIzZIDLu16QBU/2Fi9VtMaZwArxVizxiTuihKGevkn+t
IbYcU3ErzPkh1cBvmlkRlkpWSduNaIeDX8AQbdj+/lZ7uc1HDbc/JwWl3vy/mrDY
NJgSNkjzI4sOaezUqoHlN5ZXd3UxHcHLfAprD7SfqzlovLZD1KwIs7DAxKN7dGUw
DqGltBM+tw+wFG/hT1OM81GS3U7a85E0H/3pkS07lLE3GTEU6J9PuHL1ow+jz03F
X8zL8eOd9EAuYFXAHBBHPBqLStV3w5ysLDsDkVCdW9o6BgLJG9YVumdcNAEkEfTx
UA5wC8h3HrVlorEuAofVbRSCzA4LeNAQ7GExaI3+9N+6ETEcalErXNvlWvrgb7a0
0t3mB7rodKV++Ky3BiUEKL/4cmmFH/K8SpevvcpeNgbfB/dVsbeGanbVUC3vODgk
5cg3tsJN11TvtAanR6Px8sVjpYeZvMYhB4JSDZgH7+O/AY3Wb0JlKD2JEcTL6Nlr
FuSoetuEE0nJ760QF8UXmrFiSG7o0b6F+3jW6J0aL2yESSjesIR0gHX0L3sEuqAM
AyixWk9QpcBB3yM0/VFK5dYGFr3uATQMZsPQvoHVKn2BIBnSC9jMB98F8hahp1+M
e7QIwrI/j73dIj3It32qHjdI68oT7XUcWgSiUjIvDo0Zeobc4c2/alvfguVMnRj7
guqS2lk+XdKtIDWmAGE/LJsf9EtZQIMgURPItPkKB2pJTP9z8ZwDoz+aiG5zg8yy
yszRuLBC+bjgfk4EasxBem8vilyNaPAxaCn/KoexsTUgdw8XLQJeCYyINkSIeInF
cuXei8bZZuTLKBW6lmX+OVHGbNdG2LNdHbYIM3fIZFo6MkXgSnL8B7G5JfZWtNHZ
/8ldoR8oB7lvap644urk9vUZzyNIPByMB92LkWxoMtzvZTaAw3Yyz1lkxNzCOL/N
ynGyLohxzjj+b0mp/nUrgc8Q9ZdKHRL8VTlaOGFOWqLUJ2+CZrdkEtpVXgBK5WP2
pZeyOxVHNFLflaThRcLI/Vf0JN/MfMEYkq+d7UrVECpJF4qfOUXjRzamqgVO9w0L
6c0FuC7KqHq5M27MSLE+3QM7s9iqLy9GX1S1In0EeZ4a9OWpDvCTPy1/eR5qBsO3
MhTlqi3tU0Cxbvnu3wtqRucDAtr/BmWhazh5uPxxi6f58nIeJUn1meiajqP6tLdQ
N3ZzvR58pgOoQtqzLzNzlloeYCbwOeQOPSOPQKjr2I4llqQwlyRBdBxRfvKQqTNq
zYEp9jFtzAGPDAbxqy3QZwgYfiNhQU2nE3/rlo8Ju2goJJonUNpLUB7znMFP7sFJ
cvXW5WpjYjw7EDsHfnxj0LUCM+M1IdrBZlvBcVjofBsvWe4ikPhlHbgpMEuem3rP
LvB+9Q8i7QRVv0LmVxDstU8sayz5MN3OXEs0avlg9Z1tWET74VD0OHjPpWDSrwmH
MO+16fg7wr/VMzlkI4K4s5QcyzJJPxtGCVph4Ga7yt0vDJhKdOloNwexy7veRSPA
KmPqQJC1IFgzY3XuVJASPCGoQUIQziY/9FuRI1umJwZhkSUD4XylLVRRupyLddEu
fRSGDLBCPZelqgao2hV7jXcdFUv7mvfQSrFjDIJNeemk87cRcbfdm6xEmWc1a5xu
w+PSkVsFC98MzvJa7r5vorllujI7VRxoQZsnH16gi5a/Gz2g8MRhYwRCUJj4TIiy
XR7OCOOA5H++P2VZzH+t4acVf6qU1YKcw7ZSdIwuwTHmLPM0LktT2NnyNnLjhye3
DIXPqaLS/kJSbR3Hj13RuKQNhgVVp9OvUOpuHdoHF1UmzwzukFww4u37n/fcrivG
zaUKCR/O5JCAq33JhsFKvKhoTITMHCE2VfQ595EojtmF+6D9qeS9Yot8xyWkRf8K
vdKC9XZlE5AU1417ePLUNMp04v7n+AzTUr2GDqDJN8ikY1yGEQSc4Xrbz3Y8llmi
Qy6npoiHZ5+RLSNzSaVUUR64TfMtqxJ86b4e57wDr7eFbQKW7hSS08gHWLeQd8X0
0E2eVCYA5CyUIqZaBAHT+yL+8ZPQeOdticbTXuQjFxm5Ctn7o45+RcuoH+e3+kNK
Tgyg64wLFCUEZMEa2lDQ7y7mWpnqHMX58R8fhiKenYm0Lr/cZRSzbptQK6Np8/q5
S/V97LuLALbb1hSx4RyF13G82LV+oDD5/SBWxcEfOzPFe6I4I5escbA7zXULu3ZH
CKVM5f/cWr7enbqpcImo1ZEMZJZ6/d42H/7Z3yQlOVJXtumDZqXHTAIe56jslmwI
04eTemuXyXI1ykuKdrdWfch1AyPiKRKtBsfGOgTGdsdIpIUjdHwBuUujMu9N9EZ8
IZNlO6t5TwHyrpN7ecS7fh6lFxTiPw+tTulrI/kcOIHShqeEpKgWazo/xlEukTbg
gUfjVxVn4plMk9X5w1MffSkVCUax2sA/ZFB7RF0bKil5CelolzLIita13aPGo4gX
lG9iZ0LadOcOgs05HM/iDgDGFNTdmPQs/fRN1qNnicMpreBK+SGXqXXj1vW+34HJ
M/7P+yJ7cPzyrenTi40tVxfUqWbO46zlxEUOdTuO0IeX91AFcgIG/qjQ3+uwe4N8
sYJM4yj4fdsThUudZ+vLKjNhTnG2+KUM2Un7tFEmPEapRP4YEBVE6B0t2xgoU90P
BM7oqvPRUE1aKtIWYHJKrGFMCh1PDRkUstseL529Y4QWSaxkP17kDrLtNb5v7c1U
jF/gX5Wx3FuUOoMUSnN6Mr9evRTLiQjoGrHYXFsXOyUs4u6lp1u3lcoQweTDcKva
Ax01nTCtbV37etgQ7q2nLg8MQH5JIuqk/d7s1A7bttNOKeGu5vK923LQXid8pvKe
F4yvinKUJAIGhWPy8/oq+LseBwJR8JvsG2X8lvlYg4YLU+WA4LXXNQRfOQ4/6lCq
lutuZkcSCLHpmZAC8BFndNOZf3FdqWq/eRBtATSOqCkimAPIykfF48lJkz4RgL2L
Rx9Vh0ssZoMeO/FuhMD0zwABlrF1Fal/I85XXJ5ZPrqt24zVgQxf5sPSn3bAS699
ujtunbBL3cy0Sg8US4k20QK72iQOVxjqYkL3jMMnhIsGBjE8XtcJkYprvYFDQVsz
CwSTUv7YrIM/DEy/DMbhiLJsc2KEpvZ1oGd8sUCsMPqsJ/opVph3K1TzDtEppM1O
7reXuv0X/5r2bYZzRNp6jvHVxn3rbpsXEPzdfA4RnByKhI2bCvm/bfCcmfyj6G2x
mgzJSYVVGUxz6ku6nlbgmFxMQ37TmJAiXC6h92t6i7/PpoopsJLv9POfpXC6EWie
AH5U41QJMj3q3XmDZBwT93awsmkj3buZF4XZG2PQtIko9kzkUit0wy+FkgGwZxtz
pQT3rqq4WtDJphZCPIgSBNCNNiR4UO4iKQwgMUVBAGWAA53dWYyZ1ADFZG9Zl3oJ
MglMw/CT658IYhOTi7I1Se/ynrB08yBGQWfI63HDSEDVO4tQCvZqdiSvZ+KnUlFj
IE9o5aSnAUYnNCbpLgSbJHNeGs7g2r+I281A4cRQSW0xiC2gduxyTfGQjL1y27DM
ExEX6DHoniQvfPmW5ZPnZNBMR73GEPv/sm9o5lRaedZ4R24BgHJq/Xis5HwIFOdd
+Z+wjkx85/qtW4WqC0KLDZFTQwZ0ROUugI6zKWwkOSBWUPgN4uxpiXxwejRgZZTW
PDSCaQj+LOPMI/qtSr4fzaMn2RTYkEj3r6exc9+zbw4FqU69mkTVO6t6hGBFcH6f
kh3vgV2JQNuVAClaS24gnzuoCdjdP7pJc/EjOQ9sJvgD0g+lp14of9dmRV/2jq7G
ZrDwX075nm74leo1SzJDfYpxDqWageSdKLr9iSfMTkIJkeV1D0wLg6okN8ILTPWQ
tExoB3MvbjUEYPHkNscmwIx3YoFbqNIaCSIe8m2tdEdv/wWEQu2PLViIwrMgymeT
+7SGpwf2xfKSjmGaNoL5BsUZ/myM4Z1idk64d6qKPI6c8xjlhLTWZiEP43XWGc3O
IKLtnQT1P2UokkRsHJA87ofWeRtdgy2gefq1xKIdzO64AO7jCSOO9BrJ/Sn/Crsl
GKJQReswc0Ctd53C6pdGw/UiaLgTVrVHsXqvJvUvV585EnFekciMP6lifREMi8YI
sPaxNafhtjSfPHxtTMoph6ZvXMuA84NluCR2DjQp24MwDaWpF1EOpAgRC79E1lic
XJn+SHCcThuy3iMgV4N56AHzVJqUmu/FYVc5PtBnDLkRNzJ1MySdRaHrvEUP+hMo
f5PLhTbOHGNGHxWL+4GeUVpk9KalZOBG4qEPm0OmGXxWIlqG/2InnkrB0BUiFHaD
6FVm7n/E/bfw2eHUWUP27bnLQNkirAZiEQPu1/KKeMHCNoWebqJKO0QrhWuv1pwW
bwt0OqyfaVcwidKjCwwqMQOORHKLh9Adm8A5pkHdP9rQ0Ym1cVYFk7XUiqvLHdON
xUyDzAZixAbq1p14x8AVabkz5tVT+awyDsqoFyvQKz9dGIfmM7UdsBoSywsTw/Kk
uhQWuv5nX7Pujab2GsJ4XEFvKWli0yCjRMLjywRh0bxAhpTYeblDdY3+pdrfNR4S
Jf7QS2AadGxXLv5tiB+4+KpmIBLc+YLyuC84Xkprg1T+qZy/g+ZGNb8DsK0/vV7h
bAegyRSsl4rkgkFKo2ga23Ych1cC2KHv3rSuFXYlUrIWxObnmRXT9YHExirKooVp
ytGOA9xrlaZQPZarhECaIRsqBsLXhwimd0Pb7YvtE4HOGfD6TIap1p/VCQiqGtO1
WTm/GIHSfu6uwEspkCACDNi6oHCsms5T9tRbCv/5UKhf9zFmbFf7doB/aMxf8l24
p0S9afuB8Xxk7IxEPg9c+HnPerA9BQSurA6v/CmiihCXTmZUQuD8FB+NMFR7vPmk
K7YeCr47hP2rYZFGMO8yX0TSseOr/DH/qgT/eBhnwlUK3yzkP6AYSbTcMJ4HvzX0
nvp+HeZ2YpKHeb8spQVUTCQaEE51ZmWO9ZzHLrs3Id/rmgYsldmPYQLA8zRgz+WT
yyKmkAL3ubJTJMOyH5R/fefTZfCrVrm8NUNp7YD/IAWkojPjDHbHkrYZVWBAsrxR
8VKXkvr/XPaPEa5RFjq/0gKmvdhDm3U0mUT2MYglY1E4GS4fbDAo8LFoCF/AImiP
DZbMk1a9mVMXc31Aotnry2wyhBU3DUn3NUjTDBJT9DQVNZSMMpZsUSyygVkM50vy
dVOBOyYycEoKoR/zC4NQggZo8VGpiSXlT/wqT6WHWaJ2WiJYctcsZeisU3yIeBds
ofDPL7mzjSrMhOzZ9djuLoMyojHV1saj6VyV/3gfDy/Ku0oTTb06Oa/J2L7DOCI3
FPZHf9xSZUicj6f7DBiNkpfrzbb8wdquZqzRViKz8wcWLdpu/Tyn02fVO4SyZe62
U0W15PLH5Cg+k8heOe3RSc3vp7pwsx8Rb07PPordAvSOzShCcNVhrt2SbXLBiyd2
ZQFIm6Q4U8qUsl/9ZY7Tdu37WNOqPff0pLBSAW4ATWMOSGjF1GH+hLE8KD2RMYPb
UGQYKKkYwPdpqgSC17OprL4x9yjF04wLjEAYVV/nBioRiMBxeRJCR+IvdCqIulU8
VYKRUlBxHF9hx5VmvEwYo+rRbL7GljzNpL8wGfKe6chQjsPCquH6gVvg0/IU6GPn
zBq0I2FjJuPfYlDnrBV8jj4j5RJFNZwqIBoul23XYQXNG27DkK7ljz8WsesWBkAe
ukaNbuua2jzlCJUjNawO+rG1W4Z2UOpHgd+cwDVojN3lvcQdMoy15T3hvG5EmxqX
lcGgDFIY8fzG5yl76jQAICcW19ZzfJ7FKPsSPLneXPCcGoCkCObrNd2b1rwfDsA7
rfCqpf2Dj44KGKWBI5HXUGf6tt/FWep9Cow9wVdfgf15o8zP9TXgNDmTZ3dLhFv1
F/gOQxfKnNbBaIYPa2KamTUWMSeihqiZcdk9/WP2TGUdnzm8PkXqjFHux23MMi4p
7XPNnWROZrhJ3OyV6YtOVlLHqe/MSraeDhbfG++hKX/MubNTiN9juIIMWGt4BcZg
oVC4vfj5CjZsdsX0kDbPCj7tsaKIKeRi7dgzV2S7dzlnEl0OWZPxhO/HH7USwPvp
Bz3jNu9PfY7mKRZoWDOHU42T8aHSI6N50g4HByeIB9eseY+jO29P972ro/i+v27Y
Ds1in68zC1YxBMCUMy1zu7lVGcAbJZ/39VjXRv3jXQxccXNTGbGpiKiH1AIioILY
BwsSkgGqSlrDuwcfOnj+W3/rTVB8Vb2x+rcliHSzs/wFm02u8kVLX1bIawOoBTcY
mZ9egKmMLbC5gi/6jEMfR/zowZqSRiKQregNPk8bmr5JRPZPwYzuJryB3ogHjaBy
7Ifg1Cb/+42oFH0GJ/bcQGN7ksRzj0awMCJkshayuLTc1syYDJLrLNbAvZfkS56T
CMoYHO1se6X8ULnWj+jIBZbiMu+E2UJvjvGUWcf5IdN7gJVuVN8vKu7cTSATaR97
LnMG7FkZ3/1woKMzqEfgxSjFtukDn4/aOWUlY23CgYdrxDeH8YYn3Ry/3EivT0fQ
b0iyI88bp/Gk/UWC71gzTRZxA2bUa7O1x9iFdWW3g7T/JHoFMcPHkubCUe80jOqJ
ui9+Wmiz5FNiDvtGvM7jWUVhU1e1lMiWhZhRjjSOyqjr8H/cYXr6w5cuUK2PNIc3
t7dozTX7vSWu+OgMWklqr98xG1tVDANmG4QnOd5sb+lDAHHKFskUzely7lcyjpel
G+XC+bUqFIeRDFBhTGfiyo6y5C1RY+sSyL20fy59/LWS8mCKxdme8PU5+vjDE/qv
6A1ke0APPff+yloAKB/fQulM5vgEwoPQ3LYlXQbVw0AVKEWD5ySVLPuJhA9Kffoq
gjUvjEGWOpUvAyMs5PNonwDDQOykqBxmU5X2ts1rZM+42Eis0Cqc+VMw+vAlO3y3
7zLFdkKiK4qgeWet3TBk8mFaF2PefJP4qBbMVv0uasY1ptofvudWzi7wV+s+P1bf
xT0mAvqvjAO6wkDIveXFXtRApYnvwu4WFerew/1d37WP6x9OX/WBI/cKMhzDagjJ
3GXoOhwibyqKWF86wZS7SgNdMcbEa8Pd6ZVR6cQyesV62kl7UBjsiICVCmJEIqSA
wH80NWxLfRKmMGtcFtPpvmInoxxK6clB+3hoEkl51p0A7Yt56ApH8EKtzuml+oFD
ITiMnQ8rQfPYWtk6jPT4mhkVaVVumirUPFrsgCIIolV5s9k+14d8Sxo4OaYAbclC
Pu9nXRtlR3ndOsAZ+mxwlSSUym+g6rJ3GpLzK3gG2tTrTu7rk4GeTDAunRNj2YzQ
42+HTmTBfB2/uXvBsoxG5PoQAcIBTwQuCTTpFQ6z9fqJZ+itmo3/8QEUtcSczDiR
mmKGIBMKwh1Fmn3UWvErgdL3eTX5g98n58ESsdWKAisPUlCIkoaIBO6+kc/QfloO
J34FHTn1W2LyChPNGmV2B+Hn/iLhf+NRcWrWRsMANtTdstDxjWMDSbf+zAZ3ZvjF
aCqlGK/lpZY6kFl0Y8tP8lpdYf3tfr3MPlbDsEWe+03HQz6uPaLwQRFxxr/Hc+c2
rueMpo1PV1/xwS5G4kjrAz4UGa+v7GAkZ8lkq3G1nGdLnWjCDtVkrLwFEgg/CHNV
5DXRmL3/Zz+JbiqjvBf/K4ATupKq4bbf0ecVKWGzAAhGlbGk5SSejPRm9o8RJZiy
cbOicFpyT/NripaAfOKuzdnwKp4P9KBzmAGNANpSpyl10cG+oAAtT73xUQMBiBKw
FPpW3D5OjyYpXyJkQa/HQuTrWHi5IxyKTE1ccq+YIV47ouzCvrzTYsBcWYi8avAV
F2ZFOCKeLXxJ85kFUZnQ6odYBQ9B1Q+QvUY5eHNpqmrhUQ40zLhIhLIX9ZMOcknv
YZKNTLOeh+iOXx3GVCKo+HIdh/zkw3/naNU9BdkCbaxRJVZRTPniFkB+6sE1TeLg
UlyPJOvthWXzsE9pspz2pGkAQec6fsoEif1ZHsPPAflR8KHidbO4ybPrht3tyhU9
eXrqtlz351jdjYu4eYWtsImYzGR9QoKjhhK2e5QAT7RC/o2VDEtiixAZFUCel4Yg
m/SbIsefuuDT3eF41QZMG5Mc7szcnqFHP8iRSjPvxTAHdOqOiNysV9h614zy94fJ
EpH1dcx8g7+Py6JMegE5Anbd3UAcayTd7SJsc/AqoGMsrrltm8+iVdQpYu+ukacP
p3RL+EdJezOBMe1uJp5z5myWlAeQ742I6UNmlsj2gcNte0ePUxlgBZ3b0UEq6Nhc
jozFp4xdEPkDBdjxRZknxJ8d5tg1wt51a9u7sm03obDwuvGP9dhqCpi3JLTjdBlj
S1yDggfpKU3NXTgJehnxdk5G7vGhbHFyDYgvRot5sUXyOOLFGgnNqEcw8d6j1FV7
XJuLTdTydGLuDSK39n20LVViC+fH3zCeeu/bnyZRCvKrjSZtu4SpoiHBbvzyp030
vvFt0iIo3lCiI+sbDqjLrsjWBg6gBCihOR6fgrl494ZtSdFBXVhiyTVwr76854gE
EkC/LV3L7WdbVrn6usFv5WNL92X3kVb8FZBR0eqKhiOCtV9ZTPJtJ3bxI15TU1+9
7g+kR4AtzlRBBw/R9/XxyLseyvPHyCx776tPBXtZUZShg6zOfqN9XYdOaxsjQt0P
ym40gfu5AtdQA2v5RtvqMQy551yog5nBEym2sU0j7MGtfBIKMRz4DoubeJ6Ew4hR
IpZF9bQMBlgDpiD7W1N5rKtwraHsm5UgeboAG5ozzFa5Zbcs9xMicWXXD9gWepp0
3lMVjdaXpKikRAJVGWj3Pei1Z/7HTRWqH1IoqBq9Co3x3ewllL8KPnlvpVl5B8MD
dckgwWRpMOUtn+XeCfnlFBRYcRT8XqNF5jYmaQch5mXCQpqdzc7xBqICZOM0+8qh
+FByN7dnAp2CE56pGyOruBWr++mcUOR2vvVdSCWUg2guxT2v18keIGaBRyAE25EG
w9f8yHDsUeXtN3c3cDEtVMQI03Mw3klxHjN5WC6dEFzblr8bfqcud0fJxTH6ZIiS
FE1WsM8sMysTnYqoPZIrs7EjKOBXRftgUnC+cCTBehHsepx8HllGaszsIBvj39kV
s4RmtYxkcEFbzypDU5pphuF/WXBYgwhDIhoi+2sVQGKG+hTAhILYZrCfSPPiVBIl
cD/nTxutBv/UHC80ZRdUtedCI2kdcecw2jkjLrBzjxCXWhrf9nfHkoGtKba/rxtA
vt9vLx/UFiSmYKuPDwsq1p2ph5546K0G3/hXMcSWVpQI4zjdF3kho3VjZJqDqeir
maoHnzqV4d+Wxbn+/Y+6w4ex47jXQAbQBntrxPFu/YvgV8LEJ7I1ADVKUIMGiKfQ
KXvJ8HBOif+eMHxIRJLczCbJpnFlFSSKwaa+Ye2Oc+YJR1hzAaTg/QKUptWcC8Sk
mx+m7la3FwdEwK0wxZTj+aPqf0pqK+T1m2ncgaFlkL/w9/icVAyVoJtwmQePmiKe
RVaNmzs5zw319I/xTY3dToOsqtwfynep2in6TcoYpBYbGrgdn2dX+2g2eGq7qZkB
BQsyV3pHWboE62GhI6Z7nWfdbB3L2Po0x4k5NSxfsPepJYqshmDCy0fP/McY+RON
qU+agVmdw8rhovoyKaDb4LzXXrcSeFOAf0rYr/VpdFPUchONHcHH7JUOogsj4n6/
RuPDDhvW6aR9sXxE5or7O3TGwfk8Eqc4Aw24Nn7leGoN3YYTtMMjb2HTDb1syZpL
JH8X3s+AaySrsR79gmdbAYcKJDtQJURDG3wNee7gfNnDBgRuAMB96MdJKW8NSQa1
syMtrNtAdMjctgB+KvVOImWLyWofxeByS1Ff2UqJI/fS7+G5QF56t3kF3xbgua9K
3Cm5KX0t1GwAiOmj0bk5tm6VCYluXYX5C06Fpqz2YMGvRyAXiaNxeOZTbEYP1j4T
VBEXr2NzRfBFyzu4Q8nimfsxoaaAxdh8QyhJFQkCyJ/q33pR4kpw9sYCLLkTfS0L
ms2LJDx+OdjhDay8HT6x5SZ05frPTHuFebxu0A6KCH4morECx14Q+Tgh2I7vXM8g
l9emCuH4OsoJnRaJS5VACg4kIsCKaMcCHE8l05uLzgBgP9mmXols9uH470FwUX6S
fQCBmJNKh+r8BNEacVVHYwFhbysEbIl/qF5bVNTXa2afqZbcVT0kuqunAA1cVafa
5mFbF1gOcalw//xjcG22bGsdpvZaISxaQznEiSOGYvCOPvQbWS/xb81Jd6qROKVT
/YSmTR+wBE9Em59vGiS12fcw98DXGZg5rX3c3x3bBTVKbEQKIiH2BPYXYMmsxQq9
6LpAJU3Ut27hnvLS8fpbdOjYViYn94ZnximCIwqmtwv/greYvvGIJu8/EbOlFOtc
NdxdoK27FWs/XRd35HMVXnYhSWMqeJasE5pHjCwiJprShBIli4bPSOBxg4+J221q
kAh1xk+ueDpnHIjBZuVL+mntrj25yetyNSV9XUGiu7hIwrLp62uC5cM76dFFFiki
NgKcwbvF3e8hcgUBpdg1mUuJIdJjL3EQQ0AAzFwx8bl53ALP8BWjupksxBUwz49U
MqNqa9XYy+TRC2KmnGoKcDjjx+vlwFCrZgrtzCwL/+El7hd43hG6CmlpZJeLhEa+
10t8ZzN7pJiFKfM92wpDALq+D+Opa+I/Z9LqviQFKC5UMzCemM3ro8VaCyELVrhY
g3Vv/lw7SzALhivAInEa4Frn84WQraSwrXRDHpT5KZc8tY3pFq+Ry1F9ukWY6zPx
htHnFV3VPLG/2rsWGmgpitXMfPi+nsWEH4m95stExYus8CwDjtB3zlwMKnKCJstf
DilgGBwcu4sPCNCK/inY95+qls088wAW1YMCHCtjmm6asq9pxIUZKF90YOeRcIEC
EyqC6sttA7WLnON/iPuGEFud5Ua8UrAHv3YuJfdePPROm2bJ+NvV0wVw3GZjsZru
EQpQ0EbbjLv9gQYU99AV19XzkTaB7eI64d47jLNcukF5btM2KHgk8vVZsipVVWi3
3B0FSgzLE1MOOg2yM3KTl8XS12B3KIpub3rfImhmGKozhiAMnC4OBn8DgOlf1LaO
OO2e8//BPP38LhHVY7TbbbNEwT+J/qnyJoeI+qznZB2Bh1ydlsDzP+qMBYRoRnEk
buVsMuxzdrbnlC2jfgoauOt/JvWT3PJdgDQFbg6CKI30hdTV1G3+0qovimBp3nR7
dw0GmoGKSj3aNlgYFfF/6JlbOoblfm40+z9yEZMTFOvPSOABgaoT+WBm20JmY/6h
RQHkW4+pt9fOSyHzt+yxIZjk74k7KQtebzQ3qO3ZkYSISX957KrCGoHNcqhWg4VD
VFQC/zMgEKYoC+MuSo61lxCAcAmypxXNBd3nydHqDmvKkSnGnzJDPu70ZVwAs3g+
6MJdSCS5zgHF2fN8eHy2rdxbF4ZD1U5OJNF1urQk3hxILHG/5Fy2241sXB3/4iCn
BSZQVak3xZbt7kP51q0rViK9E81hLIHLpPlFD1vm6lGStbtfglnddcHAsG49tsXy
VD+Rgex6hTsDfpOjCHE/WpADIdGVpqK77qX+jfS9Me41z/vE8elp+ilsoa8xXA72
hyxLmz9KaEG0t1uCFxjGFWSxGUYJAOxrrFBYEUxjxp7GFO47yxHpGtsADT+tVPhy
0DFX+MEmTVzlZcREU5c5XiDujfIMZ09Mf5y1pqB1w8zYoBLLQuAv/goe9cr3Y18J
GN9g+GGZJtY/VzME25uMom+ZybMKrQOvAY/4MJwWP7IEY2sQqr44TaihHSiAziXy
97YecyNGAIsGbZAmhdvyXAUmGLiQ1RTtWs+M3qoiU9yRx67zOJsLUwU2IIYkplBH
k2xzjQerkd2s5ogKEASckbp3GaPSAKiRN/0kxWZtVeyPwxjCF2TQp4LarSTaEmI0
z3MsfWszTCXGm21VC/oMSnLzc/87WA1A965tUFP4rVgCYudqTLvcMYhKwU4byFbr
BDRc0bz8MQ1L9hOT/BS4Bc6hyV+XucbxOFAvL4EqpETMaZ+UTOZQ11nVi2xsOtYn
pMU5806Uq3rg33BvOzdNQYKEVKMMbXOl8MqbxY6xPATAnfLUFDlRRd+0Zb2osu6f
y6t6MW0xegs4/fZ6+URh9+96yD+zTuUk+BjeK+09GBCtwaEsiK5iLdYN9rKxHN4U
mvSilTtnbfvnu3kcB5Y7s9/T8zUIZUUv26fSx+NPlOLWhlY972ISOmSK1xq3Aqn6
+m+fWWTuzveBYRxnZlRc4SP+FbGqqix9RNG+dZu8A0j7Q81NTDigjoTrgGb9qFEB
RdoWEuG7pdAmqYLZsQqjFwlzILD0W1i3yGGbY/7Rd/M+3hmtfSiE4jK8f6eELn03
3Wl5URAb5MizD47jTmxX1XzY2H/flmQqI1+6oBhEp6Jl3VbtI1Duyo7iUCrkli9Y
XSRSIHj+0Tftx+t1edbGZrclvdc/IVmkmWz6so6CJCpYeaaN75ci47ulgnC8HyYc
ecK70CNsLVKhsUESD+okw11gD10zrH4XUWWRqUMy3LkHbW7nNkLTfw0oStlIfPJT
Vaz+7/5gsb8ggUbin3QRY1pVLjVa4Wu3GrozDdFdWIwJ5J5nR07alm5yZh+g2tDJ
ZiZruRg2i9F7KTCrJuU7rUAcsNF0io8LVMEm6b6hC64w6hUpRxeD4TnIPvxZB2sZ
RDCsK+P+PQa/WKtrS6UTXLSc6ysc/hfBgidMS0vhAmAXmK0bK8A/lIUWRSWIM6wq
dhsRl1+vO88X8LD7UrWevNUcX+fV9DAzvDD68u9b7Zve2z5yUOb+xnZfUt2eso9m
JvLx0PjTlHWpxVFCzK0kStNGxH1y1qQHRs7w86K7MRjl25aFONE7TyI77yjXHhd2
RugNFz2RMxs41smBTHLaF8bcZYQnOcZJCkQC1ns/0Fc5jIUhCfQIwJejw7PoHxzM
yw3rNGTgDePx0+wpFOTqZHMsRL2RKyM3pwNiJc8+A/90glwKQazXdkNoWIL2Y25T
ujpcO7Qa+pbYqrA7mcavDNcmKu72JtQj5UuKpZUbn9vx2fKfAgVnVDoENvEDIR/R
FfrvgUhZ7UaP1fjMD8Jf3onVQhlbXj1sT/1SGSAYdbNZTHyBPDjWVeKn7MhFv7Uc
cNMWHkIVwN+0uPu9xoDHpzsFs+W4IY/2O/NQUCj9HQvaZ6G9aADETDTr7lcES1ft
olt19MJBZUtnRApYHzkqWK9g3j16QkXDgnRotiYBkiHzTYRcsKfolz5tZVK+Pb8X
k+E44BhGeRfDWx2jnDdS12IiivMUNBBIWfQzKYCc6iAVLgUUWyvRkUSs2ZTZV1EP
fJmW938ocWYNQ6zAIClni5I1vy+BZY7Vst2PslbGenDIJubnjLnvxrdRZ5acwYnE
mOqCaPPVowYQPQ0VpkwkP3mme+LPeyOWC9oCU0KGkpCY8VlT2JE10C9VchBBSWvx
2Cx1oS4Xp+0eV3WLL0qwtoVdCE23JPuAQCxD2j3yTstgKO8SewVQ1RT/WSur6tSe
dKjWa7z4MJ5CiFPEtTqphnl8fLh6ejF9phgtt7f+u6bj0uSo9K6LPmhsCvLdZFDO
+wgsybzVUw/sLY5UCc6wDeqLEJtvCUTrzwabR9ZIvYqhVEkiQYYpScvCUWN0XOD9
6ZhxeKK4C28T9+/7+sFSF2rkzAOTFWsGEWGHmPwjwa7GD/XHKwMwb3u88wpRu0YZ
+NIZQJI//eK+jXy05oZgR3ag02fIJ15WaN6S6OYOS4ifbiWtJE6ly6aPh3GeBq0m
umRTaAa0IYenTpoSaAGEFkxHm5xJWkwVPRbvOlsGa/LA4QCyaHx6c/8W4/1mieU5
IFbOHen4jEixkkD2C4ecOTen5dvVLmi1vxlWi1/43awhtuf/tVvUY351slA0PeK3
S5goqlWkJqZ2mVjFtstmtMs4k2gZHINQMqrcveaNXhCHOv5Q4in90YfI9J/STkvf
OMPrDGvDD8Z9IZGTuDxAscMaIPodnLKHmZ0guWwzkvD+2BdVX+0xuWDVhXg4YLEB
/quypiHwU7bKs0W+ephy1VGPLFNklfNdqjB8F0Wt2tKvTUQL1nlxa1c49/BFVPSJ
3L6FFpTDM9deSJjRgD3f1mdGRNR7bc0uKNYLk/wzswzO8FPLagEnI/fYIdrz/adT
XwdtubW/f6hrceI0/2DX4JSnF8Ogx7mkn1hynv5BS2oC0c7XF6araOq8hg/jo6bP
cKU4ku2Q2xdGvc5FBSz1Wtt1yXzTZMlvHwDvrY3rwrMSeAT3kfj2+Z8Du2HRFUJw
SI6jW+oF9Io8PkX/ONXBXuErMDWeiyS3iP1QkVBGGmovk3wgF+BhAKT/8ociN2Vu
P53fN0KOwJxLBPDFbrfPjK3hjD6RrX5SGCoCZePdTSSo7CTpSgBcB3ZSMm/pX2HV
Kk8T6FF4Kn+DzqIKByeueS8Vkcv0awVU7v9R/E7OCdAitaJ8zMneoSPWzNhwxwRr
5LYK22v8AW7lxu/NKDLuJfFGYm24cl7kF9f61mBcY/LPqLkYWBWUSOnb1jTqBpW0
JLsjped3yWzvxy30TE52Vi968Ri3/yHJdQ6A45x72YatKOdQkCLgo3gDuP7C+aqV
Puj+Q4jvijK58GmTBrOl4oEFT8Zt48rvAERDSVUnXwke6TE+OW6dakS6P6oVWhNA
e2rIVN3Xbjq53shaddX04ZuGNANy1iwra71/RT+0G5SfrdS5N0mzi7xslpXChW2z
NyS/MLd0y8oScmwYCmu8eJHleOp0JNyyoZ8mJSszogXwQCTjFJPe7ykRat/IW2lm
I1FgpeMWi6YeUXhsI2c8mXYmwYqd+08xW8Ez/NuNpAxK3OvrHL1INe2RzhygovAB
xjtdoOc7bDozKueTcHNnxFSJPDcWcJbt/M4f/7UPifDLSgwJwXyu6wFSwjlCgf/w
ii2x+VSa7DKJODbFZYa3/LnLIUm6H+mHoqlg3Xnj4KDunN03qxSwu9Pos9aPAhh7
dniDMYSgPoPPVOsv2ziop2Fd4pqpYiNeCktfZ1EYsaprzrD2Q4RwA3mqzOVUF26X
kMtILZ/C/m5/7Bf/jSPBdQYvbtj90nO16beJ1B8Sn4o6Dz6ZbNG8NILnoiQBV0RO
m3WTjtNXjPiYrC4fFyzYNOj0SxVMXHsMe6lTqKp8i0sM6MOcGtph+MqVcAdmIIM6
tIFtJjpgspQkHBFRGigqEFVI5Rh4lvWrR/3bH5VdfS6Z9JQGux+7d7hz25MuiAh8
7vNmLz9DP3jyFLDN7qBepLX/E9NIfFakKInA7Cva52xD/kYiCo5XUsO4j33ICUI1
oS1JfKNSRi4XP36aD9hW8RhRdoIStOUgU4RmP+iyX3hHTxo+eP+8a78St0w1TcBl
FzAIW40fQlr+GUo59TreCWx5YwZd7KneYJr52qL06xFMeiGCCQe8/ICSju8aLXgR
MtgI3drO9iajkIwR488cMU/dUsVZnGfI5Lb/IW0IyFB267aWvLWXLwpYIuWafBw6
AmSHZOYbm+ICO++MJSB9memA7UHuLIFNGIeBQYKRusQZF/v8mPAu4HbohvOi1J5W
+/HmnZvub+beEwwJIwnNQjf1VtEXRe5xRXrUBzC5Qbtz9HKQ+V8X5wEtGZn4Gw1x
jWTL3qBMmefaK5FBAd7elHZsJjY1rh6PxBMTnFtpVR0dohCvMB7Z2DEQ//N1ao5p
QdzaFlEtbvu6Q5G+0iBe1mvYKXWODu4FS9yDW4w/zwjvEO8EwaRaGKh97sI+N+kh
JJaVY7Fdg4c5I+ESGubk5Ahi1hVpkkVPl3hoFhq/GSgxpklO6NWlCeWNWr2dlSCu
3rfla7WxBhr1re/hTGqXRD2IhV0LBuiDBilcoCmXuwIILspXt3EGMwwEFStuJOzD
gl/kNmb6lkHWSdc/UC7Tw+lq7iwzTLBaaUXHbil+dvTMl/KGyh3KOjHeMLpQnxLc
Gd4xN+ZLVpTZi3FG+DPlTJquQeT1NyxqmHRDdYLjsVzkGJ3NzEEFmwKY1JU0u2xj
TPGGFKHA7Vm/TVNak1fAXMzCv1TM5kfM/YX2VER8HJ+9TQf/D9pL57k1+zi54uQc
ws8WO5P62r6M3gA9DGUfV1N1HbB4v4igna/xnW7dHu8mwhJYzOiXZoyrDVlfRai/
7dvHl3NUk2r1eEeVzayvPB9ge/HldJWXYZDU9WnznWFJBomUE/OB4ZdK9SABWYzE
Z0Y1mNZFrG5jJhXkGJTYlRiKGlMVmc41rG/Hed8QYLvl2KqAonsIqJTf3svUjuQI
XhOsVXqRbJ2OKPsvYxK+x+cD7csYTSUwHhvMC1/Xyj2dfw9jSZQyijWB2EYhqCnK
fK7VWwdZdEu5+fWsOq5y5fokviMZq61pMLhrld6Oe46zIhTh+3YCxIS++eK3y3Q1
2IdV5VEStOlOFXggwDzuAH3OoLYl4yme1kdM/cJ/ONUA6XhaQ1gw2yB60cr/U+/g
8mKHgy7L5wW6xi05FZAO+Q/4AGZ7m8tJIUw2mPUNYOm9I2nCYRiOzt5tY14Fk5xr
mgWY+lzZ/EAlqL/ehMLjoZWPfPrcdWbTvnBFNtzK94+oxyYNNk4GBeJntv5xtCNt
XlAj1VX112bvWVnYxihWXOu+nkPmWwmXfMY+AloNAanZeFWcOTY2FFKLaR0HHDhw
bu67y62uu4BBiwCvrGRovs2eh4Y3I14XFhp8itw4ierN6VjlSqHxCBASP43Or0OO
9UqSyJxlyQn8sLzf3nplvwsgN/YAXc41G5p3y8z1S9YtAfqx4m4XFkzEJzAd7jwR
dXNaIVyfV4Hx2iR98xLkeKSvKBz4xQVPIqMOcQjriqEUsIjPJjK+4ETzLDU8L7BN
H2IgpINRK5Y93xIoIuyHWZppYVCEkaZLho4+EsysyVlBsiGohhQcdWyi0wVQAQwX
E2V8b75wDKLq7cfpUEiQeOipVdu2zfWG7HMG+KGClcwpRcl9vErj7Uwk6jg79DQ2
NrcptpZ3YT56hqSP4IGLJPPjsUKc0XEwkr9QIdD00W7WXavjAqCEopJUWqd8qcme
ZpeYVLfoTMMEJj6dgyDBfyoM7eSjGjRq614Zn/4kShWiwxEOd676f2DNCnklYezW
1K95Abf9OCBvy+Q9DRDyjCoCfL+ptCjWisBm6nhvhSqgTzoD2hbhysD6pXaPi17U
ENSws4PcAz8326DzL/8pmNxhSa8lDNbW4AzGiGsoDEcyZLzVbSTQWS0QKzXSf6Jr
1xrrmfyc/0c0Q1afOLaOZDjXJlTlwdqfZs7dx5M3s0qx7aWZ19PmYvymH5bAnU3g
54WGSs6n1kBgDxCEVIOZQ5Jmqx/d0Z876R/ho/0gdxPXWtOp73dwymryAqLsZ64g
6Yty1TTynmENbN1Mep6IQwXPPJhljCLQ8QAVL0RcYLXQ8WA1c0ZVBAdeUCm5KXjy
RfbvmqN1muVFaYDX5uDOPjF3PsiCpnFjvSx1JiYpo4TYcJXzm/RXV3/TZ9Z7ZxQK
0+xy6389DYQ2prNOPwhRUOZUMw8IlBeraO2qgzK9DuDRsZJDmDtAVQvdxSPkslfO
ink75uOC3ABndja4qMYYJRwyxtpAsuWAGjNo5EnACd0FnF/n3xhPDIgzWiliILRt
CR3U6axLtD4HluXa7OzeXUBbsLWhlUfFaCk8u0+zzoPo0XhsrpaIqTcOY6z4GcVm
PVHDnBzbavGgizpWee75j5X6Qq6AzBeN38gWcSiJRWKbQkF9R9H1PdF9ZF6HjeG3
8RgYeqKSDiXJ15IyMLIv/7vg2+oyjVPkXtDA/y0xHAXO2BhYaKmd0Y54hu+RHkcJ
Syq+zUnR7dGTkQqFeBPOUFtO7L0ZRp/TYh5Hwx8VdWGp3nQ71j1IT5xMuYUIZGH1
ew+uBJb1U3m89zHSf7VodBkbFvm6NRr9wN/hgA9efjfbKGUaAhSKi/1Lh85G31Fe
4y+CNHI7jq6RNKuJ/TT7sbHVIriBueld1oj4e6P29YZ+5ML6YB4DMxaLE1+Yx97q
8nWUb8WIv+fwfAAoaHbbDtoTHna3f3fTHzwKy2R4jb1+G+20Vsr2Yq0+ajbwH58L
QxKd1L/nXOqtGIohoVjRzBEVyF6szhZWl/j4vxo8UwKxR8Gx17ilEMx8/vdkojVi
u2NZtY+TVs1YxmRN+28npOw1/rVXh0yHt6ZZ9m3hPfHlGeqd+7AURXtGPfEjPwzm
6qaptuLK/fz0vUbS2rJ9ZSCfFg81CE2Bnx96KxTfvbFB7dSLSx9ADmdSjBQuGThz
8IzQL1K7XxIXal9u3exJxJDSscmGcu7klAZZq6/miqVUeYf11BdNKhmGCyBjW3pu
bWEwF9irnyDWSyoXRBAx9dlgpePx2Gxc2kFjfinQ12U4DhxiZP4P2t1a0y5MZcvu
p1gw9Byvx1iA1QY4WkO+O7DdMijS9Lmf6W6zZ0faWU0KsHmdGh3tym8aAYxeOoWW
BezSF1OaY/pKG3rBvj+R+zMA9Vp4BQD+M5rMyNxrPWWPraNB2GJpHcVYTJg98uok
QUZmmVZIWQeA/aOSdMeQTWwHpUGa3n1LH4UrtxUpvyX49fHIQYPDEwZlKOCay9Fk
kxO1NTjv6UP0YN/i+fKpFagorh/zQyTrQGoBt4f/RPHweTcRREPvnA2rgA5Wnk95
cLRtA+rs7wcIo+zxHiL5O7VfCOoXc+9L9pgXmPgErGr5QDop98w9gcW0ssFWpR2r
KlclDntjzFASG10HtzqZ67+PsHPDqidwQM8kBUZuxJ6Q9z2157iEXAf+Aw3tNkSa
HqwCld8T81+fAj+sFQi3CEg1Z6MHbErlF9RP7jfQagDVdP3vd3LMbT9p75o44/Uo
vEY77lA4wOHfN+pIWI1WhVMWkRgm1kviqSzWkRygpv+qPdEoDe6+UxjEnm6aAJVu
7nlA4WCCcvlkvZFCWpJtUJ67TXaRtgvDyvWWTHxaZAOfFPAIDQYgiNvJZjn1Vf+k
xrcq5xdMRxLy6YV6Z0s0gZOdrXjh6tM4ojdjb+ZZ2viNVYM83rWq765gCRvGLwMx
XLg6wQmeMFqGcqkyWOujqBIb5aSyJwzWfWVTDLSwBa3sz6ZHkUrUHRF7GxnDG4iH
mRoIL4edAIdR/vfdglCZVzX2eqlGIh2kT/ojLgUWj6TKQwGp5Z+U9gt56OQ4n/HS
AbTBEMwfbQDdxDRbg+iR3IkgRVBL83rOtHeMAJeKp5jvC8YKWa6UWlHQkV91JpIT
HbFyUiovgJc2LLBmVTOCL96MWefcpfIvRN7FvbLXUJVKLAyMIHddstWkTikliHmu
czLMAUXEtyKjEJOe/iywOrWskoPS5DvrCgmoEEeJSFxim/uEo+afNRBJrki3Ovs6
yQt/D+XahJ+M2cb2Z5uL882kvEYhGHG/UcS3MiNwCLVuo0J3D/cqx4s2AqHUIuzs
f218UchilFjzLpUmCvoiC9D/bdQxd3Q3lT77BbAKU1hx3m97oc7KqCxKH58MYFVu
wvQeBlyyEM9r0BPS+9K4/6neJibfIJ9LxKjbq3RIk9tVu3Rl9NN174fsoQLn7H5T
T6xeyYvrpJiVpEziBh0d9srisVyRFg/N9fY8NlziY9rR4/4MOLwd2HlH1bapXKjr
114xA86sfH76SxQ0ynAL4oCr1k5nCVhPs1/FXX7kfjFyMsGYsaMxWiIiLZBSHAQb
sq/N2K/Mmf//uoIya71GbnpeROOtKzwQGSzmYRKBBAQTmewlrK57NTagbm+fZv0W
OvR9cUGQ9jOEfrTLP1JAoDZXmfd7NIXMirt6hPDM0l98Jq89QuOPjbhOq6d2tubz
7urDwajDv9RN5WikzrUebOcHL+UBUwY/5LOBInVnYBlGE3s3TIQpuX2KpdA+1TBZ
USM0Mk1+rbq36/TcGovG/glPQPcWsHRrPmErchL3lUST9GapVtPqi/AJKuZiUfP7
Ymzlf/9u540Ge3zbusHaADcyKNqTKrvM12/MiO6IFKUb78EQYf5UGUKRBz2t5Kw+
JEBI+InMvOpiS0UUzDaVoLO0qFR4GygAj3x9T6DoulEZLqphrhmU/etxoEAPsTQd
5zCa88Ta8cESKCUOjOn2PdGOwAmeHp0mG4xwb18NQEijoDGlp2wzYUoDyI59WAUz
m6ScBXdl/NDBOi+oe5Gk6sAaAGUJHgTaDIdaw82b7Qf+qXnFlte9cecUv5bUtSMm
Dfj6rekBe9qG6LftZJVAOpW51QNYHS8uuBDJMIl9TdfCqXz54PddBfM6+lpjZod/
9uHXzWL9LeSWpokYq9MmyOpNMSwzqfYQAo3m2eY/H1eMoC5VsJOZhHakvq+58O4v
qPC/daCFtylouAjaqwYUprTzv2Cve2MqJ0WVNlkQl8OmeIS7K3EeowFj3wmo/AK4
TYUhd7D6fZf6wmn7Nx/LajMA884yGMccHB29lezr7fI1rp5yg5clXfjzrGLrl+IM
b4BwJyrN1wvglbmX1yLzKfzWgcoMqum8w5i/PU9AXeS4fJ1ho4USVSv200j8YF/n
7CsaWHa+qG2aSFxY6tTgNw3SxxzgVRFDkqYGD7vyklWNZDe3r+QSCcW2zoBhDAtH
D5fLH063X/9CD4yHkXzmhJhCI6+c9T5vHQ7CNrVQZ4Z6QUdn612JZEYwNh59bKFH
C6hQ8ThTJUWSh6+MAajYXimzYVKonw0FSRryjMURGeED/5cpINyca8k+B0fc6HZ6
il7xKFBoOMOwe8bddGOA/hZ8/25IVF9EdoJFS+wKisd03FZENWdGuPqkE9BxVU9w
8zxISVrmCluLF+4ln/IdDZ72sk4m7jhPMZGGvvmGsNYck9xaPctm8TvA+4vuqYWM
cldPNI2vSomTfmyhNB7svOwuO4aVShXQ86CoPJksDzpKfM7OSO31JxZrlEMHAKoK
XuHOm6o/lEGneJFkT3/9A/w7hwQ6CGyqCKs4s0JbEZ046nQj0cRGoKTx8GZNpfM4
M7EjBvYsxKRSovdbUK/r7i27ibSoEVrWWc4v5DqFg5/tIRtukBMqNaeOgzjPu1CU
MlX6nmNgS4ZUWX0a+piIqr82uHusX6BYAPG41ORoGnQsCf31k0nMXqwBtQdz9Wc4
HsT3G1865UX/BBB2eW4/c3QJw126LEd0H9cukvy2G7FHCAqbgALMQmYeD2Mqrio+
jwR5HIStU5oJfFRmsx02Y5BbYsU9bsydhccWr+dHOx8WMuzz+GH0WWBtt2NzGYHt
l0zCop5qjSufM+EQJyLijASRkfdH/JEZq4eQ4B2Kt0PJjkV7SEtUPOy2UWJ9fPkk
3QMF02gxc0Dfb2ZVBCJSIBdefvNmCV/4JLqIW6YdXY1ANV0wTN0Kj7u5A5qU2PEz
cCfAEdtVC+XokQAZz9dmYpPllEr1Wg74BWzQP5H9wBarF9qLOGRYAQrkOGtvgxYz
bAWA3NZwSeBnuJJczcLOIGy/JyF3Lcq7KVcYm8SGkETQSx/d270j3vuYAUS3YBiy
QeXXDcN1pgl56fdV7bjVe8P4lzJLcI5neJMH3MmijUH1fJiynbE2VBno1LSKn5uQ
JIZ2tq54UlW8AeoajuABRKnL4a2cJjfMQPOZlo7ABbJH+XTOck2V1kbwmXkqmnEe
Co+hC1CD9Sqb0GZd7B4r+1VQP3Dry2pO8FacY1f87LUl8Kr6nb6EJuh6eZZaJBaR
Z120pJK1RnHpKwf9NPiyfJrCYuB3+l6toLQDB1X+kz4tqK3zSI2MMwZkBWTIcTZA
/wv2EDNypIDl4Zzwh6QnUzkV+sN4iS3M3QTIsGM8eNcQPJpy2/DjFpA8b/VBEBP+
Ok8AAmTEWLrHN+Y7gUr+zbra79nS6NHYXW0DvZkTbKtHs0aYIj6CNbDVyJCs3EAb
0K2ZNFpJWC8wRZb+dgwiZuPC3XjAD69U/7gK0g7/t7OgcUV6TJgCZBFhhzNyijjJ
u+kEt5QBawH/TzoTquyXwFmCnvBlAqDk/WLGUaZ/Rph/NWKSzG9j+GloTxtjusaN
LSXo7XExv78AC6oqEnHkuIGnMUDO7b71Nwm/gOT7boDyNDU4worRYGpcynKmal2+
Oh+yg3wsnbN8htlWpKohsEwTiK6J4HaDou6j0bX9ne74/WoDPwSI3eQ8EZmCphjb
QymkJSOtyEOrr6nYmIRBqmG9gVsThgVNWqftOPTQXeBKrFxaWSUR5dLW9CGYVPsX
s3BHKmLGwtHxsF9Pa5jqtikNtv6JWadCMDjMkbeNlglZJjGAWpO986ekEp7ljVz/
i2Rj1q0DSIm5EnN3LXdco5H/Z9vuQFZbUfFCkHqTUHHsN9EQAvAPWYaY14xBfbti
ruuaTG4duY/XcLwnIAlm3ztf6H+NjikCARgYSV9IFTR2IDVATQ9LGsCUt9tOS8w8
4WHHYcDfPn3IigPhG/3kkK2LEzvg9qTBYgapEHhk5/sewP1ifs8dzCM9vTebi98q
bb5znq/Ku5eno3lIuPmPcjgkCU6F3Ffk9EXWFVDSLHFuXpL5UaC8gPtuxchQ5qXk
dB9lQgZPI+ZZj8wWJV0IJOPZcVi6bnGN5DD7OsWbMJJ80GNO2YXZQZ2I3XAsXW+c
5PR4HO/qGLoogUw0ezLMmJQRSIUKWORQJoOss4EPNVMHApj4wS+6Uy1H/Iy7vT0+
8ijDOS45dXnI12cyyBmaXod0i3B3kDE2sE7ISTP4CFiA35gouYpmfGBuyLsQqgBV
9OZjXd5kTU/t91TzomejZ3URXhfA6FH1dOsIZ7XH1ARRo8DiG3rBPQnKUcbJnOQt
qSxCHJ5xv1o7gVVJF98WeG6FCHGdK1DLh8E5hdHLqqCHvxPerA9bWAkeBixcE68V
FIE4aRx9sI9xKHh8OjZV6/xcM/qX5XqtAfcQcL8Cq8NXlfN9eHdhJt9sklfztY8w
Xn4wcXnZS1q8IRie2KgChTVt7Ke0DZQRHI969uPbRbfn5gSI6/BZ9/cXAGdkBvnE
iPLgdQO/zJfyv7DHZ69HFpu8aiJHhEm/Ulzym/fPKjnvXW045GhF8IxmWdurEP5R
keVgjA7/rJvnHaj7GHzamT8yTt8TNwBOhEgPMRphFxulZU4Sn4Q3XhlpVcczQ43U
9yOfgcgL59op5TTc3Wcesqk8pfx+OfXD2XQ95LIlzef+cBN72OCmccfHcXu/4NLQ
/r0IX0aXvKuh5qlllKvAAq6DAJDhXqSwwwFKhDRkkm4ju4vP1Km+ANn50Qf0u6C7
7MGocl8/98kJJCPuI8jOeyN/PeDpascDQGZUEi7f3s9/pWUgMy5OjJ4wz6plgKXq
TLvowgayXIOYvSeXj+2x/ZNwH5AEprbTOvYbFy6JRZuziFISRbPhLaow0tF0lGKz
FVDDXcCg49PIpukEwVDaxaLsL0gjIXAyWxNoU/v5DSAKRJVzCsvX68vv1NQ6MOxG
j2wToWvzgRNKNVG4Guho/tavTuspR71ZxP69frIU5pnEqBmmD+x0TFmrmJXLNBLR
6/4wgixIscRap64Rpb0q2/HnSD5BIx0169LIRDtV0jH/QjfjQ2baFHlESufdxu0x
f4xuUBeumSeGuqMv7VlQNFF7tYeVwoPZjVSoGla/5kKt2ersXET676LYpS8r405e
vW12HL1m8XMcVMp+yCCnS/6Q2nSST9CT5lcZZ9uxlEz02ZR1DEHij5TICUbBIS/v
2HEDySLnNDPcF0gti4jwpFEG/6/eig2pOVgyX37urRqCvYqlRMxRQfF1PKejCzXM
9MUo1jBFtIiAXgtbBXLKlmCNPFqI/6i5sy8DdV+PvnhJGZm9eijZmgq0oNBW5IJE
W9IeID0Et/pPmEhgmB0F4vJdLnDAwkGbdlmcdpTGgNd9NuPwnbYJvY7tVP1wQKbH
e32L2vn54u/72/nDdOZYh+MOhaM4guJXOK+AY9CUL28xA2LOb3Zl0peUYOjwVitJ
xkkPf18Vj9YJvSqQ+iYWqsTv11Gjgkyv6q18vD3QVQQzRwIq9qdV6OGF12U5RM3a
k8A0l5+e8KEKMY5IPlJROKWLfG6sLoRK7TmaHBxI58g8pbOlxsijXlU7eNHvPNv8
bMX/3dnx2qVUiRipXyPlJ/+MZs+wVqAHXrgEwrnAffDFU1Y2QzG6k1PbaLtrBP4T
zYfYlNw9SkCbAAqctz6hwlZASJLLAvcceXjFCFPcUMEInEwYP8F73ICh+LzEafM7
TWrHq7+1D32EgO5Asb5XakYyfTiBGS0pZUFl85OOVg24c3+ETuJDLqDJq0HDTZ2V
FQ4xfvKyImyABvzf4xbx926BdlS4DyQLDtT7pgyqfS9x/JNvSIaBmsX5Cny8QCDT
7qVBjV5Uw8MSl1WXGM4v28YE4kwAzleO4gGVHH2mCtxdexVywcAeFZbrCG3eOqoh
mpPXMsy8EUXHcbysdLcqmqi4H1xHxZavUDaAHeydVONUnnx/eqw4hFyyrxWzCYMw
Lt1RGBytymx7zB/AMwRHIDRtd80Fc0eAPN8YCd6+Di4i/8jFSHtUKpkiBzbW5Mx0
KRMfKeZIElZQp+1Z1sRCPLKNa1xtFIfqbTmyZi6WN+6tD20ooegzxR0RpesDE3gY
L4urOUHUjanvws/mvlqJcW4T5A3L94OcyNotg6KnIhfRySiydVkc90iW4Ltfa/jO
9ufrytl6xjUn3RUFFDINw/14F4WrvDKOteQccJhmEbOTmFDIIVdL9y3+Kha/Yal5
lWHj81M8Kfq6yeujRyzcJQ4t8f2cGR+9b8DXF1+MD+WMptUSdsIsM6OMe9bgCRLb
Qpj2xC1b/Di+QiM1fWY6pV9r0jgK2nBw2TjiIgkgQ2JVeORhtu2pnN/7P6tuPuD7
971qNICc6gybMW0R53F7DZov3SaJC+abTq3sFs3RohikxdvCqEFY1NvRs3z2F+pR
HZJcYhtQ4egqh60zEAeoYiRY66tPsfuThxFTuHFdcF5XdghsjMqfLwzHfrNKtRHS
6QJ9B92JBf33vTivcEXrogoRzVgf+tvvYlVAavkz1Rywww/h2lsjDTtjf6ebp1fZ
8WzLtvMvUAYAwUNcnrkkFC/6dD2pW3j8FgVRuzsWKdya4l7oqVabeCUJv4LUVvgc
NKuuoS+yCv+MR3bRrDaujtbccgRCs5gkXsqePoOR96Pv9dw3Dr/NqKFAbGgcBph9
Zcu/xkmpxghni5IcQlb/2KlVQ8iEMCnD6CmP8ojRDwzU5qXMzatXzJp2mJB0gYk3
LBJ7YdIp7HMzMvSn30q/sU3u+dCBHvWRm9sGjrmnELEj28uNdjQonCKjQIZVL3Xt
iDemqUZrT7zs2HaUVZ09qlqPKR0wSZOMfrojEgJc3kiJmAwvasRPAZxCHjyJjHL6
5wPyD+vARUNMFdcEDmDxH5MEoeyicXDATfby4w2pHECuTqAChexXr938OrPDNGIq
OX2jeVl2tHJHVfv3YJvJjQRLG/VO8tFmGK0AG/en4neFp3/BDBQG5I4KTOALm9yL
8gd4Mnsan/IvTAhtXp1yCXi4oQNLOnqyW++gO6nrObmtN3chrjV9PgNydbaCYlSQ
CK8ckWY0eJjDfG1hSbU7Uj6oMTqAxiL3FSW49ZCih7kzkyfqkTwS2Ioa1Ak+4px4
wW0S6xjSYRW9nogTAchvYpdF3Kv/0y7ZZoiX+y4rOlr9OwPh9NTzA25Trqu9t9TA
1OhbYY2z8oBJIwpFdGvkFUHQshl3Kygav1YPmmThFmk+e9+gb/bA76zeBZ1ACGW8
zroIsSVeiaIY9TmBXbrB3zCSCfpczU6lgxmgrvy91KIhcF/+bNsuS4ae+PMkTmME
oxI96WWSUoS1SWD6V+W15sjkThnRUWHMpz8fnAOyyQzzR8dQ0EWVmiUqYBBB1/DF
NVeq28M+Tk3uL2Z5r6DVVltSCfkWgs6OsGPPlaFxhBQM/hyqM+JW62AOSfKu244l
WnFgk5wqqXR2yFfjgffV9VQ5BGVog2dXiFtTPA32hT4AZeNucdMNIkVXcvUd11AS
XfitP8O8bPs0P0VGj5ZCdP7ME0Vn40Txlrv/2D1rdSV5BoUM4F4QaKXV4sUPDDrE
8DGis5yHXYePgeZPA0FV+qZGccnH57Z0HK+O/z9RUq7QevPZyCRFF7Mu8xv6SeUc
uhqDhBmDiIp0vGYLw1eWmqQSlOfAc5oO6tAb5ft6IXtGG2SHyr9D888zOewlojnN
qEooFo2mhKGfKE87n1NTtRR0B8rTLB2DpiOvBbfhGeRHChcL0gALpbN7h3iuV1y8
5REJpEhO6SjE1pntZwgFB/PehzhfyqOgK+oG7UqZp4yWnbDqB8llAv7Xb+BUM5kj
4OcblEx5CDgSwP93P3ttsJlvShHlrWpVgxnVuswFSbYhVK884Gfr/9B4ECQ6UpYe
R4t6cB2Eg9v4h7COIiTvF1v7QYc4jzE0aWGZ4cCpAsQYJ4JYZguDivAPGVppSG/0
p2mtEHC1l15wKhhwxOonevxZmGH7xzMtPrEw+rW8rrtAxhAhBPUy4jm8650Uxz3+
s2QGYKiU2WQ9a1DAA3Q0tqSNDgkz/s11EeMtewCRS0ltL7R+SaaXMRzQJhflrqoV
4tB/Ys55sUrr93LSTc+cMm6b4CVUg0rfdLzpBChUt96ANH3Gis/sM08WNwvsfoEm
tsJDRG7Z8yRhNm0fZD+RxmSs4fC08psyLtji0pHQzVqqTSjNxZ6rXWoAK29Sdcgp
5NSL9XEPRtH4RBUZs0jyjZN4WORuwbhZ+acc5Ju2PEh1Ncym1ThjrLWOQ1zcDVaC
3JCJYJ+c5I++6yZ7d8xppCRDFgaIQc9gRxnPNsBbzP99njZh5pEUJkgq2qp/XAJx
605QFbLSSwJoZ/J7yfAg+Qjy/Snv9rChnr53k+8xPzfStvgMzuNas9/7rZsMIdqt
EXfa+EHjVmf3/KnJnvc7jg/W6OXvSuJXT+R2Un6WvpFfcbwIQHMd23T21trNavMs
NwwJ3Erhpqz03Xu5IdMZk+bHUqpwXNOL6haLvI4aQ2yGt13zkGZImkU8QcXwDlY7
w6fXY+in+vzAb11OncyDPVSoTwwujZ10wcl4gT6RFZDtBOSydR0KCpc1hqyw3EBT
GzU8aGgrfTtssjMURsUx6xKqblo7VArK8gQQ0ktpeR21K1qIEmam0dVV+OERt0N3
LQ1JnIVB2FM7ll2uhx/CxRTjhK3hWfASFzsVYrFrRm8stH3CuHEiCj+vt8SI5OsU
+HBwSE8qXWWoeB0HQJ4t856zteKxqnjRNrPGx4/b7uITaK7yyIQNZYFqxe1oDbQ5
9MSEpyyz3thyIdHqmgt00yUji2I+PIoSYjXXdKnilm2xgohx10UxwuMPziIKxcfl
m09l4W6YSCQmwmx4odNxE7KPgVA1b+nPC8t8engNusMMOqZyaLNYP8VtAeX3oPeV
ffsJ+OEgZcOXzeWZrn0hb7RB9phA8q38lFu9Imw1ew+s7CyOFg+EH6sKWIDBjTVs
HLHnbLExBQHUlZbPZ6Kf3oGC6JQncm59Qwrd1GW5yZ3HrM5BK/iGa4sctgNl4oCQ
D0CnwNo7/xBgHRL6OXffZ+ZM/SOIe8QpU+fdLrSjEM6Oqcl55deR/QhVZuAye2jX
hOhhsfdu7K9hg0mfX4XNsuHpeFOOoHC8PMo3UAq/gWH7jx+JKweUjxe1KO1WAaLz
9VQ1bfpefqK+yBCxI8e4rsOPIXXP0pE7K7r3LMofIp5ioTpmrEDUm1RCPqM3hq09
tRLlMO3lKxEsGU6R8s21jwna7c+NB4ntUJGTR5VdDAMs9bBteIMRvpeE7HlAEe9I
vA/WoZ3eyWOEiyG+rvY0LMMTzp/iuQmvJLWe7YOHliwERrw0nAZ3qLrt/OLnJgCI
1x2JrvpVZGVBX3l6Xy3f46Gjo1qCo74hxhiokfusazYHJhxciV3OtpODvx8sZDBb
DhUv067OKekJ6r15T4gPPaxb+zLfRtqW6VkoKEulSHT1sGQuqInFMVg68EWGm0VG
BFdJI8fRB8FdSAd9WO2xCJK9iX4UMS8IyrOr1lVSXTC9ZeR6c1lMJTSF1V02GAgC
xX9DgTfiepVRs9IMkNg/wuoAKERCViuK+MuB3gea9k2FAEQ0WAyNHPl2i+wn2D+z
TMVfb2R22+hOtInIHIjB3ObCLC9o07kycKr2Un6f/sCPq4Y7fSPryyiUTxMfAx4L
WlNv2lkNld/P2lDnPlzhd390gZGJfASEHz5CFqQ8wS4xlhUJvVyYLSnHfKEy/ani
1iC4/9DG8LDVQGJn8Y9+aq4Onw0khqCnEaI0F5aGZbWJ9otXiIP5xtzJoRotooyg
NF//zttGrsZvZIMruh9NVhl/uZOII3Ks6sOwA94G77e3JsYtoqFeehMCinFlO1Lh
ujUxicykIjY/vcb3w0vI0jkZSWgSbjvlEwnF+e66Fa66fe6Jh8IsnfxH7PC3Wv2Y
DGDmGiQGXx97wR9V54lAkLITJd/fCzzrLHqJk/Slo+NcnthPUkvofT7u4qLzkfbZ
K1RznbcWoXnOC+F453MjuXlBkIogLLnH2QipqCmje0stCgoYxL7syPnfvHg0ISzf
6FM92fpyo99AAhAtp6TDR7O6ATESm0K27TQzDPkSM+FeQhQlL+xQp7F6vX3zHdjZ
7eOKopce+eaLVPBpxq6q4xWe4Ey4ZEm0cy2v43Asb9yz/ncYaN/adqvb54O8x/qD
olZ9rcVvsUsZK+BDrTavZ3aB3382c4l0tnXvDpClfoy35Paq8rsoubJjLk4ZyTqo
ABZ3UQZZ956zRNuPVUf1p8sD0rti+xZEv54Y3BJbpHShbZveDVZVtrWMOl/zdYDI
lDs3DDvJEYwRca72xe9HENxqNi2IpdqaKbRbDZywIf53KMW5zbjIt0GtKEixHnkP
vubtZoFwB0jtT3XXoEGpUmUaomhhsPBEOFRH8MjaYT/jix2gZJSIMAzKIH5nG/lN
8oIz+jWZYL+jPCChfVjPBhxlNMbvOdaEIpISQS0e/WTKulh0h41Z5WpzOyKaTwcq
iRRUy+0v75uOBWSnIla/80EcL97+4hrT0jJ7UHMco9MyLNZoraNtZvf7j6S3MnC7
SatgESCzBpG+uSLAWflHz/CRZAeNfzNFTpA/ubIhtYOwKsq/zkYqnrsyVvU944UY
4/z6Pdyi29MxJqgJN6RZlXCcmn4LW2Rk5n9cgtwk79TKn4HsC+uJeGnf6eQLgHpJ
tQ/+uD7G0aXQwiRd/WErKW+QUItYkCwTO11wCm4zofiMkj8GVz18gfC2r4qp9AKF
nZQHy3m3fl1rq5NKLDmg2LHsmpGUmXgjOiXIIOLWvp1mga8fYVRgD48wUxnDTvMc
tFFjO026vn09sPPHSbqJGfGDX3kDKjW2EOKgGI9FACH4JXrab5nlGaMHQn8/BMjT
cCX6T18AMQqF5wbGTqc7g3g7jFOnZ1vE+w7gjNYA5oUX3fgtJf3LPdVmtv9KKKDP
q3Urg4QPuv9tatMbZKbCkVNtLwS1BuLBwRkvEdAJHFxPcwe09meJiWTfcoE0rN/U
oS5unSLDdQJWfccKaXCZmsh5010b16/DHDV7Pg2EFBmYk1YVLGQRTCiCBvH5fOPx
zUxRPQ0WstaVt4L0xBU0Aguqv+6mpOVcml7dC33MBNGIDGm7SG00/n2e8LEhnUnN
QH3ZBSk39qVpT0DbAtiX+B9rh2vp1/ymrnBwsZlYevz+E3xZrT5IvBezvQVKjH6p
9i5V0XUnkwABcowrWHi7+4OhqOtTAMrMTPvoxZww+nQ02Nme7d0rZioPQBiXvX01
wFGdJeb89ymdOA+DxJ7WEkSJk5C3zENMClSBrPRjRj7UEQW4EvUS7PhVPdvEbACm
vOz0PRBY2eTuFCZUpg66lan2RzFyaHJF60K0dr4QtxP34Ovum6C7D0RO6+5gar9l
5R6vrLdytXWuECDMPMLbMLknoHRby/X1895SYJLNqzqkbfKgLCSqFyxdQtqhFXnK
BN/sKO0aAbE6vUoW65uA/au/jm1tLONQnRIIghwhWojzYY7HVzEceN48MgjPJtuy
eEH6B8u08XJiG5dc5229wwZO3ERGgmQQ39cpiXuGUmG32zhAa+K1oINIzMxoHur5
fvjIo/HAnabSnsCCthK6e4pt1+V9gaFwwwrkkYO6gOwRSImVZxo/z8Oasweceal5
xnf4diYhiwVSHWCmgshHjBCGMyFHmE8hrFXyR4OnCAq5uZ1Fcgm3DfU45+YPA1Zi
NkcIOn2YyLA0xlrMI3DzYWR8yl/tztGcPUJd7BcHmmrPi+FXKxNAeQCl1FCmKhx2
CzSdVzMkviyMxqWY2IhxXoCHN/ufVZSRZkPO8Rj2VJw0nQprCeb4qVYu/msl9i1c
WKvRsKWxrhg4wYGQjVkGcd6ywDOKP5fV+4nT43mPKFe6+qz9W9gH3t81oYfabdcF
rSGrn/10/6TkTFS51Mw/Dc0cCy6rou/t1gYcgIDEftk5fYdEEEaPTlEwjLLoTUvz
2/1fimsBumPIg+nKnl7bhqSMvMi+2kUkOSTFeU02R1Ed8HNRt7kC5SyWCH/r79PJ
sBfpzsH9N4nR172riguEW3IY4m02tWDhPgh/k1s/3HXiKIgmWCOk8UJwYyNPtE9x
NFnO6/n1bJrB22r97rCkxC1IMrBY+Qp31hCu/8skMRWgcbT31uDd5r62+9W07tbG
l3Jc10163BUQycufaS+5503F/nVRAEPXQqTGOAV6CmKuoHE1q1ATKn7EGLt/YQ4j
C/6VZe4RFuNO81ym7d+54nJNULTT7jxootdlAVTeuA6cjlwsAu6eMYRhDE1RYPqi
mDCb0OdeEr8Ww/vutDetVpW0JgawA+nai+EvGq7Wj+w1hRCsksFfqCQ4WRGZsKJD
WxWqOhvZQ6TT0K0M0U8kMEfUf/ntE8WPFbF7jZ2OVG93NdAUuu5DrZIPblSQ4xDz
UXw+1yDRSP+wuTEcgti5WhvfojNfnDDfcYa/UvVwnXt7DxtRhGCrtbrTR2Gzo+fV
2E7t6bezU+qhrtyejBhK9sdEbEAdcz7xe1XzgvUgqSOfQeaCtrEkVDacf498ppxh
w/9fKTRNIw5GvfFGcYU1heWxVO/p0N03kakkNJ5l+jrEQCNgWD9ypaWCuhT5PRiX
S3+x9EKRcBB6A4uHGkmZMJd6exaA3lVhrnoB7hRx7Q+M0xZ7iSRRD+KUvoq62fcV
AB6c/1127eC8qMl8RFOg5f2kFkeMk+F9SF8gmSuA6qTXYQrS0PwzICVuzRPadgUb
8Rx7I5aj1GBy5kn/+IrjMBl8Yzd1caV0r689NgazrGjOuLlccut01iotfYgFlQk+
KMLdS0Hd18Gr4qXcLRPB8Z7rdLyB4g7V2i1MRP4z/LECd+/giXF18xIjXnVInanb
FtMuDOlNhVUZSWBP4S3CGkaWyW00V+cXz64DT2TWxEJJZomp65CTYXIG/VIBRiXq
GzfMCRaNu4sEHhpL0MMd92IKPsB7n/WiPV7qNNuJhGU7Kl/61uD17emgV9XSCT1X
QbOjuh2i7dWleB9Bp1ZQqgvPKi0SXfA1v4gcW+ZA24xOxF9IDleVNybbVCQhVf83
TkfBWSBWSzD0HzuD8KvCDzYtCpweT0LBPu62ugt3F9Y1Zg5cCUqp8W2fVq6f2uln
+Q/GEEJl6i1WZfPrMRhpRlMLm8/2pmDMCL+omZO1pidx+0jqIgzOrl++3Sb0bn8n
k313AUo4jX4mB/3XoxB+kzfeB2lxo8ogP+tjbjz3QErPSO5fU61s4jJO0GcF7mMF
p1MTUlFkEQWzrMUtNdRQ3tvzZJ6dGfQyEzX7zEJVaUTsLOA8wa7himhZKfhC6NcJ
Kjru68pr68eVOd4hesrMlNkhkqO43VVCDSIe96eacgNPQ+skjwhDmdzMKwF6fg5P
Yh2lbv1j9ntXUB1wpJJVTASDEu3vlLkrtBh/xrHEIM+BPnj2Ho08ML9fOUiyPblR
HClD60dyMWIXGDKWvQUixaCzLvORY0GFP638sX5JOlKzlYu+67o4f9LkMkQVJEOi
OhmMtzIXu/Vd3r9eriwFt2FgCsL0Uvie7boHadOK9IUWAa76FedZNIJeVWdLvLb5
5x9yI/TBWOxRo+kGWNJSbl9JY/WaQC98xW0GtpOLR5xmU6kaW6aVy/pdXEUvIHEH
7y7EGEbWu8aRgCxeoL7T2XA16p4iK5jDCW6uLr5oGn2F8NMT1lfaomLQ/cwHbjnt
XukONLv3lavVNrly7NjQwYvxmSVyKyfA+60xase3ArtIwEhCyxLQ1OUy4nLKNttE
SAEzukld4leYl52uGQabdE/ycZyHrXzqbFCwJ/VdTNXELtgF9kNGq37t37UBIzAT
aah+upqX33zDgMe8LKOkW5sJME6nY8tC2FTUWXf7rg2gZW2yF5QdT8p2UL/bwIbd
38F/GkKjWoEfAkQXVwcqyoGqyy1sxj7d0WWnpNPtgCNX2FJfI972PQ7YnbdITHJn
TUYCM+xlJArUodwN8mEyFruaSVFqFbwab5SsUso2R4G3uoriQ3YAZuNsuM4C7GNP
+y/CH8izeunZ0evlWyZv16zH0GC3FmEHzo1A6X4aoE0W19H6k3SshCw9zPhPP7Ol
989aRO18xm3UZh/9Ss4hJu1k+U6nXTVivAtCUyc3R9AKGFGGYl6lNRDbNAH51pVt
SJkqbRvIVzEA4MwCud03fV2eR533KR8dudRzOW7ChopPbPj23arXf7iiY6nK+EYL
NbiAk0S68iMPRFaNeXnpVLDkaLzD5Fi3+M1KavD/EI+j3HT98Hoh88zYk6AkPXzy
ggISYGMTi995pxK+EBjMLmEtGMF8ITrpBNjefhfPBazhzvBzC+RYnRmG1KQA2qxY
iVEZtvYwOmR++1j0SS6gg9r4+kPzNYLD+jK6FGcPmddIhZnkxdJobe32SZqDLdWM
O1r4ei2l+CR+n5nR/Z3BVYDuTsYUFz9tvKEMN9HHRtNXDurn5a8h0EXZWkqN07J9
EftZYSJjGxq4buy1J5qLKMa8cahdt275c9cwi2fbx7cqw+z8cF4cxMHkHzNFBzXl
hiHOR3vmnW8vuPxGdOyIebGOK4H7KIieyvkXQRXrWeK7bx94WFNikwHHMl4fHzG4
nCgeZlNDQi5vOMEuqgYmqSQI0UM5VuYeDf8p3/7N2c3DvgMn+GbDvse/J1XmICCN
wccw2fim2YITlSFEniOEGYr9+FHXWQ59AKvWpw2iy/4u7iFWpsNKKqBAN+HQfOXi
UheoKB5VPk02D3czeFMcZZu6Ulu/PRx0niPHJBUBTVuybq5tJ8OuMWn6OHEB7Jqu
Ttb/jaGO5IXM9aePjMKALRX9N4fYC5kNfMOrRikVNp1ZVwQcmeiyXvTL4qyl4Yh0
98S67GbLNqYoddL/qRq4vC+r5scLCPThbpsJJ0vuDw3XU5hpNum5/hrriU1SOW4Z
YSmiBpnXK5DlQY+MICEq7xZ1U+8aB+Df/GbIVV9fsqzwbFfHUGQ90fUrhDUAc7pp
BQ5pzZbokJarFtD5b4+wPCSuwbcieEu2xAofUWflQ7bliYSSICxfBUxbIzVuW/0J
kqMOJbsUuj8iEvlae9Tw5LlSPVsl81sMvjaw/laqHdlkim3CucSA2qhJOaczU/iX
IlRwuRfnQ5bx+Z61b1pJQg+qNb8uwvVvZwHvjr4MKDAeeKpfqW3Oyfm1VaAHmOAh
s+nCCQatL5mC3TMTQt1GgNdcP3r7AbY8rO4xgQI1NJL/vuYnTPVuijZiFEe5Y/wO
EcT2PS3BhqvIWybrjinClJPEkAddnBlPURfKcUo1TXkAavTU51cgyDJJsJylw0gC
tMV57vrNHv7nRzMFJNFcldNeYsk34+LSkUUazAe5BVKFLku7aClD23k15oyuH3nc
3rbw4veTYUwXneaan7++zYYmSjJ+J/ONq7wpf9s+vBB3yFhekvB5oY7nFtgYeY3T
0iki4ndM/sg+1unEAf5p0fAKLrlSGrBhX4C0fPDtv3sKb/raDH76SIdgV41zN5Av
Ec6uVxCJRo6BjV1d4HCIUllD2N1qtyoAfs/zBXWx7foQ+cxxu3QRcXwSHBYPBbHj
oNLLhChkDNoqvYLMSx6c2VLfZ7XvJiDYm4iTGj+d3+so8nCXhRsgf/BQsPsU6bwL
Q10jaoQO2zWF7LTOn5Mk84QZ/+FX3fKEkkDGEUWPOGQ/oQ0uxEJwXo7maJUrKr3T
cZv8f284GdWgPA3Ikz/nHfmFEJxx8m/j+uU8ldlF+t4TTDfYkgmE8M1qYnFEMpbZ
1sNQgNaBzZe5bMyPQXHL8eWX0okHY6xWEh/2STVETn/WTyKbWTvTjfQUGfOc5q1o
h604MpOZDJlbTZeRJjj/PZDDf8GyolVe9FV4i9eRhXySCyCpN3oA9p6hm4GBe543
HrDoPHNKrMpw6xVkpR6qIJQvG8UkGyDm08WuWEWZrLScLny7KiVJOKSq4feQxND2
NUu0hgj7CTKWSsTPxlFG5NQePH0EzK4S31lnFyrG0QFsWJnc5tXZkNDmr04E/YBA
EhUfbhNsKzxxsukckxvbgt3g+tBPROLyE0bQlPR/LbCRXDc3tEtFBMj84EJIhsZK
HLg5qUp8WDbflJLgvYTwiEevSt9KPyEU6KZ6vf3xlCYmsJgatyI/eWUs1EqiXRTj
BPHRaL0q7gN7OOfwOK2T/T5eaNCxBy39oyYfTBnQrQBtUXsElfLjdMl6qMZE70AS
WdwPpXxIQ6iywEMdEcyes2PxLRXeQVrFfXnL5g1p9iPQ0vvRk917RPCqlCt2G0Wd
Sx+iE9qzdgJvV65oB4Az5SZIdRavO7aAxIPvhgblfGMyfVJcqOgWJqzJxk2LujGN
ZQTD4LaipTvk17Fr4Vlf0jCzgbaP90OxITzmSGsTqYiJoHl4MkWi6GgCfmLVPbZC
JdFCI0Jqd5DZPQVzxUjL0ZipiDKwikscdfWamEscbbGbgr2TppDMb6go8pLgRnqZ
nwTrd3PakV5GQ9VhVr4u8YVU22SwMD0ylBVZEiaFc9bbCzW+WASkLIcwJrZlviJ7
8Y9Y32MhizoNQDZ1ezeywUp64oZu/ra5RwDyq1ol6SRI90OSWFTgfVqJeekxBC9k
gSgl+j0k8qUugCPoU8VXxXRq7NpL6NxyPY0eq5WT1NTxNaaftRX0UR9XdP7UmB1+
qcjD2MzG2tTq7X04B8z4e+kbWHIjWOGBnaym1D1mcIFfNTlYA01xPJCoFOi64H4N
KV+XesplfaqmaOhOjhILoiB423spSNof8dsGoqHOS7/Jkzjc0lLl+jtOnTfOMrtj
9TarT+afWLDH+PWW2mBqvtZUnHGtqjDOLPfiEEMQ5BDuuH97Gde6LcXeD/mcvEQI
bNxameSl5pf0oySrIAVV/F0CvppGboVx8RnmsEuFLHEZg5t4XrzfrTmxYejSF5fw
CulDJ8y7qnMUyIDYlp7KaJxxF+tLqfIqlhL1c/YThZ9jxSFUcm3YpJhYPAVxdnvc
QjW/bZTkOLbFrmvBZ3CT9nlFXxluE1QFYqSVvFgjMW3Ox66o7RsNIw9a/LT1g9YA
KqM+G9u3EFvzOq2rJLw1w95d5qg6FHMRv3fH8Nz8IQN83AXPCpqUc5lNXtVi41BZ
OPSWjM+LXhQfkMOTnlrkLtISG0UusXnL/jesBXVSJEpptHUQWPSZxdDzknV/iQpm
5QXOZNcuzJvwoWIBbAcgZcNXvFTlu+dsQwJBsRYcXqXPCW+klj5BUnIc9fKHmWmt
HPrWvgb/qoPo+oZQ2v02GjVW6czhntt96A3Rhryh2YpawzYfuVNKSpPgzfoFk6NB
uvDmRkzsgxz+pqeL7Kj/4dkKq/rBqu2vLNuvO9dar31uk59UwFms9BKlBUNH8bpS
szFT8Hia9pCgfw/0mHohj6LNIBf75SIn1hmDq4bs7/wfAnA5ILBtQ81snWtHJVxU
CvRxZsP5bhs9FjpbiUaplzmmYvOCWjkJyraDGs2tzrWe+HVFlguRrCopVOyM+7Re
73HF/rbXz1EYZieTkpe/QthpuriGAgca6spH3HyBdtyW5/5LdIw4jv4TMoVBLIW+
Ar4gSed13odw0lgYl489bYgQSnAqTAr4DgRmw8QwfEZIttnayOOx5bK08F4el48T
rswWI3cv+E0DTpxaSz/tiTGxqHKBZGyfrnzG/dnGFVV6+sVdAnxM4Bho7F3uhhLB
25q2EsdVUHuJZ0T1xgJyzpqR5tPqcykAWyZDhGv/uRycUTTvfF0UZDkBbIqvQ+Ap
0CVXo4cbi4OIgUWUBpfYeK3gRi38kk3sbnR2s/FDh3uKhNfXewzDVkD7TjDfRHmH
mERZiOIuFz3zJxZWY1gskPaRVImQJQcKA6yi3aFNxy42fBywIjVPU8RuSay/4zt3
jDiUP9iRgbmzdHDYjh62pA3LmcFITKaLiImuW8ucHXOW5JcrxsrzM/uY+ckcc48x
ODRsB3xdJOZYjrhFbj7Z7F/SI+etEdACvdJkhu1PRRXz37t1qd5afbTuLjC25r8c
FJY6aUIVfwhQ7tasLq4oUsYAreWldFrEvARr6NWkot5tA07OWBbtREccMVei7fdI
YXVKwmLkVALeg6nnobIsrPOW9KDoCqtj/HPp+WfXJQfWSm/oBe9X2pzgTCluoqF8
Ws0W2uXcb136jMKopLtOmv5hWJAJ6pT6yTTMA6yZJct3NnbR21hq1sHnUBaS/H9r
ZShJ7WOM1xxISypHCmihxCeCrrF93ebyYcHEZacEWrYdp5gvD1i56IXMRLYhEYQD
LOlkK03VdEAxaFwNHU6wNekD95pXCcNqgwr/qe0ev3vt7b23NnhZbX/XOjaduJBe
qqEkxMRlh21DXA4yI9NtG2zFA4yrIBgmXbP+JL1vygWVehtXVMcB1yoRO78F7HVL
I3593OktE09Wlvm2wkZmYsByVAJ6Qeck6fFVQIKp2Kp4pUrrRedoM+FDvqqV75ZC
SKVWl/T8OnV0X448IPXtQ35HhlMaZNapBKQ9DaVH6fO3Uwpp59Bx4Llu1gTo43Uo
lhC9i0JdRWSwFiQWAJIzsZ7aUNu0XFVOlXa34j2w0HS07szCcJ92kg3ROp89WRFT
R39gRcbOVYQW5zlucPTLxvnkGgkG4hbztpuuxOTRHC7C18VAWLdGZH7HpIMxtn9/
tIUUUSzjTtUrT+ELXGTOgE6NZV2yqJYAowdAlP8uxfahJuFoRs8S66Kgz5eWpDOk
LaZA7aaMhVDeO1AO+l5tgZi4tOTC6EYHFYAdC8bbLlxZ9zXcDMR/qFPV9iyFizPI
domadU6Feo/qXnZ5gpH4CKZfvBJPq+Gg/q8CdjB3us4fnRj3ekckoLAD6UKx0Mup
bgM8QuizOgAvnmSj14cMcfdUVEdVeylpmDi+NtnkSm769mQxlTqfMoJh/mwGx/R0
rl3h4LtejGi3LRwAId+nZ075kLAFG4+T+53mVNp1t5+RbfRqXukgoQ/wNL5FZSSj
3putrVD9+ehbLXQUORW7bbwv1LvlDBEBwMpAsRVADOXvRsXhre+3X9KWMZkNqtz0
AB+05Qu3yzAS+pA40Jlr9Qqpe6iOF24ik42Bv9Ej3vq8XEIAXS7qKnJZAXZro7Vz
sF0f56Gx+h+z8geXVMu6wKhPeiONNt4HFuCsXAPh30B9Ea/Kx1wc1Cg22qXWe3Mu
LPrbrugRM3J/EUHvTKVyRbXsxQHB2mMF3L31iAtj/L4oIgSn0GZ3gPbwPvLPRbXv
uHbZ0bIDOY+BuyKqM1UrReHMtptRUDY1ENOXjbILIEDxxaW2CgpgZhJXC9ijgmao
4m8scumc7fJ1g94frO7MacT2NdqlePa6N5tvgqJcUeAIz8gmxVQ60pMqYXIKpngj
Sd8m/XJdmQE/UVBAP9kttxE353GkTIYZGANTFYEU7sQN/rVKfb8gVfOiw7X/sNz1
9AjROayubg6Ptecx3v/6pjinprNX1g2a6MVa8ZA/m3V8cXYz+nn+OjsHcBaXbo9P
9giXxc2Td6ANTRzfzwc+RcJzBx5bIa1FiAdkqktluCz5+GnjSZ1qyQoHyxYYaYzA
Em+5o9uhKCwKRyrW0rkR0Af8ZHIUXt0VlSNzKIL3Djihb/p+EkOK8q1JAKd/Lr+0
ZOuhxtWIEfx7bctE0MyilSjQy/teDZNyIzHGK5ztNXLKXxoa4wI6o0HsjsHIRQn5
I0Q/5iClKuiAFpyFzmztptZJ6pxuipRh2U/oKBG5puAgzNjmPscARNwIGOLF75eY
1+1Ov3TmemV92F/C2tHMJWl5mxMXRt5VwYGqR3Kc5rkvGe25m8TQEGCmFA/q/G0U
GDWPu7yaIXfCQDW8o+5utRV7XyzWwxDoa5PKi0/PWe/4W8HkkKw8P1Ez0FE1m+G+
M/jPJYhkEVU3XqfuXwYlyIyIeU/h8VVzPxrfJuwJOWwsGqgtGvi2YXgC/WEh7IJI
DKnwqS5JhLeLc58BoVKJvLClUrBdaHie1m16knbsVBY0aG1y5DWGMhIx8q+ehtdF
WFrN0jReDi226ObNcCAycd2lgrpL3YPGLPUeC99Xs2cfgwnbMXGsjlss6NOnIljT
umHU39zfQ3tgPysZZ9Qn2Sgrykxz6yZvnLlys8oce+HTgWnbES8QzhdGPRdMEo+7
CBh7ivNnu9rjz11Tqc4fjl5l5AGmxNfHrahgrj6jFiXruGSa3Y5XyKFf7gSR5HYa
LXWg5UkPVmG0M+xl70vJewYBAtKs+oVeRVHRJHOtDGCZ+EQqR/4rJhzJVDTFR30r
Drj9wF23t188SOvNsPBwwBUq52zilvYTcsX+QAWVd/SqkCqid6aIPYKPtlIHRndE
motaxMmJhPNXeiZuvzyVLKql0VV3U7BAlI0hIJ5DoA4DWiK2tGKA5B4Xgk9XYMnJ
hJ9OW84dB7DKuawX8ar6i4ZIWfWAHLFRSyTStN/3s7l5qhH9dCVznHr5mbjoPjvd
zjSjd7vHLqb/pHwDGS7RNP5sStgsTf5yODxHbo8Ah5kXDr8RYZP6U4pBRIJllJOM
oYZvUPMadXJGBiMYQrxqHSNJHgUDbCGCYCYy+s97vzW2Cxf/JhU1wC8kNdX+5DoV
ORoeUwW2EJbC+fBKxGamU/GGfxErLjU1aKgut6vRlMej8tR96ggNAah+Hg9O//tV
yD2GissewafOKJ0efdBb0VqcFa+sOPBdlEMqejCOv5Be1JreRYYLRt45E8lZIWcX
U3tLhLNJmSyMeUGhKBP6qx0Z2skIWoI4ENeUwd2VdbJQJttfJCAAcofWe5CPi87I
vcfU4fY4P2llUpzYED9x5384Ai4fX9Ck/0z9YCvSmu4eLrSVFIIJKbGgwjvNIuCp
CbZ5W+ff6nSTy8/uw3CTltLMUrWyxqOb8gqzMOgp3YlynBw2BCSWtO0fKGRv1kEX
9F4cpyHTyEa+G4M0Dfb7iiVteP7l1Y+Stih9Q55s5qNT7fCKkLJhB2d050nkdYZt
q5mctLlTkwR9imZzxaoO2aRS+CRc7XSprqegPoUVzfR6xCfSKXuFkW92JmmxJX9n
2LFpaAol4H0Te1Iq0LRIFxShAsnHmIH5H5RzCcw61tREMMgE+VmckySMpDoa5EJt
sVYgIt9qdZj1AmbHeD2JPEVlsTDta8d+aT3CJIH/EFO9EQZ2MW1d7l96BTEMGqMK
N8O6O67zdD/f7S06Yib05MhC150pWK1iWxpb1tpvwOAQ0UX19OQWtugjxjLQsxiu
0zfa7IxE9P5sLHXahd/WLoiy3ySXIRc7s0oYJ1kTOsp49tdrkqQ2KtkrPiVGPVjL
PzDyCNgKULfck12VSPfwNQWr/Fhy65JPdtnJrC+m2ktOZ0qw/z4jnNXc6VNc48g9
VMxY5k+sx/W1+/TDObHhzt7WthQoz1pi4mGe2RUtRPP1fzuSwNvOh2VBDBaaMGW2
zPD9INYP1aOCrjDKaxuh/xDi5Y9sppUAQkLIwawb4yWfF59wy6HpziFzFJ4TFQa9
F8O1VME+36SfCL35kR1ZVs4B4VpSgsWF73/fR/xUG580LDh8DhMxwnzAeVBMVw3J
AlsmJEGOpAVU1AC7VPompZ7a2IGIelQj9vKU/H1a0kcle4xsnkQ0tygFixUHsP5n
Bdpfv0KfKTyP+aqXYYDkhZepctgRgO50KChwHwj3v6iklayw470OJrHKVYnGyp3R
h2uKO/78PmanVOvyDKgAa1ggSSv81DHy58lgYwyhEocMqdOlxcn2pn2q70oJG44K
R43fZN+hgA1Gkufbx7ooF2YFMibHtW0juTtPzAYodP6zs8HaJ355VX8Y0gfKXcZv
32prHi8J+ZKu5QB10yGHwY0eETLqIijeBZTfIOm/FVk9yp5Gl1geowEKJeO9R98I
WoAU3y3+NJIanEUZ9fsxGlmzvnwbydCVSrIzLXB3GRtl6GbLd+4fhBSMwqKZKeun
zY0Vi/eHDqTnWCQooGoD8Hu0tAu3/p9gbl//H6l6i/FdLr7ABINh9dltV1Cmgdi2
pgvbEe4iauIGwYvg3MZDQXJ5ZV8f2wJGndqppDFwA7Bsp/hn65JgrWd1U+uxWvSQ
V1rPGjdW9dcx9o+0xcCI8TsI+X1I9XyV92LElXi2sTnOHP4js9IA+54xsHZamazq
c87zKqRzKLo7jB4/ztV2l1NCQwipQ1VfsA0fW4M1jkujFu6hgsGNSn56YqKUKzq1
LBCcOgLeHNZYvKVdMaHgeSY3q4vBE8KwNl5yeG8qMcgvltygtbWE19+Q7G00hprv
ncrgW8CSxhgalHQhzI5K4iZDjILqlBCpfOpTE6kX6BgDEU1vatYnnl9YaDBz1lJz
XXP6xqQQjbgSKOuf+hOFfgMqzsVYK44uuQB4BRKsnsdwCMEq3Gsg3SMjpzchI453
5ykIAobBD26yEeMH3aNM51dWiU3dMYJkG0v9dtDm4D6nQ/0Ehs+HblSYrRvWTsmR
VBzdqpXLSJqO0i7Az1jHIg5uPfX7Vb0mve9nk8qRJUF8Qab3+D3ls8t+DpWFo5GD
CqyXrVmOXcGT52ckvJIUOs6Mf9/e2CzINzHn2b7SoVWWKjtSN+nD6YYQDOlHxXEI
0EmpdoJCemiAa0uDjs78NJ3IBxFjuY901o+yJK+IrtXP7oWQEdXdioFcgDuIMsoC
/dVwyDi4a6p6YYy9L2u+jfNqoL1ciaMDQlgLNw2iZzjDu+p3quyVkx9QxXtVRfYn
/slwj4gjSD+RVtpjUhRjjsKSFaLr009bztz4oTJyEmf6kr2OatT4nFztT0eAY9TO
DXBduAAl9CK+PG+OImr4/4EOsW/k8XkbK6U7QxtmBM26q9E6tzl//Vwtl/dm2LC1
MzdwFeR0fjO4Q3A0l9sS8+gxfz8XKUQnWqQeVwAQOw3CKBNLhNv++z9EXkIC6Y7z
ttyoLIMkczhLNt2ySxgKI8SRwZ/qmLswjQzOeu37tw+b7wntZyDMJZ7SQIPw+Xbn
3XB3jgezWzbgRUb8g6Oj5KaGx06Kz59Qn54ueRxMJvhF267tnf/Fe5oDJEULK3Nk
6CVbs0IWGQvdbVQvhxbcNccM96Ai2msU2Kv7wUXGAg7Kc0EsozXpRm9YivsFT/HZ
d41cXcNDwQXkIhW/QUhTGeKNT6heazofJenozw6sVHYUoyaMBUokHm4n9WhnkPqc
pLFlc9062b38rSLw6DGB8XNY+lMa79Zhsx8jqSXx6Aqu8nx3oM3cdlQYiAIE2zLB
wBdvD4TrlzgJJaJpVCO8ODwZ1enxFX15wsf3n7wUs7fGc/WDd0yViUJaPoZ75G0M
kYVsvhebHhc+1Jvwc/zwwAOXlWO0LUWO2oGlIZ5fDRI+2B7NLEGJVsmnwReIPKCL
QdUMhsdkadpYEdzzgsuLX7MYYcz77bFma5su12etoo5zmgeLbRAUIT3pUB+LUYtG
rNZ1693cbYtDkiyKeyDVQnclXBIC6IlvL1bSNAyI4VapAsQc7pHrQ3PZMN73godv
CbQVP5VuaYsT5+TCk/ohCruluNImSmFg3Po9vUcdxpmxZk5EE3eEGvv2slqCXZll
2ymhBfWBzZGPJpDfVFMXxPYdHlYuCSOxyyYlEZUQqhrvMdIx4cTzqL3gxbqjKXtd
Cz+Euh8qlcb3IS6uGBRgvaUF6nlieJ2j5v7VMVxywbgGcKeq6bhX89MjPu4fTKoq
sA1Q04Y2/xoyIaLTAKozQw8ja3YncnmClqi6ATyqwm/Hjd5V817jCnSXR4ulaU38
7ewklomV3Lpc6BvvvZD09WH8CKSz0C4mM1dacxD3/ngYTucBHfGePX/MYL0/rMvJ
OSzTIAXIJgCSQb7JO2CY7BIGxv7CI/alqQQ/L3HDvqTQfMmlGcbJ3XCCy2ribvgP
RabiewOTThNAndHf7Z/Ljp46JtAT1RlflLyYc2vkdyJXnlCuqBrkoa0rD9ajltvV
3KZZEaQeeUDnGqL6Rr7KAM7LRERFfpWrThYle1guqo4GOX7yB4d4QTYmrno+4kTX
TPpqzpC6j3Plv2p7gMOcwliwaAj2azOGoivY3H61L4/HQDZruqtfLPTg+4SmPy70
7I4LPyzk0PjTgUHxcizIeap3AjsyOrTAXNaeU5xMjHro6VJrsWyKhc/zbhwd+vfB
4xIt4Lsauy5lhlVw9Oq8kFLHmxJOeno0U8cRKPZaTY5kI9DeVmrwpwNieIIUckK2
eOhs5VbzmwBM8bzLUmFkg3kycsrtHplG+c+gfeLq/Bf/h11rtjMEqXPxkEj0ooLy
AufJEcxQ+9WMKUkVbAFTFYkVqTxWz9i6CvZS6t5T9Wf/UCYOA2QvjWvALb2vz3qf
CDNPpbZvc4mmixL7/+N1qJFKR77b9+vZSBg9pJoOw2QyR1qbxRQQuPdPjsWhh1aU
9W0MEN+qXlcoOIpGumIUpWFlU5g9WRwZJOihj/5VrLuI2o5eoYXVybJWBh2AqWg7
MMQ5cPM6SkrZcsNlv+eC/A5VnuDLp0IEFoeigUVRj5kBjaCPWfYtllJ5d92rLDyR
beOtkB/qrxP54ZzVTCh3VJOzUmVUHMhO7gFlfGXO1+3tTAioSIenmH9bdN4DAeJh
oZhZ3p5dPXbHMAPVQnczdDUrDalVizlOO42DXfqDIYFiOZIdHNVwNIJCLSlC4mJa
EkHSj9TbU5pDjcQ/0T10uhA/EmLbgDy2SDnHb1DskPfrYJdcU8Q+XgvpI7djesyz
25uCx26quVF8yyz0DlFp+fHzs2vrHUJXLcI69pGLqJ0mZLUzs7SID1U6A4ypiFkH
uf9aO49LexNOboy2p715IMwQBNoOQWrJK70VqJpuEWqCP4MvrBLMGL1CVC/6now+
1lSk5J4dbUBFFgt6OE4TqZyZefsrrlJCtcycob9h9RCktgfVwIictEvMKltF7lGg
Ft78Z+FB/h3gA/UpXM15RKeM6McCN2UpNuB8wzMBdpwGiedlQxqF/FkJmARIQsWt
GnutnOHDOXULb5i633zou1q8TGzPk5tk6sHj+eyywHQgY0l7qydaNrbUkXWOZnUc
IIrvuCK+1bQ6Ao0kTSl8uERgAJFMvTsD41cRkSik23z5m2uwJ64IRq4FdYmWksFX
NqLQOcbyAaN7UGF6cB6wvM3RkfwkrdnOII0v6PBLkLQo9blaRtC6fx0jJ++VXTlm
Zf5xSmALG3s1sVUhi3EeKuwmv2u0XVvW7i9aY1saqbkvFsooq6admgLgr0/4AuDj
iVGy6bwAxsAMGuQvRHGie6clHju1klcoIX37axqaj+ps8N4zOkeKxed5+1zp7hFN
grnoPZ5W6CqmfS1DuOZbQnhQyx2vYwG7nlaKB3E78hL3V10sq5dPzGcgFcIl+zTi
LMg2Iz+yirAFq/nEj1Xy8XdZaWOP7ss7c3d8u84Rd3m+THvsYsC/J8QLNNN456bP
Roc5zkkIxOLnM9FSp3FUEdrHdrb4/ERRQeSfFpDHPV47if301ht3H6rh29ag0RIg
cvt6u06AxaK4FFLppx0pBfoJaYY1CJxpsYSsIu+EpR2gJ8jTZEt6GPOxMGEcxk3W
QU4duHDQi7CnzrfmVCy/mGDxAqPsHYQ/XYx7/sLAVFhZ4iMD+scA3JEORyGFXNxj
oaFgjl9zLSYhbB+f52jke2Vt86fUzArfTyOjWimGT43EFIdHB3VdTuV3foiLMxFA
NUIC46te7Ode/zmtf7jvWsqfqI2NKUjXbb1i1gUFcAbr1QMQkksIFv7CO1cTl8XJ
aZryc8W8dheJ8FW0spSrQ8AW50T9yQTE7+xfUwIDDXiZjiVjomr/nVnczAlzNvrX
X+LX4D/fplY7igOhv8T5gEI8Uk1t+bxzSFD6h0Q5x9qJ1bFXu30LnuxMkTXtGyjS
+PlGNtT0WnTUoSZ+RUr2Fv1hSk+8JQZYUSP3FctqLDhV13dHJEoMSIPIJoQvuXCE
1i2i3ku3jX7UIqgxQZqRHdYqKq9aEBIJ6X61VBgHTLXAfypkWkTpK5KpPd/DFEK4
eSXeUHzsQYQ6BW77v8BNYcQ9ttPd2x/NYC2E7kVDSomJRY1D6HRne2+M8sOcQG9A
qyUFoOK0ssMaWn7gV2QS0Gf8D3lMTAgkHiHzsWgNqha0xHyIJuua8lB4n/CrF3o8
xz4AQZ+qBJZW0roX//5qCz8x7jxcuCkOM7j4v0SefzQU/xZakh5XWIMlruQjdhxi
F18Nc1YEQaKhRvZjaheymMAdawTb3pDNPuapJUC+JPcFzDxkEgloITVYVlfp/NXu
991rOfUR9hRp763HQE4b5/7YzvQ53WY+ftNdsfH7J0GNmjU7MHQdXkPO5IgbJsnc
Sli9PkOv6M7S1zISjZ23dw+sycWcFZv+XDVT7a1Y4nU1gX39Wt7YF19zpgGvLJcQ
WPFP1EYKeRNZ7iyINB1SsrhnHcwFatffyqhPdL4xdzQ8RwMWTk0I7HYYSzncraQu
woyOMokeJgdacejwLKD3T7+Vh/DYwiGhrjosgI1lQMCd52H+7vkWyV6cz1MVoP/i
3YKj33gNlgCtx0Q40Vq1ny5mfwc8DnrRT95gQ06w4v+/v+vkEReNrNl7Bwamm8oW
alcHwcA/mUU37K5EHSeJXEbi9lQwE0BJFraaTfN9D91BDA4ZGtOtkW4QA7r7xZaA
EZjNlwSK0P6NqnIA5eH09mu+cPPdEocQF3Bf/QBP9gEjbCrqJCC7o6KuNHdBOkQM
orKy3el5vUvDbvNDPmR1W37e3puMeKNz04GUKRICcPQ4IuKLrVf0sytnNFtMj8h2
96JdqO/QRp73m3JZd6/rDbmR/5rN+vBH6qxXFlUhulTTEXyih7ARs5ScnkqYDeTU
viHc5VNX5KJiJ11WHLmDo4RzjCvFWQvrAXQtnbBZ31I/yczG5gvdIv0Txd7CEvOw
QYY68riOq/fy20i/ejUKBc1aH7ds2LVKuAXeQcM14k7bQOIyCdcaZYAcwV6On8SJ
JfwM4diSrhp4rS4BYRS8coo6pCkdlT2odDMm8mep7tdQb5VZrVa+prdvoN9h2gA0
o6ycDShzaKdWov4JnNJj5WbQlZKepI4e5kQyxA0+CrZTgMRirYxqTqJgZvWKi62c
jlBVSBuqazjLw1fvyqoAS0W4EOkpYTve55bza9JGMB6/5EnJZ65treIOpFTDcvG4
ryk6oLcpB2TyRQRutzV44y+MD5hUDcg4lpZQq2GpfEnIRsRm5TaQfmG7uDpVjh1c
MNhR12ldcrXCDTMSGEVWAZ9lvYDCwAvrINnBPvaNUuKpqUybfE9SL2VxnVEQ+e6/
8jEkvv5yP+UgjJcAW4mC3v0Hg2rjuLItTevUHgS/R04NkNeuwTujkdXBfwt8oNCq
ihE7UeyJqbkMoR5oB7RpFHBb3oVGvzVMUW619y/lhzKgqY2s9Jw8szhh78djAJGm
kH6Yic9j3SrlE+53DNM0YeuaAesrbfpwfBZOHb5+ohtPloV0kuTEQjZpce2yH72I
MUwVXllj0sP/ZxNcJI6JL7NGDh4M/tf9ZC+ui0d94a9T60VoSX2/QsGqXigEOzZD
xZGKjwwhxYl9DqFG9YNXC6xvAZXW1WAX6/HbM5anWGWbLwaE4A/J1dbxjbsr/lmf
x9c4/rY2E2ULebgkRtTPYVZu+NpaOiTPe2GE/yuvRW5+izsMVa+d2sUGpLcfWjej
b/DJauwLvwXNPOODRqab0LQ1I/dYopHTZuJqJxemz7c5gF06ocdSus/WP+KB/0Bc
RZmBVLGjtY7zNBDWszLS/y1gGmeFo6G5Vdx7E8I65l4e+7z53u8i/pl/MOD7mYZW
8+lGRBEwJ+nIV5HBzpC+FNsgryu+8IBIAxg9tGFH+vVSw/st7leeeE0sNK1XE6Eo
aWcyqwKP3n2fiOg3IWHdweHA0WIwcjVWRfKE0+2kADyOeJkI0BxSB512DT07nlXk
U/yIrsd3koyMtgifosFRXF+r5G8lPx+WKvVu1Zb2LpfYL5eaCy9Aou8qgbG0VyU4
MbdXeLdHLfLLjk6a/hisZ9/+AsQEIR0QxZ0mHGCwcdl27d5OGDFPk44bTJI/eDdR
MMkcwrEg8GTSvpt7vQEtFLFIB204p2LMEnEO0tOLEgeSATaQat+TY8fIcC/WoR+D
G0MPAupdJ0x2svXePtxkgzVVdUMgl9as0OVFNB1C4NFoOfgRJmEOLw3oiWAbT0fS
zVy+4ksOIQH3p6phRNe0+m0ebzsqCm7HfT9lpSidCzmDGjUrybHPV2FD4qaPRbyE
fGQZkI38DRCJIIyCuKntRxXpJEqdbi/bySyt+LheHktpw61xwMEWsKiRnXwyrxTd
Ww5fctQUHvp+JTi7/hnvVGGHQ5X/CbaHLqhv/59d0xlnmgSHRkVLcQVu023Nz1my
nvdSRK4qYtbQBBUiiIphWKYti/B6O+FjWEY+/jWfk4qDr0RrFXDHQDWoyYTEwR+U
R3PEd9sMwL1eftEvjOhlJiChXApQPa2YBt1g5TJzQK6Pie0JZeIZSvJvXkS6dXvI
2vOy/UoW7cuZAuKBTCWyMY7BTHsyTHfcxowRNIdGfrtGxGOxduKfGabN2KMdFBTE
MnhV0tn7bQd16MVBpol5XFf26HZv5pBymlkWldf4kUc9lj3gZjpnwGy5QHqaSkJb
29I+xL1XN40c9yux+6s5Di2W52kzjJKg0AOQDKig8epZ6IK4+kcm71SwktvvROf7
jxJb7lmxMvBE08RbuZf5+jAHbM0a/zeqrCtuOrQrgobwx5Buxl0G6zG2G/d3RI9w
NVWE0S496zdOoN8KkuwVUQzI2yyRLVGJFZy9wWAve+c8BX/PpmzOlRDmH/hrpgVh
rkiP5UCY6ll7l12gwfLy44tQvE+Y5IwGhL79M7WOuDHiYikOhzXJIVDTckqwYqfn
XhS0pHCOQ9EB50M4gD4HBZO4Ej+Ds7sn2sISgy78az0bCEOisXiiEY4j/V0Cz499
DBkEpK0h4rGOU6patC6TbXsgoVs+NP8xXNxd2IapZoLR1rw/D1uZvbjjvpIoRUO9
ldklWEn6AK+LOUHsiIguebnR9UiWKTxhZ83B15V2TDiQFcgfHXRNFJnf1J0QXarz
iPX2WsfgxD633uWFFpeHb6Z+mW4BHVjqR7eUoov4Y/wA1wbStg2Khthyn8Ehc/Vq
cmcPR9rPGgwDo2nfEVXiGhlsV4IpfNSWYw+4Cl5WWdx5488MsOZqk44kderxWiZz
ACBC9TAEsDAxD8r8Gk7Er9NZOXz7Gm5TDc7XG3XJBZRAMT4qlWM/mk3ZDMkis+tN
t9fCoCwnjouF/xZ69f2jHk74WWjoNk3E+Q07JRcKYl4jmFK63mjNm2KgPF6v6eGI
/vFB1FK8pRyf3QY2EirynxU+9icCzaJ3VrA7OlrrZbzHTj+WTJL2Wqb446o6cFTk
2jA70a7476ZpnOhCOzMvsn1ZpwZkj3mv89nVi4qX7P6lxxI61hDhA9BFd2ROiA2y
edtj9Z5LujMlfRQxoL1bFqkftAm8quoCh+5GzPFDi62cPxV9yoDJv4VZ7WeU95EX
yQxQxRXP8+g50d+azYonBuvVXc0LI91nja8QzAT8eYIthSqui/QgW37ocSqpLu1I
mJjEKBoRvdBZCzyhmkft/6YsDVbzCqUwmHQMTD8dHvpCLWd3r5ECLJa3sDTmu4LO
MQFo4XXvwlWaFwGpbD8UFIL3j7BBKDFNCN41//gWQ6kVxJaSQiMaUy4YIIYraG6X
BO92+J63oYYZr2wGky2r3emfnTP0znGKUVAfa3AysCn8KEo+hM0H8/2iB3kQN92D
uTGb+k11KjHdBcyw+qZxIVRmuiYU/ZwBn3qYWeKdYoDu3QxRTNmxS/X/KxJiQTEN
mgUCvI2AmSA3RwocQHiiILY4fGwUuK2+L4RctOLqNN8u7+Dg23Cu97AsLvrAGygl
VEQJAWth58bC518is2+AvvRJqZK/pPp0o+dONkSQBAGTfaCmTehF3mzjZ9S3l2fY
gz5e7sW2kKttKC2d8+9Mo+TnoyO4sya3t2eU5R2uuXUqd6NP25Jm37XaYudR93rm
+1WSGt4z07UyJhWdPjbQoz9EJ53myPXYB67+w/K7RRLZxDBzA+GWxQBKeygyjS63
crEd41RwOEZFXjNjH8P5XsfjcUdRkmzbNEjDr2BiS8x8g3DIuP1dJW3+Jc/yj3jb
9G/xU2c4MoahUhuyxsNbG5lrawq3gsKxL7b8waxxhfaaVQRtO23b3dqclyJgo1p7
aYRJdB5QUsVj14fR0HC8OF9uWO8/z5bBD3U22ch7wUscAvhvKD3zWHhP8OJhr5Vm
zsy7Uz+B5ZWXZDhmYfWkrtONp4L8nq+9QX2T8L4cNtZZR0unXaam/5fC6zBOKG4F
wEHC6yhh2KUpwO5T+s4NXmvT1l2QYeDSC3r9XAZQ2zy8H4v6NSabugRN9WJOPoW0
x5ZZtBkEalNjciiaGnzLBVr9TeQJbi5E1RUvv7dkTlX0cdQObqeIpp+gh54rgZb4
3wxwwpOxI3gPV0jVwagpjxOYzr88ZebOAlqZMUbE2oJ2yUCOwqQHEo4Q05xVxVVZ
hr5TIO4xx1sFXuJPeA+x8s+GGX4zKiOXgLQJt/i7VIqAp8jn01oZ1XQXB7g1vhxb
lxwCbR3z1DQdEzGQOHbHeZDqRYmMtuunQCU4CNtapiWl8EsA1DByXWdIMqq7YFdd
ZYKd1bJ02jdIe9cvoOS1kmsyvTllkJiZzq4c05SGsbFSfO1CrL+cpBnPL1j7EWC5
+QG13BhM4L3cKpBwsEB3dY3wYphQAaNn8WLeHDj8RiHPXp8oPLel6c90W9nJK1r5
QwPWq2ctHewdNK9BrPySgT29yqfbk+XMeKXY4UrFCY5KggHsKOkLdaMMJgKDK1YZ
v/3+Nlsdj2lxE4SKV3nN+X0xZqANjKKPMUa8OS+pL3Olt8M0ULdOpoTJGjl7CDay
t27i8guxARCIA4iVQkiwxMC+4q5ToLHRQI+wj4f1iMoBlbszTvF0YQyov4ODa8X7
geNb/QDS+4J4VqqQpdFiVqo6FbIP7AK3YoQ7zlHjYCYZuZZfe87vJpSHe+IsYDCz
zLAUX2JwNktvhqlJXfI1E+WW9R0ve7vS46Z3/crenXxZ0gXPnpGgymBgTqC0Cw39
mlNfSjCKI7xWp3PEDKXW26Q/B3PgulYP6mnrCVncy89HdShC3ypM+6thBTxeEUIN
XSjNKQp0WizPhkCWydvarGXWcPlThzq8EXmrVYmYb6LB+5aZzYxfnhjJmS9HqUgs
R4Nwlw5WHScRWlTU0SziSS4Kf4ohZ2DCal4RBPDuXkk5UBBE50/1VYycEgxyyJg3
sfBpJqxcAE1C4ld641C74sa/Kvtvld1BloJ5bRKw87EBvIKEdNacjdpUOOjr3Yfo
iYbV0WTJ/sWLxArRk9KXjPranlsqcITEAczmg1UklNA7d+pyLWOap5ukoKnUdjeb
vD9kKc3yEUWm8HmsjBxhy6ekFSsEwEBsOuG2oejiTWzjWaRD9JkJ1XpY8o120ALk
2HtnZR6/OSFHgTHkS5qnTDZvZA2stiFKeSewWlvJzqEaWGeKBLuldy0EKo+PMnLA
jzr2+eAEgn2ExczJgGTyvQS3LzOpyqCh0nXodEXBo21nuvNOVOcaS1QkucQCawRO
7J6gRpOXI2eOp5cBRzjpK1hYiiHvjMZb/FAspYIV0302hht8QISttfU0uEyUiVFK
Zr+5ox6D7/fZoqS7175xbM9M+JuVZrluKQw3AFULFckDVNL18l9DhNeQMeb+nqBh
ki7+Hc4XXiEPt21iPVnKqg8Aq9Tx9jxsm6dgetS1+BSs8ACQx1rxXC8h65AiEjAd
S5/C9EnLRfpN0s+AEivKcze4UO3ScNjkCqw0h4fNXOiz/Y5U+arRBHWccRlah+5h
TvxTRLzwpuBr6tnSpaTXXJNVdMnidvxqITWhkMNEreUm1pi/AkpAyC2IQmUKHRIc
NpsRq4HoFa1p/KCHwmyEU1dbZjGhLJLhaTnt6HO1unRqYU2PJlypHzzFd5z8euDW
dHNiyqAavUqrU7Tm+YCoSHKo9zlgkaJhbRnpn9acKHkP7MU49sxj8TfpWs4VXkeA
Xu5VW3j1s1EYgiLERSrrD5EQY9XjSFLN86CJQiftWwNkiWvQe5TZ909lgwlJ+gxP
UJwvy/tBxBJ02b8MePmxkpyXl/zVTOhR/PVXDEfD4jqES/szWy6mBxoJprVW46kX
rHhAbW/6Yqu53tH/11UfullGw0lIg3X5wnZfdzmoB+nnmEXJGdGb/7p/7tC03ecL
xnZFAS5AV7UndtMUjJG4aMWXOrgeZoGRxU4Blphl6Udt7M8xe/M3UQypsXa0v/ql
Mj/5sw9Npgr2gtm7xY92ScVLRkxn6lagT7VyAfwx9EDbJhi6xHwlTjBAwuK/jX5k
p4E68bbVKlsWKWY/akINjCx4rFxaFtPg0w3hH0+PgKmg7mVjjrYuhfQ1+cw9AEpz
324hjRBnZYmpY24meIanswYb6g949UdcnML8Adyl8xlpuGYOrFutwQlRB93cdPIh
DK6TZo8TwNwtmqnktmqOqZU812wS2NqTuDdp42jm9evnB2cot5NhneO/KBCcVUK/
I6X4zh5L7Mkc9PzbryiN2ggjpIcrgKrsLFk3fceY+1hSOY9fIWYdjA1cMPplC1x+
rODKeQs4kXbJqNdY/7ySAiW3hj7Ae71Gcc459x26hcVaDE3v/91pTL0WsDpqMIem
1SYp2RMgdss3PP3mYIVzrdRf05idGz+oReFzisJtqpPqpI7yCCmwadcos51dBH5Q
L73bIoVFH3ZY+YHsxRLBVRI1TaCECGkjCohI/Lh//MjphtqqAXx3MxxYWicAoDZX
uJmR0Oc34KV8qU7pwq7NGQAvu2vEQ/IwjcDMemeWmvp8kmRvGKBI6HF+E7K/Vg1Z
nKySftFh8VUlEynpjdhP1gdBJyZCk1MxwSse+uohJSrv1Z2rja26pB0w6Oii22Cu
cp4uk0Ijvwl6MhCEGtAnADq12r3l+/J10HoOJyD1rPgcrWc9POwCIg0H8dipLVJH
ADo5IRwiBx+CuAsD8sDZBD8NTtB3kaZPifvAA1BHC9L3aM37PPI9Iu7F6Mv/glPh
AcCgrmONNW3EyuhAzHg3k8UvKh5Mu0N3HAaVbda3vfN3xWfr5lnJQ6tFKcgqvMEX
xq7ET2c8xyGfHhmClCXvgZbuJFH9W5pHKj707Cw9nR3q18vktmnh23JjGvaALdzf
ejPdp+jDtw8guzTJ4LajaXggaGUMYAgPXbWcPYjoDOhwO2J2P/LGIu6UzYlxa5AQ
80IiczJ715W5euvJtpcPrnFfUZ/uTHQQPBl92zUQbZe6YxpQOlHxxmg9ViNGrXR8
gyBOv8obvs1a+06LmyCk6835MyT4cL8s0h+RiEojEy3IqQ+s4F0nUulvp1TGXgC/
zo/ac4aSfaE76mVswFWtwspWkx+yHCBo1adQyDivJdpPmEXKLt1OxZGwE30p7v6Z
iOgrxkVxCqDzD9ByjN8xepDwEKtoHD6NekObcnTQlD01xAMn4qpbefZr7W+aLPv2
WatWUcj3dywlvoMKdnzWh28NFXSxZWDEI3FqZ4JSb/oCp55+D0/xK8SN6OUaL2EH
gdKyNILhlWHzqarAR9JRaBoOdRPK91hCCUkPMgMm34Jj3JaSAtMwiKo+AME0SorR
K1IZT+knMSJ6SpEFQ5nVJ/mTLluCIYU3qtQd9yUOZZIJq0eLe0lgZObrB8qA65K+
s7sqq+R9ZJI9wkMnlh4OJ21ZP7wATSnTwPY0AX0GHs0c00sbEKf46orjZIxnPkZk
nVs3SJAElmElcCVEND9hRiqp/aqbLyAY54vuEXhekmNKzdpoxbmQdQGncCawTQEN
BFUfX+2U9ts2B688yK+GagOTuHdBqexyX9PFhz504tJ12TPKVxanwAN2v1bdekRE
qjikjU9bifKAhQ5a2VXREilmDH/uaKzefEydFTbudHpbb7WLEdXdFDCpRXrlYliM
TR9vuPXQ3Ire9G6zLnzI1wu8RilBApyFj6zeasqsAnmFcGggNHwq/5KUB4ABJTZe
zBizbEyncg8rvGRlXcAS3o2d9nrBj9BYVTXcUKCZ4TfrWGhefFSVByC1nL4jLp8I
Jdmd4DIJiWYbg7kUgP9KW8vgNRudQqf9b1YrLQQ0hagjo1kOvfx+tnq3znh13U/4
rTD7k+ySItKRu+HZw0a216Q0YiPRax3pKWmTNHhub/etEG6lFiJPArRl4/41tp1y
o0ce/7kgBoem2kmR4M8I3sm1Hbz+1megFSuxjUbRqX0N8SK7/2qQJZV261Qyqp6H
wFhwhNjQ20mK5psDPJY6o6F5kOGs4iUA2F5JfXVdCxlxoAVJQg1vwbUcqvM96AiZ
3xKGCG+8nPDPJGOAokt5GNaoOSQL2Q4N/JlJAenEaUEwxwTuTvqO6/YSjNIC/vld
uc/cMvrtf31zPJuqSZaJd1BEp5GMVFGaQl8D8EhBRwh7S1vUHt2pkqtqkxmus8mr
Yen1ynJx4k29+YdUFwc0bc0xlrmdjCOrfL1m12w7CvNXQL7KuAXmKQ9XykHGaAMr
SyF+/pKyCZhPPIxIHn7iI3c0cKuqQYDlxrC3+SE9KvyggVAxr5TsBowLP4qMVBBK
a9rCfbfjtFA5WM6Ir1aRhG1pCiFgtaXdzzV07JkExo9UD+zPF9TTrbfjFb9L/tOF
JyYx1FsFIlF0FF1+sOW2XzcC762ywnZZGtsDrzXVIHurgl9Oj+wHUAkB3P5tuMqb
yY7+mIV0nr9VfhZFI6UCtPhoS6PPpcQxCQXQGmbE9FeH0KuGBiUAS0XOOc35XESi
Aew2eUc9Pw7tUhAxTlQOqc2cIUKfg9aA+R09NXEV+TXWcbyQuLc37MX0ZaeUotKg
IyquycFP21ztSwfAXkcbibOZxqtrpThmJxWc6fB+bJsPUiKP7pQF1OMjKjzrJ7zc
Bzz+/shA9kDbTZZCd3gLOqFDO44vax0dssLPYyT4Kp7GXPJTMLA43M1Rvj0MNEnt
8fPRvgLqYmO67ye/4c6pgMp4zULdMjwp4JRL/MSRjL1WlVfkd7vyiDrfsnxHspZb
smGbEcUkr6HArXcLqYGK+7xi3eFhlMEycPJ3sT3+RZHJPpO9vF5LtEkjbREkMe0x
n6m6KTjWpDGI4x6etrk97+xCGN5PBjz1FhqXknJb48mK57zPbZJbYyOroAvjTRub
oX0BkuPvgym4NIHQZgXP7SOn5L2o330dIve07UevlmATI80SXqHvFGVuRW3/8LTI
2D/T8tWUpPlezOnG5R9VcKwzsmCXIf6W8ZYZnSn298GrAQkzu+kCkLlW3WKzEnd6
m020yTM8blwCRPe6RHHtzouNfguGxGdiEcwQ83Twk5nau8UKysUHu0BmTakrjgH9
d604siUx7SGCtFQk5GGcZxeommNC7JVutE0AiHdE6n3aoP+W8MZ8I0Nx8o3A39UO
zvYmq3mooaooVo7ydwE5iV6L+Fgpwcc0m+kaLQ/B7nnpTCRixOYRHhQr8B04Ym6t
RDbzUes5ID2NniCJYfQI5vP3LaZ9fQh4hT1naAERw7/cTjYy+kt1Nwa7MQJ4IMQl
2/rHZ+Et/qmJvEwwuCWZGUl+VNiEtRM2ZSrLI0tEYPMFPKMWvXx8IcYkIJeSunwN
k/4a4Gf8n5fV8xx4HvcMtLQWRVmvu5lq1UM4SuD6Pg8QdfhuFnFWXIScZjmk/Mfr
1/XVJyEfOraoz2VSWCl3VdcGCvuCHV7fNw6csnyOyAP23GQYtakbXgDBnsAKp1pc
yUt1QgmoQ7rjKMQi0sQA3/Tatc+JS0pGd5sO9Yngna3eXd7hgo11oyxJz0l0HHBs
aDZJVWCXlwzZyXq0XS0U+HM2ohaeRVjZOtD2KpkVazmspq7psZhsjlDrKx7MlnmV
Xws1nyKGJ+OYi9MHfhvAlsJseogdiNZVCpSkPfqqRhv/AdCe0LoQCyBpaDAXcYni
CjQQKqxxGBi3ajL2LCUxWMquXSV0l3BwF23b5biqo8bRm/8Uw2yklr7BFLtGgmFC
X7rZH+QTjjODU0xhXJp7xIPHG0Lejf1yCTFoIDvFwAqPO2I0f4HqsQR+HGaQILAF
3P5jL7gpOb0IZUAgEQ1i/YyS/fek++LycNX1rRe+I0wDSqqEx1adzWQsDIHRi4qH
lgQ20nfQSUA5nuoavKMEQGmReXgh2QCmr8+PyOzzpBPicSJdYpzGXlCOR/K27k6q
4Z8OfNh5jWq0A3jcd+AkL6Ktc1yM/ZuJQ3VRAzL+BSg+MtHMd4O2lJkDKXZoMhPW
edI9xxYiPVNXRZshLZIZGdxCgDut1RrswbfkqODnwTPZB58opgs8mIausGPST5Y2
vWYCB1dJbJGf1f1AUx5gDiZdib+WmSr4damEMJabKrbJ/loFxEhOi7Ej0saticdw
AjVQeCR+oiRFjwreHYVvy2goxo6G//OSOHVaD0BbbzaNJhy/mrK+xM+0/s5pIq7I
W2e6InIN1UuO8UHrbdZWmOqO5nn8iM8cc1q0i1wmKAhpXeNqGkwuJa0CqiVKaemr
P9khttQxIGBUjj+7LFV+6NfmJXPHmkIwSFQ0UkSlroGHQ0kmxAxsqq982+chr1pt
HZ/nWszEPa0uwmUGqBe9jsJvc0eoaQe76DhBBcagQfNPFiHgH8cEWPMaJpyudNlX
5eRT260WaRSMyAYUJBqIV/sIo8z8WTEN8FzTbEATCLmx76+OXR26sgvakEdNSXxQ
3aPl/68eKzMy0l6EwexXvOpEk1iLFTDXwRya3azyX96xgE3KEeJTAj2ajyUqGFRA
fEgmrhqXKFt+TG4k8ifjYDv0rAFulgzF4iceYs4c6/PJlkcXebAYd2R02wPrHASx
wvV//NdHLf4qgtMTsuTmW7V997tUlgaE8oADhbL81lB5rd3HAQxHyWZXVDBzfBsS
+SNXB2rzuBwJ5h3qGUQ32rEfmnnVxj4c6Gsb+mpyzcwo1WylEwQ40aBsgV3zVRpG
IbgT4mmqlFnhrYniQD9IBv/lhRpB5D3eqlAjq2avS6eACoklBbUhNxp9VC96h1cg
G6OrHX2DoKNyf7OK650ViL8QWgBmNPIQqOG24VQL52te3DWNkVHh5/WMarrrsOzn
/yL041HaDfuwpjEdy93Z55cdWH7WMTdizzg6S6Zdj59fMCACySFjBqd1z89XiTxg
2ivNLEvjOba4hP/W6swY4NUC7UyZpd5jSV3eVkXXTeFrJVBGT1kdvhzGGeVC7yVY
17SDlIR9WzFZvr83foh9em67wTtxzpp1J/K5Bl9dc0B9/Y+vQTEpJLtJ5B+/TUqa
M21PLsCgn1G+TiirjR9KuUeJW9m2FV3VSgxiWyrBc0vbCWBeCLMP4NjX0SIGFtXY
yDc0x4GdcoiRPHsawqASYP/sb7ER5GOTnlVN6OVAD2ychPR5iX212LFU6r3Cd433
KcSyjhV9we4jDl/wgV7/euIkzxGU7nC3/QSQz6I+65OV1xadLbQ7u6uXd9iXTeZw
+Ckm6GALfZGMcV/noweHbZ1Thfee5bmqrPjJVQZoW6dV1B4u8NhvKtIaJpAt6lWG
uGgOtFWCHnjZANuisICxBJmNHX5nEiPQrQoSBG8etzt/zpL85VayE3MYOCSZ/Mol
MBV4P7jfltxzfpVwN0bXZeGWT6WZT06hyCuQTQCnKrTwlhtaSd854tVsNpqqZmgv
k053BVR6cEeUjYgJIeRlwhieI6g0M46j1wPEdESvirKHQ3XboZ03qB5yzOvXjHY8
P47hs8UgLxP/BNM7o4vy8/v/bHdJKdo20cbqkb8XuFQpfoH0ukY5uQ6N/NkgRLjv
Sm/YdVJri/JnjzluOhujNQZ+qTPKIAW1SxriliCfFsrzttaha9VwDLN9jglMJLwG
hzJrtwO9jiKdYHOe5C+ycR/6WXLg2VNaigbBRo5Mwxt88Plho9r/1rtKF6ayU7W2
b41G25qmCVYGUDGqfMAxwerAlyBGg3huk1zz7nwv4jfDb/UHPLrgH4SX6mS0WLSI
CWO//BvNHTfQ+0qKIxd0xEYfT3wItPKqGa2lGEvq8qWgpn9BLMrpoHI46ICRfs5U
7JBdzHKDI+r2cOvwFYSV+aFArq5Yx4x4eS/0M7NOtl8pjpimIXFTsEkOHJ6nEcc2
vvvJMeXPNLoeen96r+4QjwqNejBEqBJsijVt3ilWKt0X+DIMHIjwPGg7oWeZKEBu
8lSdsS38rFVNU8Xh2eCQjr+tPay4kO5VwF1bbpF2+a5Uz/yk9wqEI9wkkxO2L3nF
SDE3b4ZISnY7vYK0gMdYOth4iC5M89BoaHr2DzCcZ+sHJcpB4Zeb7zw/UwSFjX8c
LJSOSbRin27h94z0bg7V8Glb7+x212yUhQ045RqRUeeIVyNcO4m6X6Eq2BlM2QbA
leRViLsruO8kA4mAC/Kjky6W2kRm6uXBrTGlzTlwMk4aBinYVwY12KnrJ8ad853H
ZHCghwN698W4NFWUyInp+n2JyJf/3mYtBhdV1Oee7fso7zX4mjLYAol0o1PDr/M9
UqgnZJ3GrBx0cWwRJuUK3WXty4ghKmdZArnVt/OOR+ka8kpnngKGugMe84Dmq28n
VACrRThs5a7yyXISoGbSKBdcvc/ePM33j4PnYWZ1PnbfrDfw+ROcuFLS8li/FohW
r6T9zf4oR35wCkrPgz/PH5wkKQQ3P4vZXridli6g7YYTzejDWFU+znidLX7Hx99h
jjo4Q33DD/KoerILzMLuV0GAJiLV5AuFwd3ET09BMO0PEQU8bNUtoiinQ/5Va9gh
pbK+m8/mSGztoEA1sKipYm1fJtTq51aaDiYeOKDkYdF5zNfqhMSnPoY075JcFxWA
VtwNexN0/en2geSJg0jtMVi8IBWWMbTueGNYOY5HgPPidzJT3PB1D4Y2KPY9SJD8
PYxtENk4YUyTopmRj+vA927aJHezHGI4s2z8jXc7IYEihRe+H40GAJ0eKkz78AAO
ZdicPnloxHvJ1PmVImE8sedfEkmHRib3RNYL3z4FqM69QFxRwGW9x+coWuLIfBnB
Ew1Ig6db0JjUXeRSw+4d7iiz5aGLsUn5o+g2a6O8kBRRIUbu44SKz+U1ORxVP9MU
XThzRzXOQ1mQ9lmdV/E15neu5hVKcJwlU1Uza+6XI6Q2kDgpZxw7QK4TaRvwgQL9
M0Oouq+iKcgmRkDyVG5mXClgn6WML0yvz+fsbKvpNzDkF9voMxPLecbZbvuiLp7j
BSGOyfQf0VR1ExkmWvEbp1x5e4m4rAmaAiNkzo0kIq2oUTPJY2opqrR6ccOAlp3u
5k6tyn2Uw1Ew3eOSzKDTBp3g1YTGBirinYjSXxcJrunrDjyhf5Q8obx6QUsePhb/
tP4xvGX0/lAVklO9bM0NFUvOkTo2h2p52jFtYqKQwQXU1oc2Liy5rNHuaPw0ISPf
tTxq4M0B+0qHvxLrWS+nipZ04BSZaArmlmhbJKqw07LPQbp4cKhzfacYGu7ntEGM
EQev510co88cvNfQxL9ahSUyMPG9VFJJx23o0CG2rfYlCnFrwpnSOgBImX3TmkFo
+4e82X533/6zRYSmfUvuPFW5LQ0qmm+lhDG4BAOjRoZtsAAuIsXk06tVTUHbymCl
rStUnbtiQZDiuOCsjRpW/4VLOBHMIMk5weIj6SKEYdYY8OvI0eDX4AKW5QdLMp4I
EY11edqSZbzo+iyyE7Oa9nek1uwh0+HmiELLa+9L5T/6K04JvbhaF5dRT/i7ERBd
4mF0ICeGqPxiX5sJK0CUWcqoTXdm1WQ/5KnBEBGNtZYL1RMJLfYwycKlRtievyEn
rxn3+rxFAW6UcthFyCnjqN8UGkPWeea420BVkr4T2uWvnLY2WAc83HxxLGjKCYS8
5Cs50ADAUm9MOiFFBkl7xhJs9qSbW2uPQDNlJc4EDiTD6XsB/5kX/+0vDyphwAz6
WjleLLVe4R40IvWtuRsw2gubunMxVPzCq5xG06p0WzE7/Ji/zA2otaHiyyffALpY
61u/9cffb0sn6f2X2uiRbjUDKNRz1e4DR4VMD6eUnPm1pnK0cxa48XelaJ2ilmYJ
u7/QNHelmPpqKMuaL/Yf96c7ocgJHOP3QZ/bHAyyc61ydTEtaI5UxpJatEN1kXth
pAhaR6PAAYE/ztAQTfC6UfYeV+wQ/Ds2RaFaIvNKF+HHeLYxHPL3wc0UlNAPxzTR
k6jVZ42oYk4aljbzckUyqzW8vqhF7nDHRyyHuqIZBoq+v9dmLTLZLDY2q5ZktAwz
jfVaolIHB80l9mQjJ5radSkaGJzU+zmhKx+s10Wf8rhMd3eA9XC9Hbx1gGwSZhFu
Q5ls7oaKw5quzmjdFu15eqVi1uNqmBza4JqvJcDa1vxsWweUIN+fWI+VbDgzPaIl
e5HVzMp9WVc6MIBCe7PsdR54vjXeIXYNrgY2JR3LTuvPNCmkvyqABFcfWyVjQDdy
YzljHnGwa60tKMHPvmzFoteTQA9UZjMu2fBCifwaPx3nTiKMJEuEP4uYzfT70FBA
f16xCACCNjqDkxHrllPtU8ajoNVQGYoBsN3/6mvuth9lUMd7yMMnQf6RFIhYpZ6n
vsEWmdJsyuEprKIaE0xmsitbQie7/7uHuEGyptkkr/YN1fhsg+SWo0ZA35OO+bds
5rKoMhW5VOBC0SI2kj2SVYv7hdk8wTkuoB4u41JN08J6LFRM7x3sWZD59CByVP3a
Z0EhLK1a9kUYO6y6kqNFOTMxMNQvAkEHl1AcPW0d8sx17SBZtrRvVwPEPJNdM8pH
itjDT2rMtZHfv3NfBmhwrQvdMq+woAqC1QxvKphklyNw0klwhXGSrj+Uj5HI7QcZ
cYKup1yzuKeuu1LF/cH43Tz3XdyiGzvnSHWh+cRc2l3tSyA0tqaOUS3TflfdzF95
2CLHmdQNqE1OWDLxpdQwra4dQez8qDopC+wzyiNcYh0ZSqhUlW2c891xtCQa8PJw
V6ivhbwZwu6trT4IsIueQf7gmhME7BRLm888WrLWuPx9GB+ZS5HQ6tWzKsg6OhAQ
0c9uwOec5v5R7qggpKJhoOwg7WQwPRvRx+vEYBLbcrSzors8+vhBnZBDXThu5B1j
5+khuIJ4cH9U1CCloi/TyanRv40mj+wzB1AzXpHIb/sM/9bCBsT2XjS7TNhv8gig
LiKTNQcyDJllQuxyxJFabBCUT0fSv5cPCjUQqKQQThLdKEdZkLciVEK8Hf8CYW1y
zTaueVIAYwFN08/91lF5TEnlqGPoiw6qB+m7Xr71vB4m8viqn++lGpOW2csKKVeX
Ts8wDY6cwIxQn+kBNcBN8rDzwhSx+QyAsCQnZvkdUdqhGL5icJFwchl38yP/4hXu
bpJUBysXfdinUp7+yAv2PMlLB2Y4nziiv452OgRp+D+9V1PgdMyJet4KzH74MaD6
Ys+ODThXfUYLpokWgOoZqwFfuvUTTP9FOfNZdg4h+6C00Hca5LO/zjKDJ4beMGjj
A00ssiutvlsuPHP+BsVo2DHGvtIfj2uXb0OIyvW2XzthE1vnVuKmHBfk/l4MP1W3
/kW6fquYEe05tdU7gjCrPuvkhc1il2qSRFOGRZbOli7wJWqbp757Q+yoj6hvqs2X
WODsPfUQuKcOeUrQ6ZptgRUc6UyMF41a9/8iSAQzjqRjkX1gaLwRkwHOCAmv4tij
Q0BHStoug5Dc3w7+PUNKJBm2/tlbZKbJTtxrisrhvacD+ZT4j4JeQ6RgJ9RaEGSQ
IWJT3d3V7k67PTxjfiT5UUKcTz9bnSSKtWzWZJaXPIgTxt78w1oAaE39J7QceZcz
d0CO5PP+MKjaptenhghRaM9V89ygGA8pGcpsGdEWYFP3WlUZrjleMBHIKQg7ZyER
sxK0ZV0w1QIb9eCGNX9Ex0njKlPffQ1JZbqlCFiwyqR8KBJzCK73UF0KS9Rj9+lQ
a0Q1yoCT+VKOAMqCrrcA7BkdeIOWA4Jb1Cdse8LUsbKIibrqhoNS4ZLYQB4ka7Z8
Sxea8QO1U2gZewvXKTmifDjF0p+yAmVdwoOSR69zRzS3wOsRllplJ+O7bksLwI3h
FJ2pOvo8zeytNFIZtFZCjYZGR5ShdN8l6FUW9S2UOJusuOc5i2U+5Y/khH3yIYiF
dgrFrJy0TE5GmAtz6k0wSCIR23ZSVtDraCSkFMyntth4UQEx70ev51CkAtt+w6hu
TDK0LXQzannWuvq4jxQXaxTsTnlQH4exlLmudg/tvDSEcwfBVCQeWYPnzpqmf0Ex
2H0zLeKGKofOGlE9YEX+tKPySpneRGbx4jRAf2MTArtmilfD1VQJ0KhoQ6ue84fA
+huFB/ttEeQtfsQGCCqYEJFV5hKJn3ztAkWNJgiUXih/aDPO6B+V3CHqEPvPB+ca
wbJ7GjiVf9BTigvroDvg10lY3/fG7WzGPf3d+VNP7Uk0vpLHe+TRribD2ikVqQGA
GyaXaHnkk9t06Lha9ZaqNA16aX55lmcCruRdUaoyfpfPRjJ8CTjC3MVfgBJlN5IL
ew8B1eLY5yP84HY0LPt190VSHqy0z2hsReMk9bp4CZeJhrRQrXB9Pu5FwwADnQg9
ECAKwnAS+pi2Vv0IcuSODIehZ4iCX6RtRViDsNeSi3KfpBJzhA7xIiiZa+gYwV7H
WTWjikXemaMHN+6s7tnFcAix8/hdoAeDaz5b93KDFy9h9TEnyxcr5Nsa3TZMdx7O
81Ib5IT6HjmH22hvV0zh5dlsGtypc9jVb2qZmn3X+2byWo9M0Wku1Ey4tW5KDTMa
GU6ww8uG5TlNM6b8He8fdrQMqvnSg4QT+JbNFABH0D2HjkRxCYnwi4xO/PM2TjtC
FNzRtE59H7u5v+aq9HGVjgooECktvP/gAxrac6SdQdJ35c7G4XynlXBR7qH6P3/E
mpLRiL6E09FVjlSKuJtQTvWvo0B2TvZk/TL3mJSWn6NEywaE4RWS6GV+bpSlWWdc
OzEc3bBm0RoFN0wWWsIsCnGsnDIOkY5RNT2Q2MZHlBApmWMlNJdq51NOOuWYChsC
cVWqPMFGwRv3PRhgJ62bRQiiDD2222npNEVQso+HUaxqpcActyBpJwMjDfXQ2isQ
DGR1kTsA7wM6zXyY2J1g2WLLtwQl4FZ77p5ZbOo/pc6uCF/w3EHTwhaINIKqCY4P
4GxyCjt34f+JME3jKKUWsPuGNiRvqq0k1NuQ1NMQG16Dzx60Dg+2XL9uXui+a8bc
rA1TdoC6+/TvIhpPtE0hn0DbOGVJmxTrOlZ8uW9TBzZldb1Z6T7KNVfoQdrOtVtY
6dRca7h2i5SiE59igkiKkwkpBiKNz4oEqDVBsdGhSaa0pcsrVP5mGyyHTfgSn5N4
zODe2s5fEpj5tlJuB/39nXzEZoLlS7M5L5bdnAIV5Lf8ergBp+GhI7+fIQyAJXsY
Sa+vLBESbi+QTB0eoo8A/Okgc4bAukfMjdfd2qkJoV45ayD4/r+0gFUgrkOOzVsu
h/olsa6tzlrOpt2ipg9V1ywXBejEiIujNHE88658zDTI5TqOpesW2R/m5WMIT+Fe
syEHAi6oRO7PL4Vw+rp8cTheo5rh/5tWREH+uTy1W81NLNuynGGeC1Mmqz7iX7nX
eXMVCYyfthlM7JJXttA866FCJ/KBK9yEK09j/pQI63L0pE+KVFMib2tzYKtaMjwR
xjPEGXGG4fcd6JE3lwGAwFtVjJrh08413KczWswzBpUDMvtVhUp3u7gN77T4kzqz
s8tC8IKkkJGSDtwS9Jv6pOBhbIEn7KzAcMjsL4N/E06+JdUIkwbp6XmkdESxMY2q
2y096SD5uuwY4NAaiCoYDzMV2VsUS7Mxl8JPzqbeAqoo3GE51cdrnUm16XCUg79B
OmaoDU5K6cfH5BNnyMIr7cd127rFT/vXwlIk/5OTPl0KoYcd1gLRE3HCb027zG4c
9yv8V9kiib/FsCC0ulP5hZFUpxezLuuQQ74upuSsHhDDlFQST4iHXIsnNHze8LwW
vOmkvF+YdF/1VjbcbwRC4pVsWHtSOm5XcwSpe4YKr0u/W7Q9So7QfDFOYHV7nKIL
pMo9758F+fIDs0zvRLOyhFaHlxZ4xToHEEczW7ahSbEBKmF8GW5S2mYtI4MpHgpk
pTF4MbX4ZvdJUG4DIdSTVp/oqvEbdNocKU2zWDSX/O7mA0+Fhza6Vbtjc8OzuWj2
EbASYG3nxm0JZ93Ooil2zJLY7eVA63FHoof5sFTd8aLH0F6ir2F7mBiTNSODDHlS
q50X46OzMn6/Wc6ImDQ/aJXqrhnLFo+VIBetOTQs2Wl8ZS+ik7qASsP0mb7TnpWG
vBzZiQOpOyDxB/Nvk8TWSPUt9EDXfRAphIt+B9qGBEOAE3BU7ermfwkwOLMiyDc/
7hB6rwDS99oxqJqsZKdDSEo8NsDD1OGnx3r70euWHCRT5pLxx7kjsj9ExscjRv7x
gKuTCLmieGvbEKBDk1BKgvEEydNb5MiaP4uH1UXr5iVFeaU+3M2W9r2gQMkAZGeW
SqcTVyNspnj4jOk93nuH8DheCb2VHnMSDDgBeTG+VQy/BsLWDmJ3TF0K5ClKSWHu
rA/rDSKU68BqXGQzg52sQgBn7q0c+BwoThtFaEsv0tL66TUX4oqm9S/eS3FDO3Cc
Hu1LzwsTev9G7LTXckga9rawOEFZWRLAHAC8Lr5LxcGe3b1aUiEDVd8lPIBdS0rH
zPKm1h8tow3gzIfFwzbEsClZMkEhVJroAi8bI7n3rXf3n0+UNYZIkU0RiDsNSgN7
/oDy4cZnVW7M9Y//3jXv3wD4JQrmGM3BRVrwUtg1iSMt6nQHpXYoy2e4d+6W3lr6
i3aqpuuiEjh1rhcJbyxB7HmI/1vyiEeP4NbJLMUQ4YSi0UaA2qwYfZZVNA1lBdqC
zjfR789FS/L3wOQPYrLSz7ss6YupObLw4M55bHf3Imt/cEat/BBOGTEwz6zjZrkX
SBP71m1UpTykigiuVsAOQLlx6rOe8MJAC73YzF5+sgiLr4Q7UxP7uQXAAVdZEIhl
sjrKeapbboTZdy03NSKxrimVG0NAEC/8ncVmSes/NbY1/1Bj4IPOrL6OS/GvCfmU
yFuqx4trmwy3PEoEVFjwWKYcggFkO+cgyQ4xaXya9Nyb5BwOslu0RP7RTokYOlS9
J2JFM5GSraDMe+XosU/o/vUZEeBGagtL6OZOGt6/y77Euf6xOWBup7f6TNm7p6KH
kVrau8YHBMajCeHV60aJKwSlEcwBC9nAptvRpnSi57niErbAqGoFBHQdnJpyhiwg
NypooSYkmp0qt4n/zaLGDOVEmpS+avrXxnei6BEZqro2VbvI5oHKi7GMyLaZaJ8j
buvyVIRDcIaTwqhzOeID3+KMAnSljBct7l0dsOrRB0TYoviN4/+w/NfXPaTbq20b
i6DJ1qchU9LbtnFBxS18VeXr0w0LOwnJ/jUKQgSs/lW+ldNcfG0rUDeteC0nZxe/
6KNnqnNCNDSBpIiO6n769aE9uM4pxDIh4KfVwP6w4noocRMEOjmyffU+E0QTw4Sj
FkZYeq3Ic8xSM0Z3qSOpV/flIbpSSvhOBOjjpWDV06gOUc+ojhf2CzdIhj2yq3Gy
Ld30/MXnq1eh15rG130qgul8/PiZq4AjLQMr2ax1gAUalZ+Aea1nGqXyUeG2O67F
0KhC3gBp2K1Lpl6EU5qK857FZXLatzXlsWRi+jo7+6PeB8qzdjNFsXdKTacCbIGL
GE0ovyMcjpmh05jHjAbEVnZE3CKh1jq5bNweMVho7/NaVG5xqjgfmSys6Bvduc5w
LlNPDu073TXoColvpom6/8Ht/cZ2tCbb9t4yt9nAU7N+bo5EpVl1GBIEJlsgUTve
yMwrDM/UJLDW2WCYV/P24UYrYey9y7oPuH1qN/Sx7VfYlHBnvwOAARaz88+N+zaF
BJ92j71IIMZGs1+VfKiPTnKZgRr/o+46H8E1PBtbecyOIRHRJe10PotOgcrz2umd
vD4rTWsrunfyE97AcHkVKa6FNJf4PuwEgTzlyEhcWorsZjM3/psIZkilDhKY+J99
LxUmX0h9VHNFo2+e+O2UTNTJUveKsUnIFJX1dZDamYzYT/Hzl77rt0YaGuweov63
Ne6lFMgtNXWF14dXH6kTeTnndH5EnBazTM3obHyq8Go0bR840XIXp6kwzTSsWYec
CA0EfPUpFJPGXDttejgeohFdU7QebFYSEK0uYmIE5Cr+GZVmz4z27d+/DBedSP4Z
4sWQnziEHrMZ9UQ5npmM3lR1Qy7UrQZ6woAuxKrF1yCMuG+BGTJ8LQLZO1dyeL2R
zLCoCBEw/Td/GcGZOPY8bIxgSsN4i3BzCDVMFnmAkd7mSTseCoc7genq9dxukoLy
`protect end_protected