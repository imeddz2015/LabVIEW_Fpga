`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 11936 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/59UwEX+aE7FohaWu0/8IpTj7mav863zUNIsgIH2BWb
Abd9opeuBjbGF/waQMI2vMJTwD1ie1YueHc3nSNpEh4OXp8P5ybZFY89uyGz3ztU
W1EsuUnchJoQgbHZ/sLbgtGRgsrAFn+ZoIeGN1d6RAF2wAESJmYP8zw+p00RvjZ5
G2ATm2jrAjm+J6bPpiDE30wrwQaPq+vMMgMQAWb4Pqbixyi95aUvqHl3j1E84SCZ
BHib6GjysEhbl1e68p5n5eWhoXmZ7s7zP7Pda3stxFKy6jnKJ2srvmu2PzkkXsSW
Op0hgBSMmI761EQ8yd26fxD/xwvEnfQ37CBQSn8jFCtW5ElenCNGOqOa/7x8dHZ/
rbWPC+6tBQ64VCC3XTpU5uynk7hh8jG12EN9zITxKavQ99cZeWObnTQXsTXwEDHQ
q6NRZpK5I1hIicRlxjgDM1UlZhoNI5H3nRszePOGFvH0Cct3kiG0WoHvrNA1bm40
/kfNGU/P0ygZP/6JaLEDsVPVaOuX+0wLyW5aCOFBMlqaWzzLhSWaFoGpr1636Kcu
nhPpi6T1CMUF+H188iYQjnr5pu7ToCFcaC0W7jBsWFKaHA7egsWtlzbOZpdEXref
8rYT2o7wej/Ecw0auKFTEf12SrkGnLJvjpVkjlcPwHa23xUe0r84luTJKTU1G30k
Gtow3t+XR0sf3TXd/ogOES/O108G8mx5x9Cbxbv/myKt1C6NWLV36sk/Un1mk6St
ubVJMUPpRk2vH1alI3H/iadLw4eggXUELM3MMmCWmuh9j8vITYvbqdyFkRQ+nfc8
0TuE1kN4sH5zX6SK0yWagw13DDSu56u611WQ70PuEJuGkOnamWaLDYUs3LNoOnD/
IVPGBEtvRVwAUP7f44K+NXBVOmwdvXpzzUWeQmkawURh9Ml9cyKMHHdZ0JJtv0je
O0J0dpfCcC170I+DCtpIqmRTfZFPgiQWwr3ZmFW2aoKDmsuM9NZIHY5G5v9WxK/m
/yxLaCP4nr5sWAgiMph/TUpyOyV3ndWPmcKBeQHzpgIxrbVcVPZrSbhhSw+csmcI
OWFmW2MD9B0O8HgbGSlkFovRQcmxcTeSFtiJU7VyB8zwDiU4VoBSdOaqTAUr3J8C
VjlObMGIGr6Eg2iGWnuo19bIod/i5g8tfF06NxoQBtu4ibC0KBZsuFxjkRo2lVkN
+8pd/eE5z3amIdakHAPL79qmjEqPHKelDf2OJoN3+almi1mSacRHTKmJaCy4D+dN
aHq+WkOr/e7OQb9AaxmWHp071dxcr4XjH9R4+iDCpn5LVwEnQYw9QnEsQcgOUKBN
1H0P/hAVNY7Vs7F74/CsefSCnkYE93/1bGZEkin1p/EoxZPjwgz55b4QAanQu7je
0jgxdgrn7BlvCh4MhHpO5g1eMbAB6RnY2vUyb1oDy2cCH68DQbIFnBkftL4JGMgi
bNMohpNxsxSd81etc8SzpVcALQv5qa6Ybz70ou9mOMc31Tat2d8xaqljUnBGehC7
UinZTEINTf+2iQORbAfS5/aBUp60GaST6VJFDq70IPIpO2pH6kphwS2KlUjM8bZ0
96aiggCIdsXg+v1FRQLaMTOwuQIhi78siC6SGECPD2equxXBlbbFKtBEhgBtOne3
bzjogC5KOEHTLZRBI7tkgjeH4ZpGVwLSo8lAc85KS0lLEm8vvJIsX8skbGsW7oCW
yg2faSVhb7m+u/+32n6gslJDlGt+rjtMmX0tVJTGpUdnLMFiaop1e9DN44qLGmmL
8l2VdlyJkp4N/TLzFJRNJiKhMFeViTzkm2r8Oli/3TumCY3InAD8XsdYbphJC8q1
ol6Po8yMwXu5/rPofq+0O/MRhoQKlVRdrhtRiQaoiHThajzjFKfy5FU0xxiDc6sH
q1FDHCfXZuKDqdQweS7FTtdb3/nOPeH/I6AcmMeV5qw2a4dFRTL691FSmQTU1Nr/
ge/igdtrTW/oeyNCb0TLPU+9JNEeV/n71nTmgvhRn7rJRJWh8/l/2AQzf54Chihy
2T6gpnAaYVwKh4chsmhyQrTmW+dfjF3Pn1jU6CmQtxt08HSBlaFKFhiIkVjBxS9B
h+S++RLRGeecCdQOBLUsV5Zz2WcO96O1bLLhzLDvvB135b7uejXVLWNRrFFvdlWL
GytWR3x3qNnIZ61kOXkbJD3dGT3hUm6zC8Plz6UAYEpIBVzDYJYfUrQ7D2kt6rNt
p36V8U6Fw5OGXQQ82lJko5LWR7O8A4C0YJICs4jqOr+UsV8X3knfRf52x5+jTmF0
4qdhR7NGiQ7kJdNMAuDzprbsLfflcV9w3xiXVyPqPF2CxYuRMs8JTHYJ3tiBBsTK
f1vC/H//aJuIYq9L0iBShPufdK3RoGy8ZzpTYKGZZQtZ3d7uOTiY09mTfqOgtIEG
zEvvKm53u1kP5UAUMP3QH5lEEmjeZIKNxoUE6nZD4b5uPyO8DpPKhem4qoiU/tsf
fK6sdJLdUud2lHDqFpUb9ZXcKeQxcnwhFGBxrud8Q00w+0bveTM96naieb6GmWiF
bQvCMMrr7/aL005g8L8MtZIWkltxUtpJtvGHRe3zZvU+u6Oh7Jr/KJlh4PXRe7f4
CNmWQJu5a1iZj7tQjou7Y1qHfZ0syulsPrjGz9o65B7tUCG89ENdfMrTmNcUpNEl
ex3FC+hwgDyajPXk/F/CXQp+tHy6xd03TzqRS94Cza7W74TOf30pMy/Mrc/77ITj
0jY4i/4C2GYmjNmuYlgqtwf6eTGumSC2f+ceEEc+4HNdEYf+unfANMKjMA1AAnAu
XGIPkZWCNMEbmHLdOjGHBKNFahsiO8sQKA58J7riK8N2qeTwOa1RrlGwgfVDoE+S
BuKR6QPy1sjnJ7DNRrSPboJeejXeono269J5GfWMxQBqZnmtvPu5ZKck7TbgwQXs
oahlpyl0A3UxwZSb+sDaKvf2aOb0Iixx2ZlVOX75/VKdpPOrVtixFEOFfPmi53hV
9SbWJMb1ancqo9MAwC0Lr17X+N2j9kkWDQ3wdW5+qHODkgarjNbQ/6TSBXv4wts4
dywTA5C60HJEADoK7q7nTsq1y+Y6ugKY5Za8SLih/PFo4f/wlZbYPDVMswHLEOjq
G02T1QeV1fJfdJUvSy4cHUBzMu4q/via05KSAl1F4FLypTBVOYe2pjihRw3GNPwO
Fygc4SAWcLTGv3euTf8u5JJFVeKY8GLYa6+3mKiix8z5QVRgHL/NbEL5alxtET0E
MAr8KxvKxu6f6M8aVnZno2yrR0P5++IhDYXdzfJKDqF3KUg6hSpolPFA6Vt+D+Fs
58T9cE3A6H4C2jce0epqHD2PyU8kpmnu3tupkDVJBpFWvnpslXHL0EhtR32OSgmN
PYH6P9HEw8m/BCWmZfBFpAbfQkumMYk2xMYY2DA54u2AymVVftrMEkkvWw0wAqBP
dd9wvYL+jJjYC0COyFWoLo2chWgtlOkD4iThp6Shg2oYHgCdQasffsEQzCosnmUg
1TMD0zx9KuWgkiMzkspA4xRhbPZ3ZR2XN56kp11vGNUx0OVw5BmAitbBFnsh0fSi
l3ufpIakNwbUtIB578jCXiCNzF1fwOvGe/eGwTuMd+kpAapZs7mu+dF6alwTeRhm
FWyPSea2sVUUMsRCzfvP8oglkp456PuUQkh7NZ+D1PKAZqoQhos+DbHOl9g3Sbc1
69AfG38esNR2d6jY5ZjjGgBUSCAXrToScCyM/toWpc7Lh3TVZAudIvxffSN9TtjP
5B9jFXG3DVavCUfsVvMfueUGfGDJXIEVjfacjmBPeIQowKoVtH1W9wd923UhEjMc
/krSi5/qO9TQ3VY6ydlMywXCJKGHFUJZq0uc8P6oqclPQYp6dTdAgGNp+ZB5f22D
7fhXpq7Vr5mQyiqgeoNHKeiPeJkwE8JZgHhzuJCr91BosXWR7vM0LOmXKd7joubS
Gvng40+HJ4AsDWMCxS/Btwxu/51k/ciGvs9u854Wd89JvwMpzyXPoRbSNgkj0UZw
bviI3nUReyTWROlb+X1sR2rIwIY8VU6Kz5kpFrFY/0J1KbFWUd3SgY7MsD30ZYhb
VPzD9swA6H25RqKmRC0zaWAPRYHOP3VAb21ZlANRI0QO/CFwe65TMOhIZMy8HHSZ
r324h3uZu2KUWyROmkhvnqsjps7++11X5cTedq8S0moYKarI3BjcdNSE6YWOAAB8
SNUnSK59STcNd+GowupATpB1vL47lBR6yxF+XJYCd0HAu/npxTHtEWJdAOOC9OlH
0M14a7VoHvRE1E7QZeLARn1PXAKO07tZwYdB+oEskZ46tFMo/WMKCgkXgd/rZ+ij
21vBJ+Y2I/PUNdba5wu/uZXSgmg3+cKq024PqOEooRBSYLss43u/mkkmFwcEZ8RJ
UPb1Y2zFLRIBoj0J9APQQBXvBAk4IU4/iKzoWb8kvcNHdzC0vAsVYPrDPb1GDYY0
YZeEyu7AZ4PyJ3n3ZlHbpEccrH9OKXiLmoYOrYZKbKm0aIMX94kwoehgsFK5HMt9
f8+hcytzEsRkqZIZqbXAfMntK2NSAt+tCAzwXpCh2otAWApSKBvswP+lIDgwRcq8
4WD25sGJsa9bZKEOqalAZluoJf1RBFBaVsWFkHlXgF03l6pTVqKIGbSkZqvTX/7p
CbryJisF0A1w8NVYV67G0eo6twEb18HigtJ5ShrTMHD0ke/HqhbIg2MwKmfcJJmk
ej/3NkwplKU52bEbsDhnjfvS3ggkAyJmRnWq90BTTcikvPsXI9zThRmNcFGdy97e
qZSpFwM7AeTP4BSPrwd9xAxbsoOqUhjwB8JnTwa4173UUt3N0e7Qz7jIuqI8luNf
5sD6yHzziiJZTXWpznERAJquDhEWOHa0nvOMkNKNwu00n63+qHmjDxfF8uE2NF5o
0P/NUPk6iIwPxaxcuLD6FQuPLGXShwNiCj14RvxWwnGxOHRpERpTSlR7pgIOGSML
cE5mcIumYLpBXJwthCtsXmcSU9W+6Q7k7kDIZWgcXPSndKYhxhhftZBGVYofmwqA
ZVPHia51mpQ8fG1wn8cj08IgfMy4X6pSsvoPttZAlTRvu8kojY0vz3RU1ljqCie+
nlWHCT7BbrvEjcEbJC66kAO8Z+haXfOxCF6ap+U7m2GfFYlphCjh38BUgZyaX+ke
L2+ytCWQYRkqUF3nlUkwfRpH/3WrVFyLG+62uy3o85wXxVHfpvvTi1dODBJISoF1
Mb5Kll2FtjfZhMbC5h9MpJMWuj5r4MTg4JH9GMIOVpFAO1PG3ibvE+hIvId4rMQe
0cXfXw92gw9Z+AkzXr8h/8rSjmXDMlRK9h2BZ9C4eQ57kEglEaz4+PoK5JeEFVcn
TGHoXjLxIQKgzEjhTUfgG4sNkg7Lk/psCXqEEd/H+B23OnCTn/eQNCMcbXECICmT
KbKvd4/RXIYtG+4CdnopscQKLUdCcgddxjkSfyK+rPG1Mpi3MHQqvs3p2VBVjj9U
qPBDdDAnuu02yaHccyawGu2D/qQ8x16JckfgZ7j2rmqtqdf/dWgcbA0+lEWzMcge
Zjs2m9aHgs8xot9raiRRlQqcqUFZJb5rIH4N31QdetwJ1PtXqx/lmQqdTVfD4xo9
3UdY5AN+i6X5QANOcEgD2s9syIDwx6ELF9UDDr+QE5qsAwzFVA0a8gAAmhOvgsrD
Tsu6EXTwyj3debY6h2hHC21NSzTqjo4efwzjDWn+C4LV97wNiXumvolHnn01G5JM
lF2TXtZnDJZmbVWYVaJU4ETX7Nsq0BrjYXAq4Z5dFjRys0XysvENCmEZmBHiEEOo
br0ukjZCKI8gpJ7njbKd00rK1pc2JGQANL/0L3wTq2MhU3J5yc6N0B4ahOwQUZhe
37u7PV9YuHT8j9OQgXjvB18tU4Ojt9wUoG7JHomtfUV5P/MLjzxhKYL/6j8v2Ti5
1zu0tis+bCmQfUkFkb+zp+JI7eoniXS1hF7m/OE2mrZNyHZusa5gtMvpquUBsV30
PyDmYGBlhKd0GXpLgx4OnexfR0PexPbmROZjf8G608C0uPmOZ3jiJr8BGAXOuLOD
TYjRQe75tcJyoXTLmyEBSSs7BBrRmwLsoSopV5ANbufD1pM/GcfpkdY64f/hJg+/
w+hworHG5YPx8kX57cmfJp3Ri9SqkxJL2YPVNbUTOxCrszdIvB4ia1ZDDu02BFD1
8qy56wLIIKr6ah/DgfUH51gcTDpQ8zHTbUNzllMLQQ0B6BEllPAMsn21efO2mM9p
L3Bm6VofQt5/sUaQm2TG+KimMj4FgQ2Hkd0JBjoMMpZRsEAXR5/RP2yCzEpNyqtm
dBuF00Oqf0v6BhDpu/UzQ+Mc1trtA+9VZYP0hoYOB5E9vTYD4Z9e34kix+cGDXav
3FnNktflTqFxP4SKezvTOcpGDaXX0KuPAf1W4H1pzC6t5avpeI+gMx1YG1zwxavC
llML18tPTtNCNcZd53pNo5p/z22SWeI8Adgsxk75wdPFNRgqAma/yVCTXJEG3Q8e
sfPZCEx/jPm/YNDcJ3ap7BVSwCTxPv+Idv6UmadxG3L3+00LGTdOAIzKuUwnW+YJ
zWkLbb5hiYaR0df1cN93tKXrXHhmk8DqvpBxHHD6BA8yu8O8phBqO9yXH6DbITx0
SwfM33xSMpEjsMKx+ZONj03H2voxWuSxlZukE7eGpai9p+msyeE8cd+jwurPrGFu
BVnX2uoxESgoHIV7Q8T0eXfNhcwREVG2oe4Dutlj6eW4R7sdOTtwvXAkEPIiRDxv
CYsQ4VOtEtq87SP+QD1RN9Idrzq/zzvSQ4CK51I10yQD0QNmS62x2I1k7TbPSSHT
Qjd5FjrUuruN2JESAlIWFi3uqKBsSfCVdeelmi2Ayyx9crGdpvf844Pxs9FuWE8f
IFvS/xPk2BItBAq//vueS2d7avQGYzHk1BgRK7/QBfLCsHghNLNYiA1vbu7AANVi
mgUQJb8n/XMTq0YjWsD10qLh7glzSGGKxj85Iwi4FUAkY+HpGu1oG11Z9u/4wWig
kiPFmbbYEHoQbGQZ3z6JvanKz3VuJ/bfrFgRvPLohLkzOm6ysz7PLqTC9SXsgqVF
Jo6vu+VtMud3zc92uvR9oZTtK9CvLvC91oJdZoFl1uo9GEdL+3BOUCDixtS18mhn
e4Snw1hpZIVvPGuoX7FgfrUM8YP+/tL5b+9hVjKPTf/UI8hZC4s/L92NC26TAHLw
GqCjLpsY/d6r4bWEdxOYmK4lQUzrCghCenKTzw9uMsnr28jn/q0ZCODATrQkM0+s
VEwJ4J1OfsZp6RsVCqDT62eFkPpBavcWqi1KHWMEI28zuE+Rhp+VEiPqxWQ+BWvX
cr86OB5gNW5RHKy0PokNdnF1pHInDYj/hpiqh4kY9wwzwn3X1yLFA4EOLia734oS
DyLo/0IV6VfNk9sIdk/bwMjFXNnevMAvqp9Kp9aQUVfDQreI3bQ52J2nnlJhmKvj
47crD8LoY+YBl9IX6BTOCOQnzbxikDQPzuLUQ1A7gQgqMtIGM+UQ1XhPEytGO9SQ
izRqwbv1sNWMZQb5iqzARaHFpIW1BnZtRpwN3hSQFfHIslF0wY0BEI2AnWn8sT12
fHHLgnruV5r80oWix4VqaMOr8XH/SAK3X6D/qJKmmNTB5Vu8/RYH6uqbyvaRNsya
8AfaCt8ASWPH+zLWWCguVK0O1oIPsMed+aHk+as03qBvdksTUm6lZLnGk0vEjp4x
KqAEMJgYw9+gQKjotyac5oTEfgqPkfB0thAD7m+lgQ121BCaohKSP4tu+JaVg92r
hO478AraPUXW3t2lv96ZbZLAhuiQfXXH38TIChzYYDQQAssCwKxIzz8PyaaP5JJV
vCQjSkHpLdrvoBbCuHElDuBymnvEC0wEyQIkeXzkvASzVjNouBLnRqKnEX5pWJ34
EBu5n+jHoXCPXt6w70X1WcuzioRgtDaPgRba0DVviReiMbzVLmueBJhM6/p+r6Hn
2ldouy+soHuAYl79nF9Ql71IheyET6oqLphn2onBo1zQVIRI9cAvvQSjH/xQBawO
l8l5K/CD6DFbv9JGG0kGk7/YcrlPNr3okXDHuOyTZ5D2r/G08/cVsbSlcu7WfdxB
XwnHUkvgnReYglQqwEvlu3fEWjpTTbJHL5/ZKeD28P2BX/liudwdoSDBevViKCEH
qMH5mnG+4NCJ+WnHpADT9MNgx32JLp+P+Sgc8ApUh1OmZAP7DWkj2Dzwi+oBsCSh
+uTT/J9uPvYDVhB3/8JOWAGVN7tF/VNhPCz0of/aZAsgJEXxUqmoSdnOCOCvWhup
HpvAVlX9lNKr96zGBPFjMnBfNJDL/FVlkbwcvLLWcQ6MO4+niPt8E6u08X4JRzpf
3mGrDveDlH0W3OLwIk4mCXD0uO7viXh/npI6tnOtE9u8cTo3rCM0k2aFQtfjP0SS
m1k3LARqvzgKlmr8Wa/egVVCp2M9iXK4wKZbGIUD9eYz48cF6FSSrGb+3cR7SiKc
G0B/2Hqi4Fbjl5p8fmQ57Ku7pWHZ4LpnAbTZjFkYP2JfvFOtzkq7fu1GCSUBmjdg
ERrj9v7M6fuVCbxzKaHRw201QjWbmhX0FwpivW7w/tNW2c4fSR3Dl3d31Ke+yAVu
OMnHy2Wlv2rFwTtflc0fluN1mvG8BhVQcu0L9zvHV0iK/cPTGfKi3MB19yOYQwdS
93rkgIcXUlk8GFr13cz2bBfOkkYpKu1WhCkldiuK08bjMws/5vjHZQz0EtBM/8Rq
2sfHUMyEc/E8ztpBb6bky3aOMEEaJ6bTtYB31mAER9LDEAxUiGhMJf3qPUmctXmn
8SwkWdXcSQv3JEWb3rvqFX1JSe+wNH3vUby62RTDpJhs1/KU5z6/arGzHgVvE5kp
1Zx7LTDyTRGGHBYUtysf69lev7KjKRYivty6cUCkVJEkVobuuu//4cLCSdJ/u94B
cgfqY+pq+fWsA3wq57cieIkUCVulcQ1cpSnPjTk67fw5yl5lV4oslZdFVlWkuy7L
9IYwB5IclIGHB3QaJfMq8fkgzWpny3fsh3zUJCGBL4hfAV+CSnbj1tVDen8+cDGN
mGzLSczQuU1Qe4shrAJ1NWseWAgwDh19PKgL6IhDi5OMf4W5AdvXPzzXxYcQJ8SO
KYB/uLH9dHjIOPdMJa+kJAAvLWHNpI27JGHuWhVNS7j/Dx7z8bsD6z7JnhZAVb4C
Gtl02iH+m1i2ggRo4jkFGd3MwIEABf9wgrnym9td5Z3DpFOvKeyChE6k+FMNxJG8
GIbjHxZB6q1A56KdbCpfyCa3CMM5w/tnkR5dpfOceQhrhbzkTaj7PmpTpGBtIkNv
gVUyVZAzLo8IuuvOiENzok1cyxP7VJgzj3c736QwbiU3aFjSD6vgaNurYfRrRDJv
ilFh4IixXXK27eriuP6libqRqOZvLuFTM9L/zllcaKTEOVw0w8LTpy2DxXeUDu2n
SjlhmVT0NtFr1M3z4PTP2E4P6QncwBzM7m5oqiKTYd9vGJ6hzmYp/0UdJ/EIbZlO
216r2Kl7BK0EXpHJrNLXXmKHUytgLNsPQIF3g/Nx/Q68XCa5yS1tyZgVfKUxv8gA
vju+Tk8+0YoY96cqHRKI/oeiHY4NcAr5MY8gGQWZdO2K2lQ4GouH0p3Vlgdz88O6
5rGs9CXCKMwxJ6G/+ZdtAHi8ba17jatiCd20ouujXo+YxR0YryjiH+BKnvQfNjIV
L/2N9OuxugxPeV6SQof/5sxzwT3PWYD325m+c5xFhdoIYcXTjhjaixaFwiEnilta
qfrcl40eV1uV/SgGMEP2vheaU2y3CLntEO/ihYkJzhFSKGTnUNa8AzLSt6pEfKSC
IgrEtqFnmbrZXE1embJRE6dcGW+5Gb7mDOkIOUXcprHqKegKRBN2NZAz0mtmVDV6
zxbxilRqmk8fP9Ee0zZIqMomnXfNozpT0SuvK+CuQXZn+q+rsVIgg32dQr3xsL3e
pn5VOklAfuPAYS1ul1QMOkLVgMBEL+JhbQN3rcB1QTo4vyvfnM8hzhLB9jx9ka1h
FBHmkU0Fa+gUL0L/ZSDoblWYa3f/tPJbLxxfRtFO/AvLs/24vzYl3uA9ojcGGd2q
vjoqCfWccsi904/H9Kalp72JFGznX2N/WSIPIP828SJG6L3bJUq8YKoHqfyKAHFO
MhrEcQY2QgMK+9arLBIGR9jpg1AgJQmENdwBeUwn2ny0pdAy2JiOHjujmkMANi0y
bvwL+2JrqAKucDpOOmpLfgPPrmg1fB26iMsW1wP/Kfc+QAkV/1fXk/qkusWjRgbT
RXYOxkKZCb9vBY88bHdLBfbAVspvUKfxprRUzRzddeH5k9FgJFw8ZEeySa0FZjje
MAp3Bnelmrjej6zR/00nTGNyDa1Jr4Mu8n1Y01FBtahk/uBIt3dRZX0K6Bbz3G+n
qBT20r/gVccHZkeIorAYJX09mdPwwhxoVPKkvpuhBVF+jRHZhTBdtj99huKRwrli
oeSclFcjogsBtHoa9iwr3ZPxF5yVi33JNAZvuYvtM6BcuWCXexXDmQOnU+z3aCT7
xmlf5PXhalIe1b82PtVgBr7Lq8mqeXvupOPMpv1lvaLgl1VRMKQJrKpZURJCpsXd
UsY5sRTt+/W+E6QLpugY/5zA8+gEZfBLd3L65FAtD2fcKAgUPqHpW4eUJkwWsB6p
rRDHRD1MbRqrpZVn+jF0vUWdT3YGks5P17OlLIr/AClv3Wf1rM2+5TUI6lIP6gAK
PCtdJt4sgEbfGnLkta7Su7Qd98VWGlatTVlKGsDpw/Mo8JVmSR6mioQNRGxCGGED
7Eg5Cj6KeNyH4MbaWMY9qd5MNnEy1ZyoLfe0BpeV4Mh86Hqo0I/nbh6F15ryEfz2
l71dfFbT3zc6Ki4a+qBB+Ut7cj97Z4Q9DMhPUTsq6l2uuAWWS6bbQPB57utXfbuV
u3OP856BCxF/w7I8cSPTBnY5mNRciu+y+T4Y9UOgjLkMPfLzT2EzGczoPE0afvak
ufw5x2QY23Eoo53NEe/JX5T34Ir2cE+JFM0ToKh7A8Mh1o5w7HuDSL06wmpADV/m
3pMsjsWvIFRP0vYpCTMYLCQtzeE5iLL4jaJNnQwKY9E6a+b838E28tf8N20Ml1iK
QaaFSF3U1xQPbORool0Jb1X2DwPZ5qMtAccsiav9l636shyl9g1PoFqVCzCqA7lb
zRq5pqQjr3WyDnpCeUNJIBgg9g2G60uKzbAfL/0a8/5XBZlJW0tW67/IlIoxD2yd
oT1yDT/szLZrueJJGUnAFbb54aqB4/PFxWQHil+fubF26eE/2BwbuLVFlrgI4Bjn
Onle/uKVGs3BL5xwpxq6IpwwnYtUoVqRK7MNij8uMObg5MF8X07f2mOr/ipacNCH
HItaiXzoLAZ+5zKlRJ/vazKAVv3Jqz2UoWg+Kz/He4Jp8yvQ1NULp3PKGwu/HNid
OkSSruJAgDWwmnE2QOzOtmn8bRZzCL9wkCLQ3YfmDXDqc1C4to9AJOHRypOkhjXR
03ebuwCpdT9EQ9iWuo2vjnXJsC5p70/jM+oqViSkfvK+UuLjJe29KnM5HliYeeL0
dNfmz1CtvwxaAsgPfhpNJa6b4i/SZgT/QUHHSB9PmbCO0KmEFLibdz1FxdcUP4MU
LxOo2Hb+fmSut9EAD0QjRsK4zsx34Ee+0U7e+FYdhWk4B49fhtPw8I/bj5ffMAh3
1bIxWTRZw91rVuKcljskbmQSfdbwSxdJNyk9qFcWD57zt4WqHsxfU2bMvkynFE4P
3KJwe89BNDOZuB9UyafyvOKP7li3rRYK694KotNYzrhMRdPYSuRccnLYZrBNPM4+
IwcUjlxuJ9O1V3M2Bc0u9jgdUlzs+604Tnp95opLwwso5jsWhWL+CWCdFFl1VikK
m08N6JN5CtsNp+ov/PCvnv65D23g0hy07K/21MHvNE8uNjJ8Gz4oulRuHA4ZZ5K7
n9eurraZJpcQlj8Ch+RV8cZ0SEx6t/PtcUbdLWnMlw9wgcyySwG7VuaT76ElIzQz
6SAM0H0gXElSmjpFY9NV3sdh/koVIjT7+Tk6G/7MLRVhbCrmnjhSTav0jN3hB9DY
9Ie4t0WRHvU7Vkuv3BUprusk6gmXdQ4QD/cWSZsKqcXgqWq5JtEEnwv5wr1qUc0x
vdhwK4iRC8m5JIu3D+R1gNQsmte2IZGuyDxYeDWp44MNyOXh9psdv/PAiXTvmdxD
nwSyvGYwSIDJSTmej6mF9ZkN3JewakHfwcTDODguojw7JuMJSc14tKjrj/CgYMms
8ySU3CX3hS4GIxRu+f9kcxvPx8JvPLAOkYzdM7vzGUa3sMFn28QJKHtYAd2A4gp0
JYAFXscZNOS1zaeinaV9EPJCKirnm43q18ijbTw6TAPqaLYvd6RPKV6TptD1ZtN9
PQwol+lgFEtdxC9ColrjQr7eOV2ITpnXAILd8cqhjXqdYusX+qAi0a0IcyBYAWHB
/HJwl9ks/RXK0tmlVBDdcdF4kbBAmA6bJCFOFa51/1M5IKwEkxZhl8ce/F0LoAyu
xCByhmbiQPtlZLrPCnNHbwaBtUbodE2rxHHao20AGasqYYd5Bv1jX8SOkIlzUDTN
JocWKIUzbcmVvGBuoXhu2W1nb/ihxoJ3D4+3ib7zMjOKEanXMQRr32x4zOQAxEvL
j3L0JjHhKO2NiDAIg+JSjx+ECNDksE+OACI4WVyIPtwZeUKxzGLXOBe0t0yqjKL8
kCJDy7TU5Y8dtc1BCnJOSEtj53KishsYw3hjPf8ZYQIBIYpmIbgrjc6Cdjfwwngj
FskjdFKSiMBTr2CTp+wUkLNoVWMLfDny66IaaOxWdEaOx7N1hAU5N8niLB0ojfru
Jkb3G03JSrh2wmjc4bumXGtX1SkAeg95vWwugrKcC4r1jdPqTiCJGqxSZhLzA0wY
okR+XSDnUtENMAo9KVGgC7SrG7mNBxu0xIqoWFSCLt1/nFyue/l6wgWbn5O8Lj14
Rvhjn40FXBAXmjBP/Mu8lUvwmuuVTdc2xOBamL7yENRXrn7sL9SrZG2fr9L1J8I2
46zAwMC3rrPKHvDhHRT6EPmOW/OgerWp0CTKT60qaLF+B5QnRjKmg5E73f/b1+XW
P+e7TUrhHxJIYT+etkZUJLZBBHJIev8un2rivOk4sxWE9Am9FwbTfEgRtILktZmH
tndK9kcthShhCbC2kNgH86otljGVnQ/bwp0DtMNxnqdYn1O8EEs3YXONzKXPm4Xg
Kfvk+gcVkxqjnrKsd41EKsDM4bo7NDKUwWquvn+mQljLxXHIfNur9HiBmLba7JxG
VzE5HbYCpoN3LGSdZFmPAc4WPxCDosXgQ6ujFdYsRKsy8rW9E8wx5Xa4b/BQ4dBG
WmWpBndwm+67WdJWD8ZQCt11RotkaMxHDXOUYiGzfsaboGW3mTRPfmyMrcqaRL/C
RnJEQeTJmllVuelhOZkZOVWdQc1O0ifKtrWFgziL8WH8CNzJSnRpwjegBwSHCFk2
7BeRCyABWEnWjmx924Py2NNXAw5uV1fnJ7o8EvEOuNoaNgyBU8Nf0ljrT4R+gXk9
Wyx93cg7sabTrXQEk1RTIlBNsQHzlX4m+sV0BypuJyPlpjJZUHTKCp4kHADVy+8A
HnJvEYMSITp4qK5Ke/3ibXClTjEMtRG8UxDh5X97ZkDfBAaoGQLQoFFmUTut4yaQ
ddWMZMdz1NALIbBVAYFKeG/KVg/K6MVMTkqFoS9np658N46YMbQEHSfsMG/h40uV
N8/0bx+p4LFXobR4Ka31dgwMnwkoR5ciSTpv+vuol6u204q4qAplzc/J5yhhtk9n
eeNHQ9YvI5T2bWFpb9JFxleGGxbsj0rDi+vt+38riDzcI5C8pim3g0DeZZ+CFWzS
HrqjKQy4Y4LIOcH2KH/MEvOPohaNf0JDMl5DAPXSke5YyQX0fuM5p4vE+nGe+d8p
rKQnsi79LS3nI4yMuxDJphGDeatrCvRiGpPWO0W2FzWVoilPieeC4bfwzjmkFxVA
ISYr9Ade/TpMm7u2trk48N4jg1lA9RPVcJ345HVEfGTlkhljKGP+b7rD4YL5DWf0
1FLm+qmmGqu9c4bxDKZL7te1IjugfGRzMghMO/b4HBpS3kmi3ut+WhhEfpXfZ9Hc
T7jkSwXgIzCnXw8/19cG0D8Qj/eiXR2ABvfs51OYfbjGF3Ehjt4notWqATsqAv6z
KcOvQGuZjJGoWBsV4C4xfVG+gf239Qr1LWiH6pOGP7rC15sjJqMKtsSVJcelM9Kc
4PM71lFY4iGUbWfMKZxuTUGQZZQK6nrj0D50SmDSMWJySsipB7aw5VhbI1lxllyq
awTJ1RWaBm4EJC67VyFiBexKR9s37cEsncDoWPGH2Zkwwy0l8C3AWFg8gnE0ugR5
53H/PDufCAWtbEs1Qz1BMirA/4BX4EGNFfQph80NSUylPsu+tSNNCvhAWU9V+iWX
gLG9m+55z+UPs1bW9x/34lp9YPSwqCyJYaW7ZHGpWThgbqm/2osrVdrLhzlN6zJm
DEgqFw/3KyB/Xwt7to3tPsdhi/WjdDuT+RxtiCCxUdNa3h6PpqfSuEGOmtQx+MM4
ntwBEweksSkqnajXV3diiuakwMYzq9PStujekxHVxEESzme5DL3B80HH/mlKDdcv
SWFOg0q19Z87ufps5MUFXWM47bbLx2unDeMLWM20FCld1Ca1QNkZFJ0mjrJPRUUk
8aiG+2c7D71gnqP45WJssqAiR9HJwTeTK36E/ua3Vorr632ny6O07YS24LJmqYAT
RgdKgKvFJhifsoDKcu1ixERn7E6I3QkVnx/p62RD22xwLV/URycafxRxH24R9z+S
o80YU51E+BO7Q1iCXd05M1ZnZ+/ogkZDW8TnhighpYXMl05hEn/OAWzYe9RBu6lU
IXG3+7Rfn8RsutZ6wEuuPainxmcYrHMJyauApeTX0BnD2y2OLs+gLywRQhnruZxK
uJusqstiRVzBXXH5RFGMaexZidf55FeLTYRO9nRn3gWdM0QIrMnAEIWIYk1gLibV
6wMz0tmJ2Dng4F4qviGfwypXNGWP40Dli0gUMJR7eyCGZeB7gX2dVBJHZw5vJpTD
vJQgzNC5UJF2yTRdmNx/wssTGoaeHH5YSePKhuMz7BaX457Cbti68QHZFVIJyrre
BBSvLPZHngp8ry0uT6Bgs1HDkEzAVrsB7n5PLulhYkAHi0S8mX/GvlkKVv0CFB++
Z5BZyhry+lnzI6FlEmP/q9zN1BQXas+kupJu/DpMtgcLCYf6C9lPLOGNuAU8nFTS
Vftvt1E0KIILhuBQWs8tmrciZDGVzbTPgP3RPxegcKnGyH7VwXzS12tvEv5UEOQO
4F/+NbZOTeVqnV9aT+Hi9Gc0wWG/d2PbfQJcqheNVokCR5BGLLTGsdK80AqMDacb
YLeiuV5Qnuj26BsIEVl0VRF3JemYikolD2bKurHLJxt0FUPs9AuLcWv1emurVsC1
w52///wphpvDSd7ipxZoshEiCl76o9bLpT/ZXkvKmbl/flECKaDv/7Izu0xSh7xc
hGuthAt8R42kzKBIqCXSHGc1GYQ0xUpR53CevIh/sn5MaRumYbxWIi7k1qpuczXu
b38cmpwW6HWcXXhcqBzv3jhcdJMlOWxajX4Nwhwfp6OzhmqagjFdFCJ3yK5eBhIJ
aFSB1a9yR7qQCwXihv+9lDLalflAgzkqnlYNTg/My0UCnlGf/1WSnJ86gM+Vi9gk
RsK5H7LJZ7cOnFXx2N1+W6gAkfL6p6LRxx1kaB1mmmeuYCXQCKj4BBja/66dYW7E
wqxEjl/VKCawaAq6QH8QcRGrID3fbTkkZoriw2O63zOxofgmmlr3mq4p4COHAPJ+
s1ebIlKyWAVEYziivRbqZ4Qev9ENsXEAtYc0dBgO+OA=
`protect end_protected