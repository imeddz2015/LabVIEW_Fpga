`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 21808 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/9huKRhRMtvnNqb3Z+UU7TahEoHV+T8U3P3ufru7l1O
3DlgtZzb9QxCbOjthp9+wDkjygH0eUfDrEl1ovhZG60TRhA3RbXZqp/OOCx+1Voc
am0wwZnA3tNCq3yDKnKcd563+CoZlX3+5EPY2/YhjgqrSXmmH/oJiK1pLrx8LTcH
+HQnjV4y2dcSuGYP3Xct7FEdwIQp/AC95UaRfG09JnBlg1ZSiwq5qjzBn8PQHlmF
nOVexy/NQlyBL5t1fcTgqSIfgYdkL7jPy4T5mAYG2HFCkLbJ4cooP5qQi2KTgk6F
Bht6RhD7N4WKgWlq42HB2Q1oBEo4qBcpplBmaVVx3JkKoXOle/xQdLfdzURmEasu
y5R4aAUOOmwYitqzyYGbjjLFFjezyDu7wnP5fkr2/UAdAVzhmNwGG0+XLvwwdDnL
m05aMPZfJJYlTnYNrdNQPNt5nxLEZW3qIISITtNAZEU7Cvhh4GEQNWsNdoDA51y7
a8jutMMIQZAyqOdNCd5TfcVrPQF1EgGTehiZgOBBeLwvCrGz9LH9JgIuCQwepnS6
va9TLDqcqwn9wB3lZrVwDz46RN+rudLvqCkcIqCdu33pqTnfeEAfgk74rVObINtr
W1m9lnzwxrKsX27yHtQvkMgZbGZAIWJDAMHseCZW72yU4u6AbOy77UHDbUE3OJl2
/3mRgJyvSwXLgg2jPdxz1VgFSZUwV6RtVF/xm7vTIYlFtzViaIxUQn+ElvL2erqL
0eIusS6XeDv+mCjKxiRiwCl/d2Pzahsq/q/rV4SIds/tm3jzB0k6xjm11aXLPHrC
cThb4MHsRngPu9ftOmgbZisvwZ208/6GoiHZZC8hqqL3F+SiIjETZmnuXh26JMDw
27hSd/f/IQce4LFCRAF3526pwHLgaTb/hwwbWXVwx2RK1W1ggfBrLAS2TXSZoDhp
8o6BJxBq4FSEUbM8HZByA90rAiRxufj0OmGte3iyrB5TRezpIAuw/V9zYVGNPtWW
U+nGpYfjxr2Di9ODWgDgXl0iAjZHVyHOWTS26fTmnGOZ5OTfgEAHGco8NBvf4l6I
V6tnF1kr3TAMm4ZR4GHGDtAyfnuKjJRDVjPHQwpeMEnXPPPkU4AvyUQVizIFvO4y
bddSEQyT+uovlPL+25yHSqicWGHQ24Uk7unp8NQOAaGCiN34kjs/xCTfjORFvn7m
Q6vLlkX0zUUSTCS16dLTUuW4OTcv+z3KhPIqwfD4MOeCUBXMUQOsggf7WQa1yPFT
5/DpW/+AhT3b/XzJyAFBmXpXNwXCUTqAkTwT0evQBR20RMtmeDVLcYlTzgaXHAVq
m0yPO0SDj0s7/aEc5uDuCqODS/eBmzfAaNdPbQCuWfLBJsnAjuIPjlibxYCF49IO
c3cT1Sp16nyC9fvbNF0WgPJvoQXwm5ZLPLVNLwKzLE2R7FDGHfGS2xdzRznrgMre
e9gWd9eAX/nk7ZccaJC/IOoMmzU4ZjkUWoX9GKWnidxVd9dBGfXAJy9y2asHZKqp
RbRUfPCienz8aWWqG0/J8z6tqCX5j7FTo1XM0z4AQ/BVxF9jzrvanv6anw0/8dG6
mdzKmSBnX4Z8w2qMxNBzvM1I+siqVkyqkGdtYS2Q0AFcgB5yRnYJGIHoXAJOn2DC
51HfGtm7T4yLMOy1lOJ8a5bGGTCNIHvFZyun1inYsNozj1b3fWqcYedJeDa39sVa
xDMZDG9oB03zu1jkN6/ph2xGSsdcyP/A6VgpbQQCY/Jn5+jd99T+0KRKhWWD6Kh8
hHckZKK+Jw8XYU9iHko2wC1Q4wPPDcG/wju2oiyZ9TExF0x0SaHdQKby07fxpv2Q
LaRRalX0KviQOW2DzTLIg11XYqEzA4KKcmrm4FbpqttYJdvunxH3+/yfLJjyus2z
S1hNxqY92+2WWolIuQjJbMUWTRN+vQflR2I5wpDjkP9neXbs+Gs3Tg2Ah/wGySvA
0cbyr9AgVbtj1n6pCkAUp5Sh3PxMS1MKqXNvOW4QKMBwRDhAL4J9U1DppiJ55qlm
Z95d2xqs636ZMADN4iBd38yI03TJoEsbYSbfIDRlDTx+XsGXDJqm1P7F/W2Hjm/R
zYMoJsUnhrcK3OUbl3Bi9UrufhnbWCfEsEnGVYUGNgDcbYLVbpZXLJMEvB1TndNy
tBJmGH2SXE053kjYj0l9/nNBYJL5cx1oPfTgxl06Urj+6dvRkuoe7xA8CiLVKxZ3
Cyw6Qt6FbSxFhHU183eB+MVgyMF/gmL4kDUgDFkzP3SbpSYJEj77dpW/HgGXz+WP
ww2ehLnVsFZFwnW/Toukwtnvc900J+NR+XFTXDVvUBVqGozGGhY/cDpPbaO4Fnk1
Um2PL72WoqCzGKx2hyGYtTMYCfRFlQIU15n2JS6nwuTKHlvrOy0w76Tb48pUGXfS
OkrEy9k8rby/K2flSPhrS2DB9SJnakkINrYttnV1JUNogj8TuXsGEvwDKoVjY/dX
uiueEe8tupLd2clNgDsgXaCa5qKDIzJjQ8VVKkZehOxE5ueu2mzDKKFvFCxAo9ci
czadnL1K3FquBRBWPCGQCk04DaFD1uQJKlvW/2yjGmggj0cAYACo8INhJYXoNEbd
yJ0bzvJS5slUD+jRE/FSc6TtMwvXG0ZpBdEzfQeyn2Q1iyB0s+2qDc7tyo7x0ijh
N9WiuUpSSCzIADK9VqOqMtK35YsAOX3q22FfNiBFSO187wrfITSH2yuJ3qryDmlE
5a5sOMYZBH/ezFjhBlAp3Qul15kQuG2K+UXL2JTzbDgVoILU4NPt7oG1yy9+uftd
FXEF3DE+RTbZwr9BmgdAiVMmSRhxSWvKl8ScgtPr70aL8RNoHLzW9VexsBtt02JY
gEexfr1+69f4Bm79j7KMEfaAgQ2ZSymM4S/WXvD4/DIVYrNsbZhZOu3J+U7FIwFj
frQgYXmK3aMOH4ZggH9daU1o+IhxMQ9ss+u7a1K7BSJDdmJjPA3icv+zTr5FKmwk
7Jf/zuA9Fw/QhsEXO3M949+mIGI4ZWIIECvTJN2lv8OzYU8NjvZ7ziu1O4z6kPYp
XTbi5BmOftq6LMq1tPGmsWQeMdcxUTY0yGwRIYeHYIrhtZ3JdoSakVck8z0umBnP
dKhoGBGq5qsvg3zuJwgAF75VsgLzHQXN9Yln9t3XOnB5DbDgKHdMPHBEnBpRWIKB
5j+nA5AWvoiV5Hf0AuomZtfcpdgX5FkcTaSAyM1aZIM6l1cW4MI0Z+0H3c7es/xo
rSc0lyNGzzFYoo4YOH5UPjmtiLdbyln8lCDOet5ZulR/kPXrBsMoJnC//go6zJQD
CkQWfQco7VSgrjD+LiyQ12XQW0q5pG/Hpu1+Mrb2vVeCEUdaSQTSTwZn2AC9XnUD
K1+wcSLwrdoPv+cyYE618351jhXVyIQlBf0BHN0Jdp6IIqkAk8HJKe8iC64tybd9
RtMbQsluitCx2V9oCDZYplLTeYz/iJeDNVUFE/btsVfajv+F7y3eHG5z/++QyhHO
4OnUFGVqiBPkmGWrBQ2QV+jbAJyA3AZ1fuULGQPx8BP/EFkeKL6UJerJ1p/Y1iSX
NLJ+zOEMwAUc9OjM7b9aDvIYa6UXxpSrxIt+GXa1djoSN7budhGDSNs3eHvtv20w
8pgJOuVxiIVwpKmX15Lq/+kP8/0prwMXbhtVaAotKyFq9MTMvVeOhRFDJGbPWN6E
bic17exj/ZBp5VsOv+ccOijSX/TCI9u0oauNd7EWB1e3DsikE/qGNPhpb6JLI6hC
56COuQjLoGb7YrxwYLBjTZWpuNTpgn/Rke4Kn4Q40Ho4Wyc/I1zDe4ay4oqkKaoi
pBjTUCvez0JD+5n2mI+8nQ2JG8TN8pSP7JE+UYEL2sCoqfelykvECEugLRvkmkPD
zYr7sMKGxv37hzGJD9OhLk2B/c1v7lk9CzuO+86fhld+0Z8GTNi84QsRcidcoJ6P
mt4eW2H3rB0gHK8jbsWkz6qjPzg8rwCObKgreUpBGkia+HXe4/mzIKxSrDBLwJRq
lQ7OvSWhmgTtxBvdKOpaI3xrML/Dcp6KI/7mJ6qScqpqGGC8U5+QxmBuwdWo5KZ6
TbAfWZ81KkFphUpnHywlg8SKeFeJfQc31kdSicy2ngSo10QxD3UCpYoZIQ/uDnAi
6yMNVrGmFOzurZLNN9LTsw2oOL0L8Iw2+ryXE0ylfQEjNs3zKdFNZumhfO3dFaCJ
KZ/mBRZ96mwF05OstJOtJKIfa0UT7KcUz8Zi6pkTy+HI+2LcIOddMF2mW20Sf8Wm
UGNlIeDwCRScnzkcmcWcJqQplsXoG+TXvtyXYldhjjupaZ5XeCc5ADxY9VljGd3K
tdK2jk9Uax/rkxH8Fcurlt4ARKSPnyBYCrKEWhNgOHtclM9d0qfENJeXDBP8YMR/
RDbu7ID/Rw8SXoNF8RjkMHfBB3NH/yEhR2LjfbtRO5tJ5my6ZrHPFLnBLstMqOgK
0xLM+ZDPJ+fJ8WomSY3Q+DVu+PWGJzvJ75BQil4hsbE5MTdz510J6zh2hsa1Z2HL
HUTVXh/JnjygNFfAqvWlpwKswxJiQvxv5Zxtu1XDq4VyScRlua9wscyIw7cIE1Rw
wgZEcwXMv0zJUlGv3hazbL8YAHO3yyQrdLeVRhl+hL/PNmOgWn89B/FHhFfTYp4Y
UujHC2oM/Ey7e9QT3CeRIp+jmc4WxsjM/ViQD2TUxpJcdXCF3Pku8pWOA6grXSmX
P7qPZfvBaU1/VrUviGlZyE0aE7PKqWlRzqBpFTioadi6QCwSGghiKzrq6oJyvgRs
1psFkthQP98FCLAV73EirvrokMUJcH1/FWihu6j9Ba6FlE8e03RqmOvN5Y6kN3mn
0LLmqgF2dMArEXj77d08FAGev9KP0wpoP4tsLj7huh668zV0EdLXm3HWrm1X6UtT
TubfIuS5v1MN9sMohDQNbCSMQ3xDc0g00zcCm+rAkiVAkrI31JJqk3ETgXC3xuAG
6evtH/+TBR7cptILJ5zZzJf/gwb5zT20t4kAxqicLULRxA7rIMBNk78U68rcQqjg
+6vOUuimrpcY0nElQaCv7WUEmVdNUwSEKqFNau/fqGDxOv0YEcfREC5NHKSrtaLB
lK+LUTZvNJeG3s2A8zRnX2FPBQMeCZ+jf9OCbRteV+TozaXGSS1aNrM2gDj63o2u
eqaBCqTNDLPj+u3AeWnF1cgteiZy7rGVXAjj5Lwt38fECycCHF2MkKn0zNLKMK3+
qrrmCpQMrz33isJqkOFlo7hA1lo4J9lvdU/xGUobnJNl222xr8a6pA5KCDEs5M4z
SDkHXd9f/lKeMMiSrCUbWfb8Q87hMyWaovk23bPm07ZYpyzOQT+RbZmQTkG7mcCO
I4N4VEknhu3Vhl81VsnLs/rHa9noIICx8eCPxFraqkVQbPtILs+YX7OHOz/APFhT
wk4Pxa5yVMEtAByTAWTgMYU22JW2u39NZEGacs51bYme9KeUFVpZ3xUzpmHHTR4C
uGfmPSALsYofzShseI+o3Pf4JM7ahSU+Ol+IQkKaZ8lPk3+wgy7a8Qd4igSYjy7c
k9ypsK7zD9XvncMZvuiW1gdn8HTMh2kSgRkZVlg9kfvPOWCmha1/bORbnPgxYvPL
iqSWKAwMd8DmRLHL2XJPU5X+g1ey9xiSRIUerqER6d/JIrBCX7YtTLG+RMvImd41
iPcE35Ovf6IweY2LNveR2j883aGtR1+oKhx+y6rdvQxwdxAWDdQVV2ZJSm5UpYdm
WLNEwF9Qazl6cQhYzhKRLK6u2E+YQU7QlEYEpWoDVyoCAGYvPkJC26PJfslkkmMl
wZqbbenHHZ9HGHuOY5+Qa49bLlI9U68/1cYgTRIlioazLZGqEDJNsoVdHLr0za8N
dyzXVcgfuv+TdpROYCiZ1pXkalPbe93Qn8HmOEtBO9gN8KTR7CQgij3syef6YD61
2/wqKwCjzozsVYqA6w43XxMxiHLo1rCiLl2y94h/kBfvFM5yo/D3tSmar9GotbrM
n/qjOYOgj7KknZv/HwbXtP8W+Fgaef6lrxcziWHX8QqX0nNLX7EUUcpRCySnGu03
8nKv9KKF112PuHgM8he9UK/cHxwqVbtLHZCyqsr+EmBILTgU+nau1J16Xaq4Zxg4
fHET6jjGj/OAw2L3rL242NHm05Zru7Li6IYIoUvgjOSJbG7GonQyzlVe3sTQDxHS
oFH0YhrJam6Hyra6T3FE4K44Nw8ApH0EFbecDPA94WIpMPFjJl9WxA6BrFCTkCLr
LDQo58Q1zrnekGLiLuoazePCzXVl/t4+FEHaeP62l/tvVBdqDANcKmB1gF0qIMth
4/VTzoSI2yh4E13psZ1OT4eo6gw8SboNsEGgeY9SjRho2wLJL0NMUFnJRiY3Mt8C
U0GEgCs8W/PfQmBWZwG5BonrLRbAhzvyYgCeYaWX0BETaKw7ZEEhmpf29+1mTBUV
DljpT8/v2lbf/B6LKHvubWdxYVVWWq5K2ZtagU50iQAJq8xHPtOlNIomBPfslW3F
8IWy9nuI20toe9xiaasgTIM3L2CKqBjIHbYY0JhhHgYnA2rN3CtqtQ2EuM4+FLC8
3Ps+tFSHNiA1m6DeyBgN8S32/JbwnyqO5RkLZ1Im33wtmU+BKXQ3vE4wfs9fDl0/
i97F/yGgRA/u4S9VCBxWOWXx5U5Z+0kM51i0rGolnzQ7b/15DWB5i0CESblIyN0S
lLwN86mIqgTgRCvorb30+KwBvarK1lrZFtQ0q3152H9kd9l0Joz6uOfA18nokW+2
PQo2++0BHQVoDbS7kT/J78ywkVNcthduethfTNbYva6ZQ8cld4k1HtxNuF1rK+Xy
T5zKm314HWfUXJWvBQ4pjei5qOWrWRYKXU1G1z5nI/P8RhhGXoSphrNZjYno5WM8
8dwXBT/NQTMzIK2i2RFYfuY3yQD/aKw8J69R5jYqRZDYpbuoJbs9AMnvmkjpwgIs
71SwJR5FDjqTL4irhPufSnYzoEg5WdaJUoRZLY8wUe7GaVmuRyLx4c/O+u/Mp1iU
nf6247f2/kFlvVXkslME54Z+ChJ9eR46lcMttY8A7FJXbX1Sm4QYvDpWRJMHtqls
sqztwpoKmbUK6C+K5iS47H80PMm4NcRREBBK1ZnZpOmVM85cOaS0oMFzdtc/TgYl
wxCM4kFIHDjhZZ3L9ybnAoZ97u+V/ZiIaGhO+AuLEGaJUiFe6iKnvXJhCnSuudve
saTtNiOdKu0O3bPoALKnsVcE5a1RcwB3HI8q+6wW547liZsX6XQpcaS+jSrMr7Qt
2itiO8EatHkgMCpdj+qqMor4Yxe/TMyiV89Qdji/Akkh0DfhHpmt6tEZRsG80dnB
tm9gfPsVPX3dQit69cJGVawsFuUQaHjEyWKHiPAJzoRAp0q+IXa6VIXDqnHkA0fx
bqq4OY5uQM9DiS1K5U/8Gf/0uMNRnuKFiTFSus6yRa9/ppL7XTzU9ZsBuUHKQLqy
EG+oJ1zxSvUkHSlNO9XIV7kmv1Ofj6G8eYVBhvF49Fo0/Ba7HSUctMKceSy78MRk
z4Skp68R1KG/09xF4CEToqyyCItILuF00DQnvJIRetRHKW6sUGx1TNrhY2g5nyXk
wieMFLqsk6d84iUEWl7bqjkJH0KQnlmTp2tyPw159mIU1VGgJU2j7SLC2WJZVnGJ
IJghPAzk+qOLMsItHilswRnwq5ufUYc0CkNo9Flth4c+ARK/qTcymjjKjc0JfRxc
D1K1FQ9TMZoS0RsNYHVAjORUvcnPyEP0cBlrDZ7mk4ooDAwuN78RjTawynsn58LW
AcO1dwGBzVKMEswyo7r7rK5I384pVITJitEu+1jtBx5TtJNPv7dl4C5MbUbG70/W
cxmpWoRqH8zsdOymTYIjuyxR/tppHsHQIlvPNQr3+VjqdRrlxx5fM+soyjFZE1mF
7wJxb2uUlcAAZYPS6lKJQnKlXv9lCRmx8WZ10H/c1o3GLEho4FuIdlnJBo5xSzvQ
Ry8sfDhU57N9B5t4N42nspcrcuRXTocau8dZcSC7EVUFlldBtNIE9XRxawhdKb55
I5f1RsNOEfxLBdMMmov1L3bLsr4TDyQ6WTKefBDgEr5J7CK9bgnBj0HSdIYoNPut
JguHWx2YoD2dCR0ydxUDr2ItNJGxVPlACQhs0uDfehdvknk+aJs0Tv4/SXm2SonH
xGmPAWRje21yAy9baZqJetXgjzZeNrzPKXTnJm5CnytFS9195uKzT1FJtsk8oxCK
dhWbe5nP2GU/CUwZJkn1G2J64WOLfYeJEY0ERcnh/rXlucYjRXbV2bnv0rPD5FRy
Ddsj494/nnYxxnIO8/toBFu0+HLtRDHvHs/RStOipFPyXxuTNzRsj2LMr0cIxEOc
15xIOSWnAzT7M9AaGfKq/Aks92oBLA3osrV84ZFRRrv7cZoUrp2pSgjWQdyEeor3
z1DbaQzPj7iwiqtlbLMnkNt9EdR64rv/fQNzBi73WkhouUoKs7LUvf0v8/VD69pb
wayzEWXn0+5CpQNQAou7YC10utfVnqtkbtsXxDj5EtDQhx3frEn7IMtx1LoNRnB+
WB/GUwXGt+sfhPOkIOfLhYyT6GjgOFyGD3EuQDk9EY5zkBm+/2ubdy74PPia3NZj
C7OaN0l91V1GEhgJnrV3EcMYB5+HgY4ZXn27Xl1Nykq/3abtzx+PpXizD8T3LPWZ
/nj/x3B7Tejmys9ltHtczddmkc+1c9PrO2tWWxqm3fqBX9FEb8k40CmK72bb3Ai0
9vp6e4+5SG7wFqOw/7fkZEJUp+1YOKwhSn6aV01DC3p4uCHL4RVIZd0G9dZ56ZT0
z1zS47GbOsB55ZgQDFKespeaZoaK1nGXJLnV8JQbFfTDQknOYmBlm5aYNHzbfEtS
AA4oL0a2ZEpoUVBjxIStYXBNpU2FXSecKaKb8TSZrJrInX3wOLPdozI4DFmD3Hhi
1i5wrAmpINdNpR581WFTtHLMBvuANAIcglqLqmmP8OGv2lBWvJiWe4zLhmpZVjxZ
j9iPnV2EuH1zGtAvKFTg0stDliZSrmlRDygIW2gkWbdLkHXJPevZJPJCgzNTRBCb
gLp0RsFCNLnqr3d1u6PYhHfutofMegOIoy0HEc11GQQcWIbSfWuNem8cYiYor0rc
JADTaraBl/3hbaZpWNyo9q+bNkQz17pT6+EXjGIgcFqmHjO+myahwYBsrtbcmj8o
CxmMRbHdR90cM6D19uWvnkEc3hTsoAbhJ+Ncyk+oXc4GSdBWDy2EjcrJAkm1PQ12
aGrV+lE9I6auzyBbcCGQBkL59bM0LuEVMoo+0PdKXWuKlTwcnqB0HLLqv6GsLTYA
ubADuP492axQkW68p67zqo405xcMXZ1v7znzEktNewG+TT0oDHEFGlG+HwBK/6o9
R6m+H/b1lj/jKt3BXbb3HLqAHM2scVcnU/thWR/Q2/SF7J9ZbTeeyJfeUF+nAGRz
FKxI75reAzgcDMjilyswdNC3F9fdJ3E+4lGL/b0VjzB+yqA9fh0UVeRQ4GrqllJk
df/NXhaWUC6d+Y8TAx+Vn4viCrFvymA+ksEjBsJInhXg/RwxCZUeoswD2MkIvjXB
5HVHgPWB5pJAKYfwvfm8UJ52tsZvT7fgKplxVJ31kATXql6fKi3srXdUr6Tqr30i
noU+DbzlcKf8iMPIi/J3z6V3TcF719LuDD5Id24IkGVXsCTNpJod8pxQ73s00tZz
bgpuLqN5WZBCmxDiwGTw4kJPjNZydHm72TlbRWj++e7aRi5YeXAE8fL9vvRRGhy8
EaIe3YL0GBQsEIFu890YkcdiB8aTwvwA3In/JLF5KqNDVVrf8Ub8yj8MCVr+ALtt
hXOSu896wPN4F/dfnAvdypj7H2VgtWcio01eb/YgiLlNka19wH53JRBpGbJUxnF7
edU5HjVMGg16eOJTnOQEeVF0jy7Pv40xnA/iUkySDB9dd1MTzPUzRDRsdbp1+HYc
anuXLyhcdJlWL5Zt+uk6lcGokhYUZCKbzzUAJu00otBCOEG2ryW4Vv2jlBSg2E+T
jGTr9LNIx5jyAkU9MlYi+PMMuQCTPjDMxKxavYIUHpMVTPZAMC0KKvo/HK8g7bIG
KIz8GfeMwGibMf794Q2rJIGzGZNf1VPph4qHVXbnJn8z6WMPSyAbAoI07499VhHx
t1H5LiuWC/lH45keBkggcFMfBzkQH9IhaAkf/wsPZrGK7UUP1W44y9Rd59xvQXLV
9qj5JsJtbjy4ixcNqXDWRE7u4sTw/F5NDht4onqi1fK+zLzg/NPMl0shLmn3tEXC
LQfWZRKWWBo0zutzSs4s6C8QHthSCZsXRIvMdPVbbuBX+GVjcfWXogaVqzj/a347
wYRF1RmSDvJejxKLyPrpVFBf0HSlUEXkv5kxmdYdWyvVA6ZE7Rvf6CYzYK02yibr
KkRicSdyyaXFb6Ci1Rs6qD4sbHmquB6V6b9WC9hbb/Yzz+Sv/ROkuf6UZr3P5YH3
+qGtbb1y16ogD6Rl6MbxWS4004uVvEHQGWjeFCghEbaZS4DWCxPRgVpq33hx9GuQ
1Ad4HGMdY6hz8Bp6Mb73YMdyFCcJFdchwTD9JR8qFFzdTGYn5FVddEAcuO5jMPIJ
pCwLXyEyWznD1E7bsUsPMsCHjdP5pO1MuETYD++Pygc9dc5YJGCnLxOWtWa9IwGW
Qcj6djmNH+uG8wMOPxU+e2aoSB6trkuF0pYS7sh07/hIFnKl02MwtJnjkyaBRrfd
eBFu8KrPmte3mzeZlTSbh/fCvcRHcYSppXrOLs1XdVeP8nv5qUAj2o5HPegeJ2dc
ifjRhPfojAqfSvQ2nChnuq4cVPMCdJJz+s/ORVhjfY73Sj38HZ15oK7gYNAgPsSN
10FJUx/Et2oTyN5v1fTX475OkeCR5IEY31vI6iUEQtcZSUCObtHEy2ZRGtKvyB/0
oQfrOW9KL5El4lvRCCBxkbg6K4jDA0HRFk2qgWY76XOQ1tu62ZNuqgA8xl6QsGMa
E4N39qrfc7U+93CiqawxKE443ATlJiVBzI7qcFNruPkdd09e52XOABm7lrHKt6+b
mxLjxxGiPgFSX0ygeImoDuQBEJMGMHFwdfp5r0EgM1s3yms4OOcQ/BgxenKt0qRy
r7eLFeVd4g3IYj5TM4+dtXyUy6uT4N7o1Gr0oerxULPaXKI60YquPnsKTNe+r7k7
ge+eZAX7Pxi9ncIOXhRUHgmXJtPfeLGxqkE28qIEEWHFFhenCR15TTP3gotyXQY3
j2g5K3LEPFVrJPmeD6xDBQyFjjNhTWDe2Rog1zNI8YKaxH4/p4uZ/Ib9tcPzQYm0
Nhclmt3uiKghaRliyimAsaEMKx80Tl2er3brNfClDv8STwm48sKvRl+52K9Kw6HU
2lGtpj1lkwULIxWTy04f6aBT4eaee5ImAGvIktOwkTPDl0nJb8jqKx6AuZDJLo9O
OZnO/k2YGaOLqyRO2ixeEgjhMI1PDBAVNONwLeVuH/yZNLzO9HRQ6Djc9bXRyUlv
bGnFKi5+LWfDgnVmUhAxrbRe4z2GiQgWX4p265KKtXQRGkWJI3RI3OB8LzWw+bHh
5faH6iDeObMstdZp4A5rmFGlM65w2dptyYNo+8N8diFHEl5pHloRUp9b/EVQ5sVM
Earjawa+sB2SJ6RPV+2UrtDaYw2voAOHIZWWLLX43N/mBv/phe9GXEehnb9kqnCu
jET9655JnAvO9iZu2ZuotXe64DeVSAVvBQub+yZAzqPFoA39pRnyepkiTCvmGTE5
qfmB3a/oqa4rBXPg6bJ6fg/iQV/ID64TvmTHPOKnQy7t7iffyUWIsa0iCo6gCHyv
6FxwM+J7uZveq7172JJ8tx9qdZ/OyleMMmA5uELesbLD4wgu0LSaL4XmJpz8bP8D
kNFAxjmMVi0RculpeR/o+nmdWM5MNx2ytPq6eNV7WgR+ncJ+t8OtHZUzAMcxwVCh
nJkqKjMLBhTEWXD1s1cytQawb8NpEBK72BU83r+vS/N8TqRICCnpypAKXLQbDvTG
xGZrWLI/iAVJyU2wWLCI6LfN3gy4IwRzIsUQp1pFBLfabPfMs6BPSJcqNt+DPfNL
y32lNnbcBR7IjcKBdC7MvRgepgWkbiZi0neXjL0bRtN/N+j3TMKmel37oPzNCHbB
dfkMTQMvBfdnStLfuhq1Fgg/yme4KBwN/HD1P7YMKbVyJI71YSa8I9fDCQP2Omlj
SIoHmiNGHRrfeNmDEyyrKp97Z1UM2Ph7n3fPn8FE1VUvVl3tDYTmJYwIWw2yqFv9
+oYAdiOYskZBVP25aZPuAu3sZzs8LRhpODaM/Q4lJuobMNZq4vcT/qnJ4pytL1B7
POqg9yY/2H040SW/Obpx4sJ29r0O2O77xRtYYCr/z1mbGF3t7xan+4bfoo08yxis
Sb4uwXU5IUqduMeMLbxDAuZoS9jh8xulwoA5OzaHcMt60vAlgARkYT4FnFaPnSQw
qt3J+AZiL1g8H7oMZsum8IBAT6b8oRqKSoeXrt6Hfnw8WANIYQ4QAtQsaH04fzgB
nK/HirkdyVbGdW67Bu7DUj0IKB3kjymxJ4pVx9HxXIh5VRuaV9a1p6fk9BjgtwaY
kwPGR3gsciODOHbqBpaeELBnS+BIUrxLRZP8GeViyRhdhgeVUVRTU3SZ4lyUEtfl
2ZGZMaV7GK9+lXo3GXYa7TX9OMvK1t+uDmw3bDj8sPks1o++2eWU8fmSJni9cOwJ
QdtoKxOB4yIZr+5i174vD+Y8c1ZguKHSTP6qQllHv3xYlEcJGJs3jUINP61mH9F/
ixUICAEwZ1wuukdw/beyimIdMaY+LlZFIJq8xxKgl27QBt3WDWTRZPd14wBfIP/V
P/V+eoDefUTfrNtOzaWJxr60nk3GO5D2tJtq1ZmlnrTvsJE/ir/zNhDI/a41ztJz
50k3zjmJmAJ5vDka0SlzWGR6SBUf/lSFqeNBcbOglpRK87rIN1sDzWHhcDk66qs2
HLuFNKqq5Xm7jgTmJWC/zlUm0r0FDQylVlm2hBnzVXxefPauqtV7kqm02VsffhJy
oCfNegPcZZ0LQ1lchSfss2IYb564WWJNxl4lta+qvpSOLzhrCw6qnCE0EZ4lfXH5
kEiQS6cR7oqe4gev6MRxS+Gzf8hBgcNShqr5eGdsVGK6HvQ1suV3Kzb4d/9QuBOB
sM91m0ljO5RzA8l1Dw+SiJsikUABh4hHowl/9Bfut4lHKjtkzEWuEjU+9Srh+fi9
Po7Uqa3SvoXo2J/HWbQlFfxnSkkcUTJMmzBM9W9I8Oh2tc5tlGWZG73G2zq1BQix
3CPvitMiA8ju5gJXjVot0/i4fjUd8ghicv6sl3WcvoD1ZkugPnUn+SBzDPQ0qTeU
cr3o/uR2fUcbT1GLb150AHT4VDaI/RJlHgco1nb0PDO0YYE9zFYO3Hi+YyjtURfN
MmAA9dgWp5p6Z3uuuEzBirjtIPdD+ZEULg8kFjVrpt74BwG2q9P0Mq2SW0Oh09br
oTSmk6zu3H6RE9ut14HFmbIdVPgrP3CoDxj+KOZdBjnrOASiCTGyRpRFO5CJ+mdS
Ange+U/THqiLK4xCRUhvnN5rwNZquTFPufQz1Rr9y5GnboNtwUbtOrGj18pvDg31
5yI4Ner/Iv10CeiAnkDhsWZQdlbbYPcXMnHLcfkCT06yr2xhp3ecR5yCmEJugMQ8
FIkn9VZKzECs8JdX62sNHw0IYOVXu05C+zqKWcJwPQ/VmmsKc4nUvfVjG/Gg7ghy
jpP3SWl292G3K70iU3LnrYT1ztidbNspOmWHKzGEXD3uLV+JIVmcLNoP5N9UMP5X
qp5y2qVAWQMd7thwNHK38acnT2aVTD3mckfsu5HDGAZA/7WUrC47P9Z1qEIBGnP8
6hWam8HxT8roYi+D8PkUGen15ChnKNmVwQ7obaUPxVq1qH4ToJu7pNH39JMsAWoa
a+JxwrLAEZvqokpAv96orbN9Q8aDszYqaeV5ybLiPEYXGtFzalmZ5edt6TQ29i2x
4a4pWsRUtUaiulJ6IJrE5lTpjYX+Fk2pxbZHv9yco1m524FgjipPHm1c729I7IXH
di8HBkzKANT1SUG4gfyS6RISKD7jHVyfk7RexDTFFZJEZsS8qqxCvsvGOKCOR184
yZ3Ap0e9awnEGkkRYG5mJahiq6CdealbMLA79gzclk20mApZhu7yxCW2QiTB+827
CTGk4MerkmPzCDUy0BJ0haSiBSzZkn1u9QqGbTbpwOOT1Gc92Rpda3g/Fb4W4rn7
2vId3RTxxLvALTSD+TPkP0Oh84zpCVHjyHLFwFM5XiDiMinvwvFjUlG0XpbEUuev
BZy6hvzXouzWrecSnUU5SrZfL4HWbBGW7G5Fu9SMvzB1u9c4g95mfGwb0nsVPDCd
5azHHorV8bnn2Udby7y61xcRqgJKpzLzNLBWgS4BdTnQLPcI9u5NfH0hxtsLVQ2d
yu1ugBb1fW01xiOPmWXlaoMcwZsH147/vc4Ve9uxAd7+fkBh3vv5QiSU1u/Fh7N8
QcEEBFj3DKjqlhqLZFRJClOGcEoPtvyjiilHfh8C3izOqBWWrSjT0wncruCkysMy
Ee8XlwHT3SrugnLXt5a2/bbDB9hkMqnxrKloOi44eH+4c+fKssst/LtMD1WWRSj5
1UpOlb4Fw4KOI/GB7lQhVbmCJOyJErZ1wAK68AncBvqiOmVIU22OlyqhZ9hd4YB3
uO4gRc8qNVS6WZ/ggiWfm8eTzEebYQcjlXyMxD6H2HXrfEE3pPp0EOhCa6MD+KUk
RkTYTpXfnLv69xE/eH9BBs1QpzRIDzXspTk0UPzfnW7SSBR4JSwE8l22gtBF9+aV
d2qPTASH8350HSuHqZpMSZGRb95m+9eJAcb65KJYttZOv7ilyxEofTt/OdaCGiAG
M4IJEhYUIdruULLgV/43hN1aokW0hMoPCDB1YNgCbtz8NqfEmWKcz9OMPIINgdfZ
AiMRq6MJSrxQ55mLK19WwdOQtxsN2E7pQXaWh1r3V+5i0ULJ4FP+7eQhHnVEuYqa
BDykmqjKSPe8aw7KE1dI8qgloWUrNbQL1Ki1sfNgncAq8NGYffttM4FPFcCwFpOD
rhyq+rxLrGaN0rq/LDUyxUsg+r6omDDKsxHGXI7Ify4pvQ3cC6K0RQpGcljgPyWq
iQ+7jNNJbQCcpOQsE6WHtSbjJ8k7CTheTTQv6BAlZn57q5yWxxSx28J/MazTDRC9
nXDnJcXMx0YEFo5gGl7AlwUzEkO9cYOIuAwPgg61MlsR+nNGlINU/vA/IuOboJ0W
fQ53SgoiNDFISyD2QWM6mWUtEVAetB2U3ETCzA9csxBVv3nGr4rEDhzttEUcOjXr
xYQ8XjEAUYO5jpDFdBPQaSWXgW6jSnM9rfRDx1s50llclyKzJcAZCzx56AzgkF1j
EmKGSUA3oaYX+uWFuGiKa+lOkVxh/tzDGgYwAyMS06hVldoTq3tcLW9fCkY+d6uY
XbA3uEs2cEhujnShrL56/haUruRvbPUMtFTP4e3BrsTx34BP3ak9otfSuY86toTZ
8cbA7q6d3YbESpbin3p3zL9mHtFNBIV1nIa6LSH/wljB8fkiern056OjSTpYlO5l
TZ0ML8jNcpRWvj/Z5gjgHjWc1hQJMxsmOTypD9G82Pu7Hb2ZM586k2do8Pouoq1Z
5AZ+Mj8vMsWvvUstC7UvCSsyGmcx1GCtU3AxEoV7DwyKWkZeeCXfXX7ysIJLhvoc
eInkcFDvTl3Bgzz4EXkEVnGxCBd6IsvDdBPXmy4jNXXoIqQovGJD8iSYJM/g8Ur8
2sMQYHoZ4Vftkka/WXSvBDTlNKNe7XebvQ2jVeThDrCHbKLCUgpwgMPafoyaeWwT
5W2Q4YMH4g9adwjub4cpQLgYRRYQ1S2hXkV2wTaY5tvgCWWEglzeZrCjVwK6FfhJ
b+0TfHMAmD899D3OriNB5xedAbmoJr5stdrHzxd65VgMTTFMCJs3CMm5BFQgoaRO
1lXPsaHKW4YRMN+vw0ykonwzA82YsiXaboPqMuAb/yLYmBM/eYyfKpengJqj2sxh
mffJNg1QWj4JRWLYZBs26ymoXp4lcplKJgSqyXXfrsb2pI7KzIwOoNbRau9f/5lr
Jrv+BjrsmYS0QAtNOwGQLHWbQbnkw5zrVdn4zVTmCGuCAHxzPa2mt92aVCO5PxLj
8RM9YsUTgQ/vFb/io92sfFHq6yCzTv8tOPUS4c1bLr1QNEU0c2R5NLj1Ug3WrebS
3c9TlqWBaA+efUll5187TDMdzUc7vZRZgFkN1ZAW4gXWqDiOcRnfXwrdjwL+8hPu
+Yz46ZYBRtyNHd/VmA8ep9yA31LeYXGPtWHP6KPsxFJ95eeEVtLA5vfd1IxAoU+R
1xLSQBey7Hu3ABZpGcoM4MXzKjLzS3MlM67301ct/W7W5M9Pj1Gb40FgGaluK/Wb
GC41ihx1umFjNOIyNgHxBk2VVPgrYck+5hv/EY9StLf4sYuyudeyMmg0VNkE0uqq
TVO8UXaX5De5GG0UICxYS1n0lYepw3DrHlQiT09QWcuqude61UGAZw/ko8LFsyGx
hkwrVdUI2OYAh4HRMZx+JKNDa1YnEanSxREpqVHylpbtCL50oiDgUh3wIwWQCjLM
q1WCX0titq4SWuUGf/4rgsEEFZI41cqu/ISY5bxrs79ocN4J5rnN9ejVCwpwNZij
vTjk9JM0lIuKVA8275ZsrmM9lYaQXukkhlhiFjTwgNnUD4BdpsifuTkir6Sn/+I/
2u46Eh+ht1jbUTFJlpYnY+6Tzoy8hRwNHEwMBSsd0q/lgatkcljv/Qa/wm1N+jXn
40ohP6127VbQur/8M7NBrCz68Aj1vg9n1PFee8XaK8VLObElreJWrIu8WXgh6SHs
IpcrU3/S7ikBsB+dB0ck5AmD7oWUdRfNvBu6kTuEa3Lx4BuCdf0jZuEOW+/fjVs3
GcnXX+5m3RPTaAQ8jmDDjQH8FJMXwxJKswcvFFQ/uQ4nyKPF6mOyyAUnLyeyzd9H
KuHxI5PikGog4os9EDOeiYgzJlaP5CicJUilQ5RAIqIEZX0j9+Auv2Cl69I+a8Bv
cv/FGlYWKRiCP6f2cDdNr9NRPxXpWXQJYVLtB2n8VElqty9ltARucrv7IRgA/ykz
Ri8PqDZ+vR7DUDhSVyx5y7JoYSIDu4K0Fn9nb6940J0j49Ntswp2/DJ71QvwyzBo
byPPBooTdiOWcCL4vdajeTtr8JRNcWluoURaTZ5d8xtfHkb3dcikISxTava244M/
XriWygiLDnMgTtA1GPCSd4shkm876eSE1rw7QmTROhWT1KltnfPnKq4ceslMQQbY
q8x2vlF33d1qMpOwzH8feoHmbtyUKTIKl3GLbtc/q+fxDVhvq3amXIYNU/AIJmej
VCp4fDqJ0DK1QqgZ+z1X81Qkb07Q4z2IeaDbSjip2jods1/nKVu6livqOQJIJGR/
6Y84vma8s0sjvkYwPykc+/LheqlShlFGlOH3ekuyTWgUIMX9GDl7DZ9S5C8JkQUE
BNUS05s7bkr4ulmBWZQAY5ZzJxhXl4iKLz/5yuhj4YYRGh6BHAiIEWYs6tKCny3Q
SZw8g3Ldco6PesOFL4dRdnY3aaWNWka3IOy+Ip5dsfTXV+A/pWqMoNPE6TvBW9h3
puajvhsxSGtPW7k3HyieXOCqiqpuJPotGSwhlnDkpi+zqvWSeag9i0zdyKX0iCUE
6IdzRTxYALWVMGrpeMGigHoJ8ql59aCOgEmSYjBL+hwG4UOaoD9ZnKv6/YUFQyMQ
Q7ByMD97f1R3tlUV2wdJq5dqpm+8U7vKuFrKsMrHTva/aP9gqbLSJw9ie7/QO7uH
OnQr7OiDihdsdMaQDIm+YRmi0ln0NKNWgezopqVrSsfltTcfy2MW8GeD+ej0uazE
gk+D+P2SSFj4LJtwBnHUSPK8ag2BEUbo5fDcEEteUwXQb9LUHUk6/ClKIW3wVE9l
o+d27AsMaaf1UFJ5cijz3oYzYYyLx5IAJUyul6Bnlbkv4bcCOPz2KpVdDSjJQ4N/
w1N59Vwjgbo5oacceH8bRd1SpgsR88k/1jB69JHtyXsq1seNPWRHcqJuwDkuqCGd
pzVToyF4JdV5rXSqdKiFxasoFeJWn8A+ChC9lmZWvn7SYOsA+czcr0aggkYMFbZ8
NPjDl0gxyYuwo6Hbra9+NnCu6l2tPaAguVGLVx/pnHRryxcxvvL7I6+R4CevwASA
dK6PYrgQLfvZeWq/XWWeXL4JYqCTqI3EtRRFkJbQwr1T2gJsgsptSC32V2nvgwTf
J4m/kC9MaIwP7jDM6r2RkJ7lmaZwLiNm942twl4OVd2m3G28BUcxzHnoIEonVwKA
/sd70o6k6vA+PUo+Suv02cWdwUtXeB29Z7uVxLMWFz0y1Yy5vNbME7SoRDo2YXtv
K6HkyJCLWR7ol9lZKpicugpUYDF5n+KWhgF5vNCFlYj1LabALXA3ZrgxROfi2EUG
8l2sqtiffd8LPMce63/4IZ24vnIu+CrAieLLiqkxrHbZ/ZxoTQblTDPHlX9UQJXa
avp766j/ggNnbHE7VcKvBUCvNX5i22S6XeWRIBgEm/paV1NdxafEL1ij0sFC3eD9
x09DCQd4FYsZX6cOBiDSBMYPB0dz4/YSM8enq9pXL4LQZokqeag/ENFX7meNoRtO
LtJkzLGHk/KcPjZBcm2YHtccNarWf5hq93Z09ENnu/UxtKY5mAZ+EANiuhecDHF8
wXsWznr42Vz19xY4/4T/dCZDJYEtwJh6Ks1VqdYzVYsD20vGA4lmKxyXeJs50G0f
lS/A7mNEN65kACPndnjbygqHuVzadDOzlstJg0VLakcPbc4RHuMrvWlEvd5Ic+FR
WclZVoI7qpaaa/vmgmwfRuesfs2l0tRoasg+vEmFru+0kj/TDZEzVypkC5PSntYd
yy39cwi03765UEYJzjzwNcRPrOYHsyMv6YOsyvfBGDHd92AG9lx7AP5A1ASuD5Me
zjqkSI18iO3ynVHt8acxZu8yVjMy9WjnYPADW8K6aNRtrItzA9VLl+aqKyHgvCAm
hJUY230RdXwI1HdMI1QhyRjs0zLsYPYknPB7b5mXiw8zvyxvONlT2wyIDyFCJ40h
J7VmbNeMUZ2JZ6eCz9s5aPjU0a6nSvsltyonDpI99YneH4H1v9nQ6wUArZcnTcdI
6L+NnUssvydZs/P1P3dQOH0ddGPtFYKog2vYrq3KJqXVAU2PkoBkdmC4+tgcy6lf
cFSMzKLPZoon7DHM3vw47b3fX+S7ah1rm5uPkswX+NhIhVX4dLRAQFitIDLNkJKv
Ia+BmAV8DjoSS4DgcMR4sup7r6T1wbQ2w8/1nfZy0XSl/83PxB5RoAmtvSTj7vq2
2zgIwe5YGwOSv4fQaQAKd35aFr4hV4ap1INDJ/3lfkPilipmAjWVpUFbXGyAApsn
Aona074w7ZEHaq1Q3Q++gPXkaPn6sH97cxSvH2DjimvUAiOtv+qWaHg4X20Ib5dx
h3uoGOhsqxvr2oo0uqohSmBUGhuayqxlMYVCEtWdW7xbpn3EQ1g+Z+qY848jJP27
dxPP98aVszXn3qHkWCWg5V8KRQlWoGUZns6bVGsyOttb2rHkTsnUgMVYyHJnA40U
6/R46Hna9n9q5YueSYhEkakhitLkqrBsbY2IF1ma2iZg70T0VvBj3G8g4RwPIsiO
JxCfapzzEvHO+A8KBjUOPF3frJdWFgSwlsemiXb6nHEXI+8ahhBgehpyMVSsMs6i
bBPmIn2QflVbqDN2z6i1Y6raEepmA+WHAe7NcePTgJIfcSZ+/6FtE6Clnf1mUFOo
o0H6/2tVzY1hhrA9giGMQu6STPORlxIJer0tof8Rlnhb4s7s8EA0Jxhy/P2i5S84
gzgrru/3dN9KQ2z/7lMTIOe45mgixpESoIIjLZi1zWHJ+12/clHZabDzCTiKveWO
u11uid1gOcAq2jQfYatEqb15GUTgzml9wewElzNJ2rkGDiTs60B89ciu2x4TQsDh
jUIFfVj0F4238CBOIHQF5xP6OJl9aSP8zKekKIfdte+zv0CK9UPZgNJsKU7wAdpX
eQQbV2xyzcNixTXJN4QqRky0ahRSIhvQE8mIcXr51aK96SYB/iMQDSuyWRLnETHI
4aYiz9JFazktWTev4j6ZLh6gm1LdJ7Njy69rqx9+8Z07WdWR/1PmHmDrv8icDnQG
U7JASl7weLqcCYrWotvs8nmKrjPhdVUeVRDsduR+5ZaFXtUNPhWJ9S/cmbj31iYF
uTauMDIa41wKdENdYfJUHIsXd3VyKnn3NFvjoqzzBdJp2tunT1fXxdjUKMzmJnb7
a+Iy6wZPLL42YIuWluQBoorKbumfLThDmeJpUG9fFnWu5pOr0NaaSBZGVjp6yFcy
yM7jRR6GOh8NGEoi9/q/F6GJWqKJaCZ1uATYKwfAwAdz6hbTZnd/euCiQwwdG0Tr
vu3c2hKJKxOltejbZoGyScVL6MFclL9F7RO0hxwlJ+y1j+VKWKsB5yYUJ46X57Rg
cgAtya4ncaile/Hr2CqyFLc02kTk43ZR7dhYuoonMiTw+D2Ie4KS78lubMwg1WMH
UPHfjw4zYn+OQL5nmyTe0QitI0Ycvxllygyj/WW7GertDhZ5SaiC6NNRuJJuZAtP
cZ7W2Yis+XIw0k1ONHM4EZ4VIyDw2zhIL9AP2gsyjASugOvRm5XR9fSF3o8xf9Tj
ZbPikBrMGoxurSvua81jMobrZkP52Hhn0jQql8vDy49xsXZehqCnFs+xTmrKNc6u
7AKAsPryvLXGFypMqgXBjywGUR1L9fH6C2gQAxXYGRSMGq12Dn27tFoFSJYWmb04
HVHUiSRDYsvYmpEDf3L+uAqSII2WX+XUGBbVagzHrpaK/wuEqk92fhMxzsR3vUfN
sOL3NBGANNCxTsaFANX7T2paNSBBgrGu77Dpu6YWijBgqRgRJIYYmfDLKSieDwBf
k3iit79RYWDWnlwIF9kekL7cQOXUNn91Gapgw7UPE+NZ4vkLXNaf9awdJkYhUNpg
jlyhKTIIprIvzNmgYvg3hMU9IeYWJe/1i5rmxzfRCAsf4QSkuTovzPW+SgUOEIjK
PGEx90Uv7EQK+/RySyOpcMPpbIcCvA2PH+3tX0QMHIbbuCDqAstIFVVXw2VwMFj5
8PLKP5TKItGoGgY+3uarm5NFyVAGAGMJPskIUMG4VdByLWK99+ZxHDRzT2mAYraZ
GGbGVkFt+VP5c8HMrlrxCXl3RtJf9zIrYqv4z2aea0RgrVm+f4UAL9rW4nUXOtKE
ZNQOoy+zvhxo0byVNCng84RcqvbxAQHKYLxcHEMRGUmQFRnO5+bGZOEMkVd3NlEu
fhGojp2vHLkDPs9Pa1Zsyxs5ssGw5o5/HsfBy54UH1yNMf5/ZtArTHb5NHhHitWl
1MREtibI2wNaRWvPCb83ffyevstGbe997yYbVzaIB8m7HVYmtzOqB7cC9pe4QR3W
BKfSMLKJyClda3ZQtKhyyMF69kciT4J3cb+kRvmi5oQzyLpIyKxHZ6VNYyt3t3Jq
qXICkX3Ny7MamEAiWOJ16jxxNU0Que9aAXao4BJScTjZEavRjRg2q0Qp/ukW3BP8
amTpc6EUidjQ50mBpUEXjv1LKXyJce4qKO8+ZsBwHuDXW77QJjEHfhN9UwJMmrOB
yZsPg2E01JG+FIX2tzAL37p4ziK+dyOAFWjyeZVBos6kHQfOTrfU8Sqmbn3tPmn5
fszUPdDkwLKSwCyiMI7Ai6zN4e/iHevA3NlFdfAjb214sJexUm0Wq+3GzUOlcAwf
eeYgOVdOcQNwXa2IJ31uypEqB6QUwh+vc3V7Uing5weeG4BECphWL/Y/LxIwHh22
28Ptqc5Aidy5t/wDY/diQx4Z3s4fmc966APMNqF/J1hlYgPn2oarXku+34nnH9n2
UUhi9Xav9UKcZMQ4cdVh3SGIXKwLJn8NG79fpUDExkapImXlYdODCS1XP3lBEg3o
esLFVfbfYGtcbd6b6DMhngwVfQxV9ZRRMybFnvUGJATXjDFlWeMUw5dvH7Z5p6Gf
kc/Lfn3HJYyAVZTM7ODkq5EpRgO8Sdfy653ogLT9NTQ7dNkqXNtkKQ37lGV7s8Ax
McNw8kmmNzAJRaV+G4KAE9c9CwD7GMCyUfB0kclp6XFsHcZwiDhNl+bmPxqKLuNC
kCla+OA9Touj0IUEWgESqwl2mxQf21kkdRRzntSdfl8l+0QEYMa0FF9WcLGcUxn0
pKIYw6+qw3KZ5lQOrTKbvdg/I4JWULZh0yFmyY+pPAQjuaKQX51+RQiHqJ87zuZy
hDcTmI/bz9b6vDGFlFKGnDWg6hFmug85c/Nz8rtY27PV+Bb2lw+NbBZhsI3WIUQG
2AIxPvvv6rd+23k80PeqdX1KNexJ+xnnGZQK5OGBTA4dcDsdC8f2d8DR8DYr/yxp
u9hPg5IinoNCDGl4RhgufA8drU/MBTnfeL75fQOD/q9O9UnqSWVmXNv2N+Qdkksk
exW1YkRD/8Lx9+nnQeyK211jJzMJZ29YjL7gdXfOA5LoSrRwIoHtcOrlxZ0P5060
NiiEGRA9H2oCkUSnfe+SMH7i8SHcZ3QTZf6QuoprIDN7qgHteveRpZe3NPoTO58h
MTA51abGe2zDVK6FTKo666pdOQ7YupSHhfVJSeEozDv9RqSZYZ327c01DGLllFBg
WoKh8waTpBwak+2nye8JX7JfFOIGHnIRV8ijKiPySvrfltUho8y/dTKVz5PM31vZ
wtqIWj39GUGs1JWnZjSxUC7HdiUjSIc33a10iog7mcF7fBi7nmJUR0qBfh4hye2Q
joplle/KiywvNSYAePuUsUTj9eqEFMeXi5bSWBHzYBnQOKT0mNpwAzaP79c2SJWf
c0mOarBsLm2goDz6QeeVWzz/wxa54E1MBThpMStjlp/jJUY/2MAgWl3w3FKesxeu
BYGde3yJb+NC1yJ27GltKvJWeor42/zdER6uWiPBNbNUmHnIdYujktF10nhYA/Qv
ZqPvDxNWbgSU8cxwUcgukZwqQ4A5RFim6amZWeQNw4pO/9+d10TIXlkAlCDTRVDk
dQirgZdkAUM2b3e9H5tfsnElY5ok4CRnspYkex6WA0HhGJReH/Y29UApQhYi4HsT
8FlyYJ3Ub5wTVoligjKSSleCzAlxTVkWxy4rt7HoFq3HgZ5X20InFZZrrpw1Wlyu
wSpPpg8LFepq2hxxgF/aepDwKmmIv2qMnEccp3zeZeSF2ydTqiEyjRWbMKDfHf62
fM+1HR12lyhpnjEpYhjOFzg6i8dAA3wO/n2Yu3OiC2vPHTvrDCdwRw2dYfslzhP8
Ym+20759GPQFqc/7ytBQ/lUW+n1KHeinfaPDg+zp+vquB6E3XjO26fCSbVy9h6YO
dFd8aNIRFzCBIXpeHw7/pQElN7E7oSUUWn0opZTKTcqzv4FuETCM6SXvFZxDvJAN
QF5hWO2So38rt5H/oR/UlbBP6UEzR9itEF2cj4QSp38Z295kd5LZE2sqwRgAJHh7
KL/lpioGOEja0UTsmPbg+Jyt73r4FzblL5Oa4CZo6enP/UUCFKFB9HCZ8PJTYmV/
xVRI8x+3qfzebYSmASm1vAbANsYH0+DD2r5rf90eDnjl2IqiM2557nkBkdMClT1J
NasNt4ntDYiv4Y9oadWMd8p4ew/gFiolW8O35yOdDnCkTDha6pU9KIyWVMBWDWI1
DRYvO9hwTmtJFFlkR7AtYXyvjN3A8ITvEKadtIvJVBqzDhxcLtXNpBPRn0JDRpOq
CpCizB8tBIDRq+HW149+BCD0QK7fln8tCbc2USUMLG8i2we1Uvw3lwuzRPWPsS/k
id15hWiazMIW+eA4wpFWi9hmGYPbPGRmxZXmIki/TCcS9zgI2fI/awEgInXn6Ij5
D3UHn0Ju1rjrcO/DVaHtUzwvU58W5EiN1P1w4vPQAymz4olqqmMgj/PZtxm4KNIx
Bc1eWyUKY61Ky+H76Lv71PBDOLGOpWHqG/1+RH9rxNkh8EzJf7+1gdGKYrFsZO2y
nkRDcYJ7w1D50KfTOTpLEcUU3vwc+iuJAc4nfIYltwb0d0qNWsYVl9UeA+Apg7Tm
w4qjCs98Cx/oDbrZsg251C+h8JAapG1z5ax7oDB5A1EdctVOyMSH7+NxLZJ2+i7N
Od8Y7NG4bCEw7szZxIPpIRgYt1KnVlTIa2ohsnTMbFK2Isx1RKMGG7Qrd16A7O5v
O+MEYtH3b7Sd3fHKtLa+tNxddQ+GRlWhnmBq+R3ddCDeOr3BLU+NajqwjvKUivmK
e6cAoDXvlESx90SBwuZahq0ZAlN/tQD6V6kR8wkmVher98rRKAjQmReIUlPJyeik
uunt0H20+ySP/7WVD+PPSosFMmFTix/u8G3BoB3kKeQdtjYKfdjEQvsYUARDMDLk
ausqQHddwDTkMYYzu+mNPvk5/GfLVcsF0p3/wnUw/ukwwurXpSgz8G8Mnb61zZz1
GVarwQg+4qWPRAnRDFRSGNdfFdOrjuw/OqZ1TiKnIcx/UaRfyqbCjFSjlJfZlHtX
z+vaDDj+tX9GGTCWCJEp3m7JJ03Sy4yVnvZ7DUN0YhBCxZfUilY9ATWA1TaHKFOB
Lf8xXU3adRaLj+pSHm1IEGlhPcC5Huty/YUAHjhX+DefA59p+my/q6oVSXvXzh6T
crz5+OW9Ww+SO/c2nvdDkbhRB/+3NkLn05IVHDQHIx0d8POehms6H64KnpW4hWvp
iEnYQzW3P4y/G1UoBaWAR2fHkTzao013l2AtRV4osRnOHgD/1xJzX4shTA9EXArW
3lVr3wMeYsw1LS5PiKl9a7WXhylMQLJ/z4MkFa8zsEkvOltT2JLwFXU3Mt0rbaAL
fgDbSEWeypirxVz34BfbQUG+32RiCMqg66tkD0yrDhgv15X2AHr5wRAKM2S4Zcjx
7MwRyVwKmZCPM4cKs+bSXii85/LekH7wuU8Zvce3EtvmNUO4+gchkkpYPIZ3XSuo
IyS20/WvXT/Uei1CdeXA+JU7QPjB6gdoRS8R3/0vo63ovAL7KcfaTM0CA1h4ymvR
7QPgwZuqMy+XntO8a5+zaB58E9lvH93ZMusQZh8MPpQGmflSYQMbu9kdjiuO9ZS1
4yLgv0q44q2LEexT4ukch2YyplL5csXtCbQ9iGrzyHBb6vrn0/B7X7SmL80EP9Ah
vXGspu6+LG8/PICLnEMovLeN/kDpaa5F/gR4LI5W4T46ShGjCrHqjSEhStOuaUOy
fCxKs41Rk7w0I8B9+9o2b/gMEcFK3L8xld3ybreoBIXhXBAhyp0KZr29KtvyY+Of
4xBXw2sjGSN9YxFrXYrymATiHYXzGjPDfF5m1yQsSEvxw0Jnh5YXYGvBVVV+VSFX
P5SsXIf4nXIuAWFKn/r+/tWTe/8Iw54BjQUWC2AE3YNnHIsDJkQRnyIGVlmU+ePb
8/gLCAQsbIngQMxh2PWgEJwbOQZfLra1uKjZhkAdoEL9hZ3IgoGxeEjUdczp1l/u
H4TPOS0Phv6WzqCT7BMavTjrP+rfW7hAOWaQhDyIknU7FC3fyjWp3+Q8D88gEq6X
axGIa3czBxOXRc/5EfRRnvQEl96yuUY0CMpjpdrhdtVBls2Sw6IUqznuREkDTbvN
2G6iq7/zA57fZtDP/bLayE3/uDNAHKC+x+fEhsOfIAe0w3Y7muwjxwiRclDq/lWP
7EYrxTDDndmaZHyamzz/mNkiydGWjA9PxiUPn1aGlk8DvrNXuv8xMdFLN3TPAm8f
3AvIPJzKYr9JzQd0VpySYKby6HEGulZCgFdD02wTHRKhZVcEWSVJgNRJgNGLwnhM
gfFBxrAz4dhAfYuNFzMWLYYsEXm//YqUSCCmPbNuxJaW/bzo3T+shTpidzNvCuoP
NyccFhQ108OJjmdaU7BFCKV/eBKNbHyb3qA4ejcZNdUCjBEL3cNqfByw3kzZt7RY
vy3Bk+U9yDkhfSy23EuuilyMjm4jBj2lPQQEX64xgmuFfFckY5t5zWkxfO69d40w
pjxz9FFXCn77okp8kPS1Rmyk1LHMBHS3nXy1vQJPlV+5zSJVIpYnlk/VSN06LCGt
QGs9IDli5TNhy2q+tWFhLrWvkIr0JPjVBlYzDnkWiOBGyvnTUmkNULgXftoZbD/8
iJXN0FDOYU24y51r/Y0hVrHaRd8B5GfAB0Bbkf2LkBiNZxd2QGEM4nYo6vmk9XCO
XXlIaCIfZezgknIcvm/ccNirIH88nYtksZSckzHoRTbky5c3hz8AvgSqgvHrNwyp
nPYq1EayLk4cyA1N5rrEoNlP3uog6MoBgFTOzWyDIBP+5R9ze4b6EuIGTG2pA0us
PRmoylJcdvAQhhYNhc/4pXE45V+J9xJGjJNj3LpypGw9cYhGavvR//C1WqZ/n2H0
VOh45XEYaxfIZQNfTuweygEBNPSEh5HhGM3k8zfjhmPhiXj7YcZKQqoE9+PZVjfu
1ThKgtV0mapRu4Q5XT1oBxGjb7I7pWmaxD2knqPG/J4PLSB04LmxZjh33j/NV3VC
xOM9exc4xtijQ/LfBaF9426yD8n0k2G8L+x3ATgbzy5xN4V2ULpoq0ZZqk+8b+zD
eyMDV+VYhAQg8HbwpNWo8p/cQQuzMhhO7fjFsYlolOOZC7eYUi04GH2Zq+iq7OMY
axM2yQMXelFJEjNeCj7dP0Q/tDHVmEAfEo0GisCN+R+AAyzyKgkqLUhxaWcaJr41
XikTLwUI1zChGmMfat+/Y5WHlnmiBb10lsrwSLRJ9vhTE/rEixwg4g+l03StGCx/
1wfe4bMYtHRw3jk8nPUQNXsh0v9/pETScxCV9S6pvGdBF/RNAFKZaPv+nKbV0HuO
slfkqtzpaICDO+/OWykeV0KU+Q9HFn1S+kGW+wwHJln8m2wuPsYQaoQCNttgEgH8
XAWB3yFpRlsehuZZSTCLhl6GZFyCEIA/smUeSoraXf17oya6u8SLQwZ7G19hMQWq
12d+1BgayMUiSGjWLhAZjMVIv+FmYwPGHDctTztQEZheERjaJrNppcP77jy8YQ1O
45P3A9wslyvuetRwy4mpBIcrGf51NrDmJ4qFbN8biwt3p+SSlIZA5MKB/7/m/rsj
MHShFj2pwkZcXtBy+d/0dhdfyvY55wtQVSUpkGt8B+WJhiIhYGDzbpZwq+vnjKqW
J6mrRIYS+L9HThGJCYcfzgHHaPVOWkW+Z8AEnx3E3hEk7HjwqURTRBtFL7XWW5kV
TCWdc9ypP0QlaYDpgvGoUGtI1okdqWb6tt2gYAIDjzgoX1c3yBheh5fh8IMe1Uf2
NiC7jAVF/m8vbjbKEnDRYCoe5zGEZU3j4AY6Ot43cryPeml3zryQyNM5fDTjDp6G
fHkDhm5jn91czgNhPaVJ0BDSTZAOkjCYFSsTWEwgldisWa7k4I4bw7adqzP574l7
dHKtjWE2DspNTc1IQbiUT4YslhIwbB8rA+8qsf0grxF2j4nXVcAOWgBYUBd1zSEX
n4iYejERlASpBnd0Vqy5Bv5VIZuyrhD0BcLXEl58+pWF74KTULzC3HI3rCHgSgWs
inRihAZf6fe10Tu1N+pVzmV7jfDWj+Z3IdVUqKDn+y3BDnWmywh9DjvOwedlRbG2
zhxOilRGnv2IJpwSqhE7cd7Rj8QFqgeq9zNJUTwIA7+wT66zRLVix7tt7Q08R8L7
O5MwBPr0TSQML3x8HlpQJbNlylbXiUobOBpZhkZX4500/fh8VdtVBpkatu+RN7vr
kPv9rA7dV3Oi8uW2WkaLjnAIPNkugp6i3gt5NasVu/do/Mc/z+zDjNj9e+CMgrtD
bthEUcGio2B3kULpHR5pq68H5MHORrbvVNzQH9MNzqjGqQd9uG/+W89o80p+ms8E
aS/QWeJSb5c1ximobvL1/613xJEwEDIWAeqYdndU8eeQM/VmujYzefHEY+l5bCLZ
0/Ny4wW+y+NwSSo3Cf8vDayKR5bN/LbovODKPlXsH/8ggnlNHVUGh/t3A5m8Keti
2UukvvXmLvOiV0ANslrRPq6IYvMU2P0dFfmuvE7IS0LYXVI+NvkMFF6IZrOzifBr
/IWvLBlYPoEOq/3QruHXrlefNIHLqF/jeidHmxDTUMnotDnaP8cKYN7pZPcI/YV5
nANLUAXmdYD264J0lGWkhf4n+mdYc4ssm0Z+vqewtRxeTunVvAvbpIiejpkx3R/A
UXMVCCQXf78DXPptVnn/stII+i7SLXKuTrYk6/Yqn84ElYYknoy9QYp4stdDDSNH
L2sdMU159DLXxNa4IS100Jp6F/PLx0fuozTMzsu0PU+srvmI9PFejkdqjOBO97bb
keL0lYwf/pTApes7IN4LQaOaNNemEupyyxyxWxPNzYC54Jl3BgESxxWjKbyX7Twr
U32/4gO15M8B4AyGTP/WNuLxsjUP4x5XHzoOKy8oEfIMZAC/enfQybnkwJzH9gux
sG7jK796ID+uybm3+hUjrfFJWCujpRjOqrvmbODd+ipNHPSgC2YtnFdLGviHRWWB
w+urgP9knO1JqnTYLwTlavek+qn1IGAfBYvSKOzHfDkKF0nty3DtrkOLO5l5loKd
RwHsCB1DgtMka2BykRgGGE6x535ePbaXoZ5bSvUXmGrfCaSW+ocgnW2/8hkgPUUi
M43NBb9PW0g8dMKke6oGuwPh1HM6o2B9t5oTl4GIOVgiNsbkmE7wxVI8/GgABI/2
vO3+67qnOfzXz8olVAJlRiKLwyvzmUdDtRw/GMdcp5t/cLGZ31+zc/a3cKB2yNYI
/k/c2eVqcFgvaUkUXFGGJovrEK+NB7X4HyLM8VHop8SgqT9Y4elvSb9aVom1QM/n
eg++XVeHd43Ba1xeWbFdg1Fwa2aiTs5zgWII6FzRXz+wKkd6Z0yxtzcYiSutNqlb
ItgONG+0wCYzyuEYrwY70iKDY4UWjO9ngnmoJUTtrepseNauG9vyOcSl7FkyHA+k
+dKGagJsjYXNlDyn8VC88okpx2I3HtNM4UNTax1W1UPZ9PuaI/8kdxwnP5/fvmMl
ugaAReJ/RbLq17L9bjMcdg==
`protect end_protected