`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 1664 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/9huKRhRMtvnNqb3Z+UU7TahEoHV+T8U3P3ufru7l1O
3DlgtZzb9QxCbOjthp9+wDkjygH0eUfDrEl1ovhZG62qmN4wNbDfzinW5GbKrflw
b3mKFB1glk7KpB39UX5PHiue8ECVD+dTO8NWn1nPOJ6aG8b1wgqS8+geQadefXju
3D+wkvCc80on0+xXYJG/tpUR/Wm9+JP4jWfFP4n9KgMbFzyU1oDznFJOtwCmYnAo
gSQi/3FiP610au7PHNNZaqc+s97FZG+yRFCRO6hJmreip6TGuNOVA2Wm9OtpFyNY
qkVEuWzqSSbQEXRrPdUObuCve2q+Ueelh3PJrgiDW0XHUgZ4YbgURgzaMbqRgrZE
VoIa24RDGIhvMEEEU9IMwkX90DGRqeDIw61UVIXnN6DgUr/GdrgfZWqr0HgbB+MZ
ttIHCEfDZ+9vyvHWysj836D67nrbRAaGGL8XwSGG79GV3RlIZqhhsSimg84rd78O
9Uv18bWET6iWAHgEJzBt/76ZFzpBst1JaxTAKOS48+00J0xxbi9ezbRY0FkyuQkI
TGNyP59AqLldKQ0xqRlaWGMo/8/Ajse7CihOJDFf/GVwKmSpr1xvJtkkyIzcwsla
3wzoKuNsVsNSQuens/sqRvL7zpwx2ZFSVNU4+LyXAuwy+IKGM/e9YqI0Z7WYaPXp
1L+kf1SD7A47Gj7cGvk8DE59Had9elLBUa/fEvJ2otw5h0+nrgignzy3mIKpEqXM
FZPc+pmjtYmwRLqc4s5etlldZTJR4wEHQ+BQjbJat6DpBISrd9w5DUuZQ0Am7pdX
8vr+lNAmw1Is4zGrMu7J5zA/N61xbHKw0+kTK4kbhqpG9aXqBwi3pkuYeTvv2p2R
fNaFKq9IwvAxABw8jsYBSGLeea3xbxAHFWep5ZjWxUEnmhJq7rw9kQgQxjl+xJdb
1oIy2ejwFkXbpJGVqZ9PBN2DPB/JfW7+iVv22H89WDFoOn2pcG3Rirv8JSzYIVv/
Q50zxFkuUaYCBSjMei6hEFZxz1wRMmE+e5nyu1G0F+yygy69ZvmTzgF4xS7TQT2R
fCvsMqFXFnIjk2/lQTSkRnhmbzCrkj6+Auj394G/GfGiZC0c0heBznfXVOVoJtWJ
JCwGIx3PcAxy+CSQoqjpEhnj0sJUkQWf+VBbYbR01i8icKDzU8W61DN80qjjjkOD
Wgo+L6xobPIEbWaaVoBbfgF37e/GelDOa2j98LVTw57JOuTp2YXIFP17eDAlr5OU
/kQvSJoua2bi24Gx3ZxwGTHrbj0g8+ASgz5tXMAj6wGg/Cow0z0fU5qnP37Ra7EL
0Ovx7SfceHC2UYx0outcPaMEYkhDHWGvE5qx9pOeNgdgOt7kp7vVSaFD67zBb/jG
I1qnhmOyeiFQk3xkXyHibVv3NoHplxBHuMqeI5zT2RrMAOcc1GOtzVUOJRaSsqn1
OcKHvEFyHtC9xgfERXTiQ5R3ZsE/GnCl7oy54dhoUgN8lUir3GD6tnRnNvn3C6yq
LvpZuNWIFNQbCxaTmkMvsOmLgCokUtJwv1zD1qo3N+YEJjmbNmx/fBXmfm07IgBG
eiGY21HXS8DcvHK3FwYY4PI05nOGLD5UurSVpZyvnG40nHxvBG7fICRaykLVmp3a
u7kdsI0RFFhI+zR/UIhpGlAz1JWQAxVxJbI2zxOTbKDhujQ3wdShrwiSNHIYu67a
IYqK1/p0n0fF9sxM6lzehXf4GRIb+EKDewepLuYNGJUPflwUgu0N8Zx5nWGIHX7L
adrEV/rdjaDTLZ5oqK2nKxvsvU9wYhOQFBbCJ5FWp05Jm23YsGF+hbt1ZloHJC6s
GQzpM1F2ACG9tuEi3wrN65BTyqiR8wqvIYGKl3vTC8WWjx2in7/uGa5HnzETlY44
z8pUY7vAqaZM0SkNAN8Vt/bXnvlolYZylPh0rPS4kFHbmZxzJx+bl9BEPQBcYDNn
NYfAgW2LyzlIJ6uP+Zs0robQ98MbPZnL3sO/i2Y26n35oVFR327BCWTVNfDdXH26
bi3x/+7Rbcc50NrAQKJYFO0dsMXcQ/HwjrPvt8am//uO/5+FUnkxV66qNryWcEdX
gl4+K1qeMz6ei0v3Dm0SB1L3d5DkjkmlsK3f/WOgjjk1WdBUIxThB7bqU45ZQexI
Jnerq7l7f6UDdW4zTX/UNWIG1yTEr2r4aPc7gj9tMLs=
`protect end_protected