`protect begin_protected
`protect version = 1
`protect encrypt_agent = "NI" , encrypt_agent_info = "1.0"
`protect key_keyowner = "Xilinx" , key_keyname = "xilinx_2014_03"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
aJ8rBNnBXqlSdSQu+M9/DYpqd770dYRDDW65r0u9FqUexGLFjbBJDxX7pkBVyW2I
o9U52aSv6YAvzjtrSjibITrJ7/qZbHqgcDAjHXN9Lwrq6o3xS8Oox9g5jGOvX/p0
S3e12h5ECqszSDH54GTrAr7D0LmYxGosqwMcwTC+hXuzDZaiQvA8S5z079eKUH9k
B0oA5dXw8g/6NZLZggtNYsXQySJbR8kVjEkrAx43pttEMH/pOQKpjZ0ZTYv/ZH8F
pipOfVrk/ptH7V5y3Ald2SXZ6mcvrjArJpzo9S3pVgF/UhiH6xYqC2bRR4mgO1co
3VNs/FJLXvxGL/2xUlIN8A==
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
hmxfTqYVgEqBNj1APNEo7B9SMhyrhRLWFqbSZdYJTYFEqgLSLI4/87n78IoKSNQ3
Xw/ws5J7RkOcTnJAzJ3Mow0O6JcP8fvhM9LN95tgDRA3vekisbNbQrW4fzzf+ixG
Hv5hGNDn7wlmxuCAgBL6y1WTGUQjN3I25tftzqFLkq4=
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 3200 )
`protect data_block
XAYzcToIY1VIPqVIYOouM/59UwEX+aE7FohaWu0/8IpTj7mav863zUNIsgIH2BWb
Abd9opeuBjbGF/waQMI2vMJTwD1ie1YueHc3nSNpEh4OXp8P5ybZFY89uyGz3ztU
W1EsuUnchJoQgbHZ/sLbgtGRgsrAFn+ZoIeGN1d6RAF2wAESJmYP8zw+p00RvjZ5
g/irlrcvR5923+bWtjXsfz/a/DCUZ8xN6/YxzYsqyHbsI/LN60u3V6g955Cft26V
r95fWj2wFgjLgbsjnGOW2XltKQpjoiHl11KhQaFUB/kFZdqT9gpgq6f8BHDueo18
5nkEFIWTvH4hCTcc+nl5NHf1PsQeHQdNLGnMZkxNjRqVMp5tUlK7Gvc8E6O7ac7h
Rsy3wgMfxJcOKB+VxKz5SHZ42OrB+EDqQ9vIa0r74j7UL9uk+ENyAC+RVHfsj6lF
J+J06WLBtJTYhvnzA9cISSH2Kqxf/a1QMGoPJ3wIOlA95I619d6Ymbe54vuiJwQN
e4TXVQqzYx2Wadql4hQfmBGdJHJBatszhXvAHZ34XUGyLKoC/vJgsZ+ylr/CCUmi
avsKRsvdOaiE/5YgngmwgYXefnt+g4mVVmouPKwjuxs+OvbLG9TJWxXRPExcTMWu
K+K3mr04TJlpubufOIhepIIkTktpP2Xgr4IALsDPHDVgTJG3dOzZq0uR4hWPfQY4
HcoviupDV9srRGcDMbuDQtOLkKcbRAj7YTBDpfJwJx2qvuVIrkZ8C/oaa5cA525Z
PTIaumTPL0xKOJxx5m3PRZtmS3vBMDGFL/5YWfSHd1mr3ySJhm0DgfS/iEBT/akm
pgWlns7wDxmfB928O97HHlsnSvoNgfuB5klXrrBpmib83l/eJwhufZA2jwSUWdMW
XxWxwvznbnlayIExwrApQUnX8us6rfhaIMtVACDzWvfkXqQvISA/Y5OI7dIINPLZ
MmwqmxqAxvEo8RjFcaMjdJ9dYDJOUuTyPvxx99MlR0Oz3AwBsxHrchLnfurIYjqF
xKBNYFY7liaF6ZXzT/XgXEvtN78uItGrsM/AzN1o3A88/mRHnp1Dmqzf2YxxLjZC
rL7Ysa5gOSfEn5kodMaMZoGMUjh/2yu112CWsGcYCG4vgD8wIJdX0dIj9RNkVhzj
ow/kmC4faGNfv9jikkS94MPZQKwSXrCm6ZIsOOBUP/Igd4QRnA9+c9edoQJ07lWE
bgps2Zc91egQ9WTk/wbI9p32qZKUjf/xyv1LqoHvS5/kAFQ/YLLG9qccUC+I3L/4
wA29CV6c0T8DQVVXgdkQbESKAYVny/haHYiZ2uN4gE9JZyfVa/+8ZcBH1jxZvJjE
5EnTSCszZZ7Ul3Q9+fkZSHMHQLtccV6HvdiGavV1cG9FXUHN/tAND8gEnzHmCJ1H
BZovAU/1MvWZug9opXAkCFb1Yf7HMzpmrHCq6uKFgJXH9dbi4bNPQF0vAoARV0j3
fhhKXu1nMhOSH6O/IqDHfYgEtBw2M/xmyoDQkHlXFva0VfBp24s8RRiBvB6wVTS4
lOZ+w7mbbWr6NQMgWGIlkG2mFIyArClVJEeHl/nB+9XHf2GRSOeRgJ3aRxuYcscl
LlwV/1EyZNsq4GWYkici6HW2ScfbKEUhiFBwZ5K9I9b0J/s2iR7w8M3T+J09Ainq
ZhKNc4PLoYvnRsBkTI7PAhEAFXFeIEqI9LoZQdXr01xdGDqUVxUk5UCDv5FEbj1G
AoFsZWyk3CP1pmQLfXGvpxkz+VzcmcKNpvCQGUFfjhV2h3fREhUzhSnUqzQVyGs8
vg96z0DFzwZ6r4YWBlHXEhBwn/BKz++mAJf/+yjrdAmmt2IO1TrKsxciK2fuEAIn
7Re/MNZpHPv9TbdRbJxpiqyGaJ135WYFm7k6uATmFAnz77S0HyO8l2CUShmT8ctO
D/Wh2hu1MHKdltAlGeEEPiQd+2LDfJGWx16k3zJwvDfjBehK5cU9OjXTIP9wTiom
vSHif7h6RhIESTWKJgxaj0gmpXBc/UnQaqvO9QwVo6OaPivjMj0D6ygXc2gr88Yu
6O7KnDlJ9l9w1wM6/A7YQbUZ8yv9biBi5sya/BFWoLfPrE2w9NstV2gPyfUKuO96
JBZ1Mb6Y2NtNlL0c+PMogfDmc4WWjLZY6gvshtuNxDxyirhxKmv7P68Njv+i2CPh
0jz5DS7jgNvH+6gTwgLwe42iLaB58+ccp+axSFM/5NjEwleWgJBC/91s0iDUez7t
YJcEB+az/cVJ7A19144KhaJrLdaFa2GycJAjppDfP1J6d33UoooYvMBHItKrZkMI
O0MCtPslrWydc/gVnfhyaZcUNVILhvbgrIjTEUkaDojjylIaSeT6rclp4oT2+bPM
3TJ1scmEAbqOqhVHBZTkG9RBcz1NGTKYZzhHLDXR0PWPnDHzggVHLprxQRM+5Q7E
6JSROy+UIv74NGVq2XYwRIevRmMVQOG7Lr/jipDubGcsor+bQ8S3OPTVaeKg28ud
123mpKTrSoYNGw9nW/Vi9La8PMzqZ4nhvF87YdJ3AElg9J+Kw3yTUVCPW5UPQ5Mq
cT+djZI3PDC4F19oDx8Ohs9ixymQS8D/HQnGX5hXxGmHmMjgeBov4aZ5RqcK5kAD
85FuOwlkpPp2U1IBMM62XFsZj9d875vfhozfDZoSUBB+nfSZRkeRaV7/zn/O5gKM
K4nJqM0gQpVLoK3jXQZqrHFX5bvTRyaJTzA89kejUEpuFfiiRvMCw/Pu6ZXpbkc8
nUvA2TYDuF5eQRp4gJdEaAH7HzDXmkF+WxgQc/KNq0joI5ijPtaHOgaGmmpnNqCo
TYD7K/B4wIMbD2YyukWIROZX4sjHrfj1vXgJaP/a9Sr2tniEXIb6jZ8RoZU3ZWOx
cXsOQpEJXNm4GsXA5wqp2izLqt1Wt1YBLc+SVsad0k9Z5DKBLT1Bx2M4qWUp58cY
+m/a6ZGu8Iec+00D+B1TEXrWEFr29Pr9+qv1ZyBP9PGcwzhwnZR2qxWoS7ODFmqN
J9CYqeDHYVSul+Uh6E1zAUBoccOXtT0j2wl/19BVDyUUyBqU45cTj/z+ADSoyJGN
5ZGnOj5SMo2srIYdrT50my6io4XA9EVdIZHNdAs3iwJxI2WBWn9IoKz6Gsz9peEe
AjwkISrl4Z66yoW7Gdf/juN6lFU9RmmCsgdR1bZ+AWclKURNYRRtywB7VQ5bHlFi
TJlcnmoL72X2cQfraCJn/JNElW55Ah7AJI4cGlOKe5/wxxW/gtcO6RZB76GraEti
vlNCZ/MNOM+EswU3ffod2bM7AExCrgc44k5hl15ksT2g+0mHHYG7WB5+tK+6lEZQ
OMCBAcnk7uMw6VUMr6o+76sau1DE4YTR+XLo5/rNWG3thRlqZrMozE2n/cTR33BD
phKv2qey4Vpm5MLnn5p5aitjA3plTKiXLZO1SIlFG+TFxaSGyykRIhzeTJGK4r/+
zRXdWKS8Vk1iIgj/zjrRuVaxMfShfWQVSSqQ7T6A5bhMS192ge667/WaoQv1AvJK
LsQVLlbP2XTJ0tdMqORG6ltQvZicGGerZQLqfUErpqa0IgwKZ47JH5qk6EaFy5um
NuQzi7KJt2dviT9GQH0JViog1gJhAev6/OW0LHoDDcdW/9DfaAwUbb5TKumKte4s
4cR2MkxlSxn5mbKRgvD5p/Qi21+mJtVCDJGo91i9APzAARbWf0J+PYkWqorZk3ca
4fhr9NZgrvlzn/hG/RsvBxCeKECPorAB+twvel3oqMpoRl3+JIFP1qiLKdmDxEXi
7DYKG0HeU0+xv3rHGAuRwP2bQiSVKUOaOCe3MWumJNecNsbV9NXTW5mqWxUsWtzS
dCg4GX14Q3ow275X7OrmrLiB8yfzB8Aq9iXBUAjHStUUo/MDib0RV6SCRphPgko8
JxgheWAFY8ve0EyR1HlQD4zVxc379+o4TeU8qMsPrCCuqQ77xhP2SCtMNjvKZcAr
TnoSuC27mnggfloX6HIhD8uB5dyafY25KhGyWo6GFgB6mj5s90n5VGekpzobuVub
3dJ/pFtrBnZiQgyc/vPfAStDVRfvC0bs/eC3aEN8uC1ECntYfsRnuPdDV08aYGBS
sAvl9bq5S7sKcPOCaTsgM2t6wnZYdcr8AigQUOFvZZ/UCbQhe0sJZCdjz8vUzXuD
lFXVQr6Ozfedw1exhSAhXCNMpjrUFBUvfBBFpqxHN6zOUTHu7kENqbt6wSeGbpfc
WZhJCPFZ2KftlcmbvFgoXR4EggodPPZSxGDAsAWvy8E=
`protect end_protected